-- no model for tie_diff
