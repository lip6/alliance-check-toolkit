test spice model
.param temp=27

.lib cornerMOSlv.lib mos_tt

.include inv_1.spice

Vgnd evss 0 0
Vdd  evdd 0 DC 1.8

Xinv in out evdd evss inv_1
.end
