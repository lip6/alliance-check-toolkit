* Filler200
.subckt Filler200 vss vdd iovss iovdd
Xbulkconn vdd vss iovdd iovss BulkConn_200WNoUp
.ends Filler200
