* and4_x1
.subckt and4_x1 vdd vss q i0 i1 i2 i3
Mi0_nmos nq i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi1_nmos _net0 i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi2_nmos _net1 i2 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi2_pmos vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi3_nmos _net2 i3 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi3_pmos nq i3 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_pd vss nq q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mq_pu vdd nq q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
.ends and4_x1
