* C4M.Sky130 logic transistors lib file

.lib tt
.include "C4M.Sky130_logic_tt_model.spice"
.endl tt
.lib ff
.include "C4M.Sky130_logic_ff_model.spice"
.endl ff
.lib ss
.include "C4M.Sky130_logic_ss_model.spice"
.endl ss
.lib fs
.include "C4M.Sky130_logic_fs_model.spice"
.endl fs
.lib sf
.include "C4M.Sky130_logic_sf_model.spice"
.endl sf
