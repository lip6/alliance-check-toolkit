* SecondaryProtection
* SecondaryProtection
.subckt SecondaryProtection iovdd iovss pad core
RR pad core 241.0
DDN iovss core sky130_fd_pr__diode_pw2nd_05v5 area=3.6875e-12 pj=13.68um
DDP core iovdd sky130_fd_pr__diode_pd2nw_05v5 area=3.6375000000000002e-12 pj=11.2um
.ends SecondaryProtection
