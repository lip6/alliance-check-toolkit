-- no model for xor2_x0
