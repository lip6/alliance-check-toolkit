* Coriolis Structural SPICE Driver
* Generated on Sep 30, 2024, 15:38
* Cell/Subckt "mac_cts_r".
* 
* INTERF vss
* INTERF vdd
* INTERF reset
* INTERF multiplier[3]
* INTERF multiplier[2]
* INTERF multiplier[1]
* INTERF multiplier[0]
* INTERF multiplicand[3]
* INTERF multiplicand[2]
* INTERF multiplicand[1]
* INTERF multiplicand[0]
* INTERF clk
* INTERF accumulator_out[7]
* INTERF accumulator_out[6]
* INTERF accumulator_out[5]
* INTERF accumulator_out[4]
* INTERF accumulator_out[3]
* INTERF accumulator_out[2]
* INTERF accumulator_out[1]
* INTERF accumulator_out[0]

* Terminal models (aka standard cells) used througout all the hierarchy.
.include tie_x0.spi
.include rowend_x0.spi
.include buf_x8.spi
.include sff1_x4.spi
.include nxr2_x1.spi
.include xr2_x4.spi
.include inv_x1.spi
.include a2_x2.spi
.include nao22_x1.spi
.include na2_x1.spi
.include na3_x1.spi
.include ao22_x2.spi
.include o2_x2.spi
.include a3_x2.spi
.include a4_x2.spi
.include na4_x1.spi
.include mx2_x2.spi
.include oa2a22_x2.spi
.include noa2a22_x1.spi
.include noa2ao222_x1.spi
.include on12_x1.spi
.include an12_x1.spi
.include oa2ao222_x2.spi
.include no2_x1.spi

* Non-terminal models (part of the user's design hierarchy).

.subckt mac_cts_r 0 1 2 11 12 13 14 15 16 17 18 72 74 75 76 77 78 79 80 81
* NET     0 = vss
* NET     1 = vdd
* NET     2 = reset
* NET     3 = partial_product[7]
* NET     4 = partial_product[6]
* NET     5 = partial_product[5]
* NET     6 = partial_product[4]
* NET     7 = partial_product[3]
* NET     8 = partial_product[2]
* NET     9 = partial_product[1]
* NET    10 = partial_product[0]
* NET    11 = multiplier[3]
* NET    12 = multiplier[2]
* NET    13 = multiplier[1]
* NET    14 = multiplier[0]
* NET    15 = multiplicand[3]
* NET    16 = multiplicand[2]
* NET    17 = multiplicand[1]
* NET    18 = multiplicand[0]
* NET    19 = clk_root_tr_tr_2
* NET    20 = clk_root_tr_tr_1
* NET    21 = clk_root_tr_tr_0
* NET    22 = clk_root_tr_tl_2
* NET    23 = clk_root_tr_tl_1
* NET    24 = clk_root_tr_tl_0
* NET    25 = clk_root_tr_br_2
* NET    26 = clk_root_tr_br_1
* NET    27 = clk_root_tr_br_0
* NET    28 = clk_root_tr_bl_2
* NET    29 = clk_root_tr_bl_1
* NET    30 = clk_root_tr_bl_0
* NET    31 = clk_root_tr_0
* NET    32 = clk_root_tl_tr_2
* NET    33 = clk_root_tl_tr_1
* NET    34 = clk_root_tl_tr_0
* NET    35 = clk_root_tl_tl_2
* NET    36 = clk_root_tl_tl_1
* NET    37 = clk_root_tl_tl_0
* NET    38 = clk_root_tl_br_2
* NET    39 = clk_root_tl_br_1
* NET    40 = clk_root_tl_br_0
* NET    41 = clk_root_tl_bl_2
* NET    42 = clk_root_tl_bl_1
* NET    43 = clk_root_tl_bl_0
* NET    44 = clk_root_tl_0
* NET    45 = clk_root_br_tr_2
* NET    46 = clk_root_br_tr_1
* NET    47 = clk_root_br_tr_0
* NET    48 = clk_root_br_tl_2
* NET    49 = clk_root_br_tl_1
* NET    50 = clk_root_br_tl_0
* NET    51 = clk_root_br_br_2
* NET    52 = clk_root_br_br_1
* NET    53 = clk_root_br_br_0
* NET    54 = clk_root_br_bl_2
* NET    55 = clk_root_br_bl_1
* NET    56 = clk_root_br_bl_0
* NET    57 = clk_root_br_0
* NET    58 = clk_root_bl_tr_2
* NET    59 = clk_root_bl_tr_1
* NET    60 = clk_root_bl_tr_0
* NET    61 = clk_root_bl_tl_2
* NET    62 = clk_root_bl_tl_1
* NET    63 = clk_root_bl_tl_0
* NET    64 = clk_root_bl_br_2
* NET    65 = clk_root_bl_br_1
* NET    66 = clk_root_bl_br_0
* NET    67 = clk_root_bl_bl_2
* NET    68 = clk_root_bl_bl_1
* NET    69 = clk_root_bl_bl_0
* NET    70 = clk_root_bl_0
* NET    71 = clk_root_0
* NET    72 = clk
* NET    73 = blockagenet
* NET    74 = accumulator_out[7]
* NET    75 = accumulator_out[6]
* NET    76 = accumulator_out[5]
* NET    77 = accumulator_out[4]
* NET    78 = accumulator_out[3]
* NET    79 = accumulator_out[2]
* NET    80 = accumulator_out[1]
* NET    81 = accumulator_out[0]
* NET    82 = abc_567_new_n99
* NET    83 = abc_567_new_n98
* NET    84 = abc_567_new_n97
* NET    85 = abc_567_new_n96
* NET    86 = abc_567_new_n95
* NET    87 = abc_567_new_n94
* NET    88 = abc_567_new_n93
* NET    89 = abc_567_new_n91
* NET    90 = abc_567_new_n90
* NET    91 = abc_567_new_n89
* NET    92 = abc_567_new_n88
* NET    93 = abc_567_new_n87
* NET    94 = abc_567_new_n86
* NET    95 = abc_567_new_n85
* NET    96 = abc_567_new_n84
* NET    97 = abc_567_new_n83
* NET    98 = abc_567_new_n82
* NET    99 = abc_567_new_n81
* NET   100 = abc_567_new_n80
* NET   101 = abc_567_new_n79
* NET   102 = abc_567_new_n78
* NET   103 = abc_567_new_n77
* NET   104 = abc_567_new_n76
* NET   105 = abc_567_new_n75
* NET   106 = abc_567_new_n74
* NET   107 = abc_567_new_n73
* NET   108 = abc_567_new_n72
* NET   109 = abc_567_new_n71
* NET   110 = abc_567_new_n70
* NET   111 = abc_567_new_n69
* NET   112 = abc_567_new_n68
* NET   113 = abc_567_new_n67
* NET   114 = abc_567_new_n66
* NET   115 = abc_567_new_n65
* NET   116 = abc_567_new_n63
* NET   117 = abc_567_new_n62
* NET   118 = abc_567_new_n61
* NET   119 = abc_567_new_n60
* NET   120 = abc_567_new_n59
* NET   121 = abc_567_new_n58
* NET   122 = abc_567_new_n57
* NET   123 = abc_567_new_n56
* NET   124 = abc_567_new_n55
* NET   125 = abc_567_new_n54
* NET   126 = abc_567_new_n52
* NET   127 = abc_567_new_n51
* NET   128 = abc_567_new_n50
* NET   129 = abc_567_new_n49
* NET   130 = abc_567_new_n47
* NET   131 = abc_567_new_n46
* NET   132 = abc_567_new_n45
* NET   133 = abc_567_new_n44
* NET   134 = abc_567_new_n43
* NET   135 = abc_567_new_n42
* NET   136 = abc_567_new_n188
* NET   137 = abc_567_new_n187
* NET   138 = abc_567_new_n186
* NET   139 = abc_567_new_n185
* NET   140 = abc_567_new_n183
* NET   141 = abc_567_new_n182
* NET   142 = abc_567_new_n181
* NET   143 = abc_567_new_n180
* NET   144 = abc_567_new_n179
* NET   145 = abc_567_new_n178
* NET   146 = abc_567_new_n177
* NET   147 = abc_567_new_n176
* NET   148 = abc_567_new_n175
* NET   149 = abc_567_new_n173
* NET   150 = abc_567_new_n172
* NET   151 = abc_567_new_n171
* NET   152 = abc_567_new_n170
* NET   153 = abc_567_new_n169
* NET   154 = abc_567_new_n168
* NET   155 = abc_567_new_n166
* NET   156 = abc_567_new_n165
* NET   157 = abc_567_new_n164
* NET   158 = abc_567_new_n163
* NET   159 = abc_567_new_n162
* NET   160 = abc_567_new_n161
* NET   161 = abc_567_new_n160
* NET   162 = abc_567_new_n159
* NET   163 = abc_567_new_n157
* NET   164 = abc_567_new_n156
* NET   165 = abc_567_new_n155
* NET   166 = abc_567_new_n154
* NET   167 = abc_567_new_n153
* NET   168 = abc_567_new_n151
* NET   169 = abc_567_new_n150
* NET   170 = abc_567_new_n149
* NET   171 = abc_567_new_n148
* NET   172 = abc_567_new_n147
* NET   173 = abc_567_new_n146
* NET   174 = abc_567_new_n144
* NET   175 = abc_567_new_n143
* NET   176 = abc_567_new_n142
* NET   177 = abc_567_new_n141
* NET   178 = abc_567_new_n139
* NET   179 = abc_567_new_n138
* NET   180 = abc_567_new_n136
* NET   181 = abc_567_new_n134
* NET   182 = abc_567_new_n133
* NET   183 = abc_567_new_n132
* NET   184 = abc_567_new_n131
* NET   185 = abc_567_new_n130
* NET   186 = abc_567_new_n129
* NET   187 = abc_567_new_n128
* NET   188 = abc_567_new_n127
* NET   189 = abc_567_new_n125
* NET   190 = abc_567_new_n124
* NET   191 = abc_567_new_n123
* NET   192 = abc_567_new_n122
* NET   193 = abc_567_new_n121
* NET   194 = abc_567_new_n120
* NET   195 = abc_567_new_n119
* NET   196 = abc_567_new_n118
* NET   197 = abc_567_new_n117
* NET   198 = abc_567_new_n116
* NET   199 = abc_567_new_n115
* NET   200 = abc_567_new_n113
* NET   201 = abc_567_new_n112
* NET   202 = abc_567_new_n111
* NET   203 = abc_567_new_n110
* NET   204 = abc_567_new_n109
* NET   205 = abc_567_new_n108
* NET   206 = abc_567_new_n107
* NET   207 = abc_567_new_n106
* NET   208 = abc_567_new_n105
* NET   209 = abc_567_new_n104
* NET   210 = abc_567_new_n103
* NET   211 = abc_567_new_n102
* NET   212 = abc_567_new_n101
* NET   213 = abc_567_new_n100
* NET   214 = abc_567_auto_rtlil_cc_2608_MuxGate_566
* NET   215 = abc_567_auto_rtlil_cc_2608_MuxGate_564
* NET   216 = abc_567_auto_rtlil_cc_2608_MuxGate_562
* NET   217 = abc_567_auto_rtlil_cc_2608_MuxGate_560
* NET   218 = abc_567_auto_rtlil_cc_2608_MuxGate_558
* NET   219 = abc_567_auto_rtlil_cc_2608_MuxGate_556
* NET   220 = abc_567_auto_rtlil_cc_2608_MuxGate_554
* NET   221 = abc_567_auto_rtlil_cc_2608_MuxGate_552
* NET   222 = abc_567_auto_rtlil_cc_2608_MuxGate_550
* NET   223 = abc_567_auto_rtlil_cc_2608_MuxGate_548
* NET   224 = abc_567_auto_rtlil_cc_2608_MuxGate_546
* NET   225 = abc_567_auto_rtlil_cc_2608_MuxGate_544
* NET   226 = abc_567_auto_rtlil_cc_2608_MuxGate_542
* NET   227 = abc_567_auto_rtlil_cc_2608_MuxGate_540
* NET   228 = abc_567_auto_rtlil_cc_2608_MuxGate_538
* NET   229 = abc_567_auto_rtlil_cc_2608_MuxGate_536

xfeed_6739 0 1 tie_x0
xfeed_6738 0 1 tie_x0
xfeed_6737 0 1 tie_x0
xfeed_6736 0 1 tie_x0
xfeed_6735 0 1 tie_x0
xfeed_6734 0 1 rowend_x0
xfeed_6733 0 1 tie_x0
xfeed_6732 0 1 tie_x0
xfeed_6731 0 1 tie_x0
xfeed_409 0 1 tie_x0
xfeed_408 0 1 tie_x0
xfeed_407 0 1 tie_x0
xfeed_406 0 1 tie_x0
xfeed_405 0 1 tie_x0
xfeed_404 0 1 tie_x0
xfeed_403 0 1 tie_x0
xfeed_402 0 1 tie_x0
xfeed_401 0 1 tie_x0
xfeed_400 0 1 tie_x0
xspare_buffer_44 0 1 50 57 buf_x8
xspare_buffer_42 0 1 51 57 buf_x8
xspare_buffer_41 0 1 52 57 buf_x8
xspare_buffer_40 0 1 53 57 buf_x8
xfeed_7276 0 1 tie_x0
xfeed_7275 0 1 tie_x0
xfeed_7274 0 1 tie_x0
xfeed_7273 0 1 tie_x0
xfeed_7272 0 1 tie_x0
xfeed_7271 0 1 tie_x0
xfeed_7270 0 1 tie_x0
xfeed_2437 0 1 tie_x0
xfeed_2436 0 1 tie_x0
xfeed_2435 0 1 tie_x0
xfeed_2434 0 1 tie_x0
xfeed_2433 0 1 tie_x0
xfeed_2432 0 1 tie_x0
xfeed_2431 0 1 tie_x0
xfeed_2430 0 1 tie_x0
xspare_buffer_49 0 1 46 57 buf_x8
xspare_buffer_48 0 1 47 57 buf_x8
xspare_buffer_46 0 1 48 57 buf_x8
xspare_buffer_45 0 1 49 57 buf_x8
xfeed_7279 0 1 tie_x0
xfeed_7278 0 1 tie_x0
xfeed_7277 0 1 tie_x0
xfeed_6749 0 1 tie_x0
xfeed_6748 0 1 tie_x0
xfeed_6747 0 1 tie_x0
xfeed_6746 0 1 tie_x0
xfeed_6745 0 1 tie_x0
xfeed_6744 0 1 tie_x0
xfeed_6743 0 1 tie_x0
xfeed_6742 0 1 tie_x0
xfeed_6741 0 1 tie_x0
xfeed_6740 0 1 tie_x0
xfeed_2439 0 1 tie_x0
xfeed_2438 0 1 tie_x0
xfeed_419 0 1 tie_x0
xfeed_418 0 1 tie_x0
xfeed_417 0 1 tie_x0
xfeed_416 0 1 tie_x0
xfeed_415 0 1 tie_x0
xfeed_414 0 1 tie_x0
xfeed_413 0 1 tie_x0
xfeed_412 0 1 tie_x0
xfeed_411 0 1 tie_x0
xfeed_410 0 1 tie_x0
xspare_buffer_50 0 1 45 57 buf_x8
xfeed_1900 0 1 tie_x0
xfeed_1901 0 1 tie_x0
xfeed_1902 0 1 rowend_x0
xfeed_1903 0 1 tie_x0
xfeed_1904 0 1 tie_x0
xfeed_1905 0 1 tie_x0
xfeed_1906 0 1 tie_x0
xfeed_1907 0 1 tie_x0
xfeed_1908 0 1 tie_x0
xfeed_1909 0 1 tie_x0
xfeed_7283 0 1 tie_x0
xfeed_7282 0 1 tie_x0
xfeed_7281 0 1 tie_x0
xfeed_7280 0 1 tie_x0
xfeed_2444 0 1 tie_x0
xfeed_2443 0 1 tie_x0
xfeed_2442 0 1 tie_x0
xfeed_2441 0 1 tie_x0
xfeed_2440 0 1 tie_x0
xspare_buffer_58 0 1 38 44 buf_x8
xspare_buffer_57 0 1 39 44 buf_x8
xspare_buffer_56 0 1 40 44 buf_x8
xspare_buffer_54 0 1 41 44 buf_x8
xspare_buffer_53 0 1 42 44 buf_x8
xspare_buffer_52 0 1 43 44 buf_x8
xfeed_7289 0 1 tie_x0
xfeed_7288 0 1 tie_x0
xfeed_7287 0 1 tie_x0
xfeed_7286 0 1 tie_x0
xfeed_7285 0 1 tie_x0
xfeed_7284 0 1 tie_x0
xfeed_6759 0 1 rowend_x0
xfeed_6758 0 1 tie_x0
xfeed_6757 0 1 tie_x0
xfeed_6756 0 1 tie_x0
xfeed_6755 0 1 tie_x0
xfeed_6754 0 1 tie_x0
xfeed_6753 0 1 tie_x0
xfeed_6752 0 1 tie_x0
xfeed_6751 0 1 tie_x0
xfeed_6750 0 1 tie_x0
xfeed_2449 0 1 tie_x0
xfeed_2448 0 1 tie_x0
xfeed_2447 0 1 tie_x0
xfeed_2446 0 1 tie_x0
xfeed_2445 0 1 tie_x0
xfeed_429 0 1 tie_x0
xfeed_428 0 1 tie_x0
xfeed_427 0 1 tie_x0
xfeed_426 0 1 tie_x0
xfeed_425 0 1 tie_x0
xfeed_424 0 1 tie_x0
xfeed_423 0 1 tie_x0
xfeed_422 0 1 tie_x0
xfeed_421 0 1 tie_x0
xfeed_420 0 1 tie_x0
xfeed_1910 0 1 tie_x0
xfeed_1911 0 1 tie_x0
xfeed_1912 0 1 tie_x0
xfeed_1913 0 1 tie_x0
xfeed_1914 0 1 tie_x0
xfeed_1915 0 1 tie_x0
xfeed_1916 0 1 tie_x0
xfeed_1917 0 1 tie_x0
xfeed_1918 0 1 tie_x0
xfeed_1919 0 1 tie_x0
xfeed_7290 0 1 tie_x0
xfeed_2451 0 1 tie_x0
xfeed_2450 0 1 tie_x0
xspare_buffer_69 0 1 29 31 buf_x8
xspare_buffer_68 0 1 30 31 buf_x8
xspare_buffer_66 0 1 32 44 buf_x8
xspare_buffer_65 0 1 33 44 buf_x8
xspare_buffer_64 0 1 34 44 buf_x8
xspare_buffer_62 0 1 35 44 buf_x8
xspare_buffer_61 0 1 36 44 buf_x8
xspare_buffer_60 0 1 37 44 buf_x8
xfeed_7299 0 1 tie_x0
xfeed_7298 0 1 tie_x0
xfeed_7297 0 1 rowend_x0
xfeed_7296 0 1 tie_x0
xfeed_7295 0 1 tie_x0
xfeed_7294 0 1 tie_x0
xfeed_7293 0 1 tie_x0
xfeed_7292 0 1 tie_x0
xfeed_7291 0 1 tie_x0
xfeed_6769 0 1 tie_x0
xfeed_6768 0 1 tie_x0
xfeed_6767 0 1 tie_x0
xfeed_6766 0 1 tie_x0
xfeed_6765 0 1 tie_x0
xfeed_6764 0 1 tie_x0
xfeed_6763 0 1 tie_x0
xfeed_6762 0 1 tie_x0
xfeed_6761 0 1 tie_x0
xfeed_6760 0 1 tie_x0
xfeed_2459 0 1 tie_x0
xfeed_2458 0 1 tie_x0
xfeed_2457 0 1 tie_x0
xfeed_2456 0 1 tie_x0
xfeed_2455 0 1 tie_x0
xfeed_2454 0 1 tie_x0
xfeed_2453 0 1 tie_x0
xfeed_2452 0 1 tie_x0
xfeed_439 0 1 tie_x0
xfeed_438 0 1 tie_x0
xfeed_437 0 1 tie_x0
xfeed_436 0 1 tie_x0
xfeed_435 0 1 tie_x0
xfeed_434 0 1 tie_x0
xfeed_433 0 1 tie_x0
xfeed_432 0 1 tie_x0
xfeed_431 0 1 tie_x0
xfeed_430 0 1 tie_x0
xfeed_1920 0 1 tie_x0
xfeed_1921 0 1 tie_x0
xfeed_1922 0 1 tie_x0
xfeed_1923 0 1 tie_x0
xfeed_1924 0 1 tie_x0
xfeed_1925 0 1 tie_x0
xfeed_1926 0 1 tie_x0
xfeed_1927 0 1 tie_x0
xfeed_1928 0 1 rowend_x0
xfeed_1929 0 1 tie_x0
xspare_buffer_77 0 1 23 31 buf_x8
xspare_buffer_76 0 1 24 31 buf_x8
xspare_buffer_74 0 1 25 31 buf_x8
xspare_buffer_73 0 1 26 31 buf_x8
xspare_buffer_72 0 1 27 31 buf_x8
xspare_buffer_70 0 1 28 31 buf_x8
xspare_buffer_78 0 1 22 31 buf_x8
xfeed_6779 0 1 tie_x0
xfeed_6778 0 1 tie_x0
xfeed_6777 0 1 tie_x0
xfeed_6776 0 1 tie_x0
xfeed_6775 0 1 tie_x0
xfeed_6774 0 1 tie_x0
xfeed_6773 0 1 tie_x0
xfeed_6772 0 1 tie_x0
xfeed_6771 0 1 tie_x0
xfeed_6770 0 1 tie_x0
xfeed_2469 0 1 tie_x0
xfeed_2468 0 1 tie_x0
xfeed_2467 0 1 tie_x0
xfeed_2466 0 1 tie_x0
xfeed_2465 0 1 tie_x0
xfeed_2464 0 1 tie_x0
xfeed_2463 0 1 tie_x0
xfeed_2462 0 1 tie_x0
xfeed_2461 0 1 tie_x0
xfeed_2460 0 1 tie_x0
xfeed_449 0 1 tie_x0
xfeed_448 0 1 tie_x0
xfeed_447 0 1 tie_x0
xfeed_446 0 1 tie_x0
xfeed_445 0 1 tie_x0
xfeed_444 0 1 tie_x0
xfeed_443 0 1 tie_x0
xfeed_442 0 1 tie_x0
xfeed_441 0 1 tie_x0
xfeed_440 0 1 tie_x0
xfeed_1930 0 1 tie_x0
xfeed_1931 0 1 tie_x0
xfeed_1932 0 1 tie_x0
xfeed_1933 0 1 tie_x0
xfeed_1934 0 1 tie_x0
xfeed_1935 0 1 tie_x0
xfeed_1936 0 1 tie_x0
xfeed_1937 0 1 tie_x0
xfeed_1938 0 1 tie_x0
xfeed_1939 0 1 tie_x0
xspare_buffer_80 0 1 21 31 buf_x8
xspare_buffer_81 0 1 20 31 buf_x8
xspare_buffer_82 0 1 19 31 buf_x8
xfeed_6789 0 1 tie_x0
xfeed_6788 0 1 tie_x0
xfeed_6787 0 1 tie_x0
xfeed_6786 0 1 tie_x0
xfeed_6785 0 1 tie_x0
xfeed_6784 0 1 tie_x0
xfeed_6783 0 1 tie_x0
xfeed_6782 0 1 tie_x0
xfeed_6781 0 1 tie_x0
xfeed_6780 0 1 tie_x0
xfeed_2479 0 1 tie_x0
xfeed_2478 0 1 tie_x0
xfeed_2477 0 1 tie_x0
xfeed_2476 0 1 tie_x0
xfeed_2475 0 1 tie_x0
xfeed_2474 0 1 tie_x0
xfeed_2473 0 1 tie_x0
xfeed_2472 0 1 tie_x0
xfeed_2471 0 1 tie_x0
xfeed_2470 0 1 tie_x0
xfeed_459 0 1 tie_x0
xfeed_458 0 1 tie_x0
xfeed_457 0 1 tie_x0
xfeed_456 0 1 tie_x0
xfeed_455 0 1 tie_x0
xfeed_454 0 1 tie_x0
xfeed_453 0 1 tie_x0
xfeed_452 0 1 tie_x0
xfeed_451 0 1 tie_x0
xfeed_450 0 1 tie_x0
xsubckt_155_sff1_x4 0 1 3 222 53 sff1_x4
xfeed_1940 0 1 tie_x0
xfeed_1941 0 1 tie_x0
xfeed_1942 0 1 tie_x0
xfeed_1943 0 1 tie_x0
xfeed_1944 0 1 tie_x0
xfeed_1945 0 1 tie_x0
xfeed_1946 0 1 tie_x0
xfeed_1947 0 1 tie_x0
xfeed_1948 0 1 tie_x0
xfeed_1949 0 1 tie_x0
xfeed_7409 0 1 tie_x0
xfeed_7408 0 1 tie_x0
xfeed_7407 0 1 tie_x0
xfeed_7406 0 1 tie_x0
xfeed_7405 0 1 tie_x0
xfeed_7404 0 1 tie_x0
xfeed_7403 0 1 tie_x0
xfeed_7402 0 1 tie_x0
xfeed_7401 0 1 tie_x0
xfeed_7400 0 1 tie_x0
xsubckt_18_nxr2_x1 0 1 119 125 120 nxr2_x1
xfeed_6799 0 1 tie_x0
xfeed_6798 0 1 tie_x0
xfeed_6797 0 1 tie_x0
xfeed_6796 0 1 tie_x0
xfeed_6795 0 1 tie_x0
xfeed_6794 0 1 tie_x0
xfeed_6793 0 1 tie_x0
xfeed_6792 0 1 tie_x0
xfeed_6791 0 1 tie_x0
xfeed_6790 0 1 tie_x0
xfeed_2489 0 1 tie_x0
xfeed_2488 0 1 tie_x0
xfeed_2487 0 1 tie_x0
xfeed_2486 0 1 tie_x0
xfeed_2485 0 1 tie_x0
xfeed_2484 0 1 tie_x0
xfeed_2483 0 1 tie_x0
xfeed_2482 0 1 tie_x0
xfeed_2481 0 1 tie_x0
xfeed_2480 0 1 tie_x0
xfeed_469 0 1 tie_x0
xfeed_468 0 1 tie_x0
xfeed_467 0 1 tie_x0
xfeed_466 0 1 tie_x0
xfeed_465 0 1 tie_x0
xfeed_464 0 1 tie_x0
xfeed_463 0 1 tie_x0
xfeed_462 0 1 tie_x0
xfeed_461 0 1 tie_x0
xfeed_460 0 1 tie_x0
xfeed_1950 0 1 tie_x0
xfeed_1951 0 1 tie_x0
xfeed_1952 0 1 tie_x0
xfeed_1953 0 1 rowend_x0
xfeed_1954 0 1 tie_x0
xfeed_1955 0 1 tie_x0
xfeed_1956 0 1 tie_x0
xfeed_1957 0 1 tie_x0
xfeed_1958 0 1 tie_x0
xfeed_1959 0 1 tie_x0
xfeed_7416 0 1 tie_x0
xfeed_7415 0 1 tie_x0
xfeed_7414 0 1 tie_x0
xfeed_7413 0 1 tie_x0
xfeed_7412 0 1 rowend_x0
xfeed_7411 0 1 tie_x0
xfeed_7410 0 1 tie_x0
xfeed_3109 0 1 tie_x0
xfeed_3108 0 1 tie_x0
xfeed_3107 0 1 tie_x0
xfeed_3106 0 1 tie_x0
xfeed_3105 0 1 tie_x0
xfeed_3104 0 1 tie_x0
xfeed_3103 0 1 tie_x0
xfeed_3102 0 1 tie_x0
xfeed_3101 0 1 tie_x0
xfeed_3100 0 1 tie_x0
xsubckt_137_xr2_x4 0 1 144 75 4 xr2_x4
xfeed_7419 0 1 tie_x0
xfeed_7418 0 1 tie_x0
xfeed_7417 0 1 tie_x0
xfeed_2499 0 1 tie_x0
xfeed_2498 0 1 tie_x0
xfeed_2497 0 1 tie_x0
xfeed_2496 0 1 tie_x0
xfeed_2495 0 1 tie_x0
xfeed_2494 0 1 tie_x0
xfeed_2493 0 1 tie_x0
xfeed_2492 0 1 tie_x0
xfeed_2491 0 1 tie_x0
xfeed_2490 0 1 tie_x0
xfeed_479 0 1 tie_x0
xfeed_478 0 1 tie_x0
xfeed_477 0 1 tie_x0
xfeed_476 0 1 tie_x0
xfeed_475 0 1 tie_x0
xfeed_474 0 1 tie_x0
xfeed_473 0 1 tie_x0
xfeed_472 0 1 tie_x0
xfeed_471 0 1 tie_x0
xfeed_470 0 1 tie_x0
xfeed_1960 0 1 tie_x0
xfeed_1961 0 1 tie_x0
xfeed_1962 0 1 tie_x0
xfeed_1963 0 1 tie_x0
xfeed_1964 0 1 tie_x0
xfeed_1965 0 1 tie_x0
xfeed_1966 0 1 tie_x0
xfeed_1967 0 1 tie_x0
xfeed_1968 0 1 tie_x0
xfeed_1969 0 1 tie_x0
xfeed_7423 0 1 tie_x0
xfeed_7422 0 1 tie_x0
xfeed_7421 0 1 tie_x0
xfeed_7420 0 1 tie_x0
xfeed_3119 0 1 tie_x0
xfeed_3118 0 1 tie_x0
xfeed_3117 0 1 tie_x0
xfeed_3116 0 1 tie_x0
xfeed_3115 0 1 tie_x0
xfeed_3114 0 1 tie_x0
xfeed_3113 0 1 tie_x0
xfeed_3112 0 1 tie_x0
xfeed_3111 0 1 tie_x0
xfeed_3110 0 1 tie_x0
xfeed_7429 0 1 tie_x0
xfeed_7428 0 1 tie_x0
xfeed_7427 0 1 tie_x0
xfeed_7426 0 1 tie_x0
xfeed_7425 0 1 tie_x0
xfeed_7424 0 1 tie_x0
xfeed_489 0 1 tie_x0
xfeed_488 0 1 tie_x0
xfeed_487 0 1 tie_x0
xfeed_486 0 1 tie_x0
xfeed_485 0 1 tie_x0
xfeed_484 0 1 tie_x0
xfeed_483 0 1 tie_x0
xfeed_482 0 1 tie_x0
xfeed_481 0 1 tie_x0
xfeed_480 0 1 tie_x0
xfeed_1970 0 1 tie_x0
xfeed_1971 0 1 tie_x0
xfeed_1972 0 1 tie_x0
xfeed_1973 0 1 tie_x0
xfeed_1974 0 1 tie_x0
xfeed_1975 0 1 tie_x0
xfeed_1976 0 1 tie_x0
xfeed_1977 0 1 tie_x0
xfeed_1978 0 1 tie_x0
xfeed_1979 0 1 tie_x0
xfeed_7430 0 1 tie_x0
xfeed_3129 0 1 tie_x0
xfeed_3128 0 1 tie_x0
xfeed_3127 0 1 tie_x0
xfeed_3126 0 1 tie_x0
xfeed_3125 0 1 tie_x0
xfeed_3124 0 1 tie_x0
xfeed_3123 0 1 tie_x0
xfeed_3122 0 1 tie_x0
xfeed_3121 0 1 tie_x0
xfeed_3120 0 1 tie_x0
xsubckt_0_inv_x1 0 1 135 78 inv_x1
xsubckt_2_inv_x1 0 1 133 11 inv_x1
xsubckt_4_inv_x1 0 1 131 2 inv_x1
xfeed_7439 0 1 tie_x0
xfeed_7438 0 1 tie_x0
xfeed_7437 0 1 tie_x0
xfeed_7436 0 1 tie_x0
xfeed_7435 0 1 tie_x0
xfeed_7434 0 1 tie_x0
xfeed_7433 0 1 tie_x0
xfeed_7432 0 1 tie_x0
xfeed_7431 0 1 tie_x0
xfeed_6909 0 1 tie_x0
xfeed_6908 0 1 tie_x0
xfeed_6907 0 1 tie_x0
xfeed_6906 0 1 tie_x0
xfeed_6905 0 1 tie_x0
xfeed_6904 0 1 tie_x0
xfeed_6903 0 1 rowend_x0
xfeed_6902 0 1 tie_x0
xfeed_6901 0 1 tie_x0
xfeed_6900 0 1 tie_x0
xfeed_499 0 1 tie_x0
xfeed_498 0 1 tie_x0
xfeed_497 0 1 tie_x0
xfeed_496 0 1 tie_x0
xfeed_495 0 1 tie_x0
xfeed_494 0 1 tie_x0
xfeed_493 0 1 tie_x0
xfeed_492 0 1 tie_x0
xfeed_491 0 1 tie_x0
xfeed_490 0 1 tie_x0
xfeed_1980 0 1 tie_x0
xfeed_1981 0 1 tie_x0
xfeed_1982 0 1 tie_x0
xfeed_1983 0 1 tie_x0
xfeed_1984 0 1 tie_x0
xfeed_1985 0 1 tie_x0
xfeed_1986 0 1 tie_x0
xfeed_1987 0 1 tie_x0
xfeed_1988 0 1 tie_x0
xfeed_1989 0 1 tie_x0
xfeed_3137 0 1 tie_x0
xfeed_3136 0 1 tie_x0
xfeed_3135 0 1 tie_x0
xfeed_3134 0 1 rowend_x0
xfeed_3133 0 1 tie_x0
xfeed_3132 0 1 tie_x0
xfeed_3131 0 1 tie_x0
xfeed_3130 0 1 tie_x0
xfeed_7449 0 1 tie_x0
xfeed_7448 0 1 tie_x0
xfeed_7447 0 1 tie_x0
xfeed_7446 0 1 tie_x0
xfeed_7445 0 1 tie_x0
xfeed_7444 0 1 tie_x0
xfeed_7443 0 1 tie_x0
xfeed_7442 0 1 tie_x0
xfeed_7441 0 1 tie_x0
xfeed_7440 0 1 tie_x0
xfeed_6919 0 1 tie_x0
xfeed_6918 0 1 tie_x0
xfeed_6917 0 1 tie_x0
xfeed_6916 0 1 tie_x0
xfeed_6915 0 1 tie_x0
xfeed_6914 0 1 tie_x0
xfeed_6913 0 1 tie_x0
xfeed_6912 0 1 tie_x0
xfeed_6911 0 1 tie_x0
xfeed_6910 0 1 tie_x0
xfeed_3139 0 1 tie_x0
xfeed_3138 0 1 tie_x0
xfeed_2609 0 1 tie_x0
xfeed_2608 0 1 tie_x0
xfeed_2607 0 1 tie_x0
xfeed_2606 0 1 tie_x0
xfeed_2605 0 1 tie_x0
xfeed_2604 0 1 tie_x0
xfeed_2603 0 1 tie_x0
xfeed_2602 0 1 tie_x0
xfeed_2601 0 1 rowend_x0
xfeed_2600 0 1 tie_x0
xsubckt_81_nxr2_x1 0 1 191 198 193 nxr2_x1
xfeed_1990 0 1 tie_x0
xfeed_1991 0 1 tie_x0
xfeed_1992 0 1 tie_x0
xfeed_1993 0 1 tie_x0
xfeed_1994 0 1 tie_x0
xfeed_1995 0 1 tie_x0
xfeed_1996 0 1 tie_x0
xfeed_1997 0 1 tie_x0
xfeed_1998 0 1 tie_x0
xfeed_1999 0 1 tie_x0
xfeed_3144 0 1 tie_x0
xfeed_3143 0 1 tie_x0
xfeed_3142 0 1 tie_x0
xfeed_3141 0 1 tie_x0
xfeed_3140 0 1 tie_x0
xsubckt_64_a2_x2 0 1 207 84 209 a2_x2
xfeed_7459 0 1 tie_x0
xfeed_7458 0 1 tie_x0
xfeed_7457 0 1 tie_x0
xfeed_7456 0 1 tie_x0
xfeed_7455 0 1 tie_x0
xfeed_7454 0 1 tie_x0
xfeed_7453 0 1 tie_x0
xfeed_7452 0 1 tie_x0
xfeed_7451 0 1 tie_x0
xfeed_7450 0 1 tie_x0
xfeed_6929 0 1 tie_x0
xfeed_6928 0 1 tie_x0
xfeed_6927 0 1 tie_x0
xfeed_6926 0 1 tie_x0
xfeed_6925 0 1 tie_x0
xfeed_6924 0 1 tie_x0
xfeed_6923 0 1 tie_x0
xfeed_6922 0 1 tie_x0
xfeed_6921 0 1 tie_x0
xfeed_6920 0 1 tie_x0
xfeed_3149 0 1 tie_x0
xfeed_3148 0 1 tie_x0
xfeed_3147 0 1 tie_x0
xfeed_3146 0 1 tie_x0
xfeed_3145 0 1 tie_x0
xfeed_2619 0 1 tie_x0
xfeed_2618 0 1 tie_x0
xfeed_2617 0 1 tie_x0
xfeed_2616 0 1 tie_x0
xfeed_2615 0 1 tie_x0
xfeed_2614 0 1 tie_x0
xfeed_2613 0 1 tie_x0
xfeed_2612 0 1 tie_x0
xfeed_2611 0 1 tie_x0
xfeed_2610 0 1 tie_x0
xsubckt_134_nao22_x1 0 1 147 151 156 159 nao22_x1
xfeed_3151 0 1 tie_x0
xfeed_3150 0 1 tie_x0
xfeed_7469 0 1 tie_x0
xfeed_7468 0 1 tie_x0
xfeed_7467 0 1 tie_x0
xfeed_7466 0 1 tie_x0
xfeed_7465 0 1 tie_x0
xfeed_7464 0 1 tie_x0
xfeed_7463 0 1 tie_x0
xfeed_7462 0 1 tie_x0
xfeed_7461 0 1 tie_x0
xfeed_7460 0 1 tie_x0
xfeed_6939 0 1 tie_x0
xfeed_6938 0 1 tie_x0
xfeed_6937 0 1 tie_x0
xfeed_6936 0 1 tie_x0
xfeed_6935 0 1 tie_x0
xfeed_6934 0 1 tie_x0
xfeed_6933 0 1 tie_x0
xfeed_6932 0 1 tie_x0
xfeed_6931 0 1 tie_x0
xfeed_6930 0 1 tie_x0
xfeed_3159 0 1 tie_x0
xfeed_3158 0 1 tie_x0
xfeed_3157 0 1 tie_x0
xfeed_3156 0 1 tie_x0
xfeed_3155 0 1 tie_x0
xfeed_3154 0 1 tie_x0
xfeed_3153 0 1 tie_x0
xfeed_3152 0 1 tie_x0
xfeed_2629 0 1 tie_x0
xfeed_2628 0 1 tie_x0
xfeed_2627 0 1 tie_x0
xfeed_2626 0 1 tie_x0
xfeed_2625 0 1 tie_x0
xfeed_2624 0 1 tie_x0
xfeed_2623 0 1 tie_x0
xfeed_2622 0 1 tie_x0
xfeed_2621 0 1 tie_x0
xfeed_2620 0 1 tie_x0
xfeed_609 0 1 tie_x0
xfeed_608 0 1 tie_x0
xfeed_607 0 1 tie_x0
xfeed_606 0 1 tie_x0
xfeed_605 0 1 tie_x0
xfeed_604 0 1 tie_x0
xfeed_603 0 1 tie_x0
xfeed_602 0 1 tie_x0
xfeed_601 0 1 tie_x0
xfeed_600 0 1 tie_x0
xfeed_7479 0 1 tie_x0
xfeed_7478 0 1 tie_x0
xfeed_7477 0 1 tie_x0
xfeed_7476 0 1 tie_x0
xfeed_7475 0 1 tie_x0
xfeed_7474 0 1 tie_x0
xfeed_7473 0 1 tie_x0
xfeed_7472 0 1 tie_x0
xfeed_7471 0 1 tie_x0
xfeed_7470 0 1 tie_x0
xfeed_6949 0 1 tie_x0
xfeed_6948 0 1 tie_x0
xfeed_6947 0 1 tie_x0
xfeed_6946 0 1 tie_x0
xfeed_6945 0 1 tie_x0
xfeed_6944 0 1 tie_x0
xfeed_6943 0 1 tie_x0
xfeed_6942 0 1 tie_x0
xfeed_6941 0 1 rowend_x0
xfeed_6940 0 1 tie_x0
xfeed_3169 0 1 tie_x0
xfeed_3168 0 1 tie_x0
xfeed_3167 0 1 tie_x0
xfeed_3166 0 1 tie_x0
xfeed_3165 0 1 tie_x0
xfeed_3164 0 1 tie_x0
xfeed_3163 0 1 tie_x0
xfeed_3162 0 1 tie_x0
xfeed_3161 0 1 tie_x0
xfeed_3160 0 1 tie_x0
xfeed_2639 0 1 tie_x0
xfeed_2638 0 1 tie_x0
xfeed_2637 0 1 tie_x0
xfeed_2636 0 1 tie_x0
xfeed_2635 0 1 tie_x0
xfeed_2634 0 1 tie_x0
xfeed_2633 0 1 tie_x0
xfeed_2632 0 1 tie_x0
xfeed_2631 0 1 tie_x0
xfeed_2630 0 1 tie_x0
xfeed_619 0 1 tie_x0
xfeed_618 0 1 tie_x0
xfeed_617 0 1 tie_x0
xfeed_616 0 1 tie_x0
xfeed_615 0 1 tie_x0
xfeed_614 0 1 tie_x0
xfeed_613 0 1 tie_x0
xfeed_612 0 1 tie_x0
xfeed_611 0 1 tie_x0
xfeed_610 0 1 tie_x0
xfeed_7489 0 1 tie_x0
xfeed_7488 0 1 tie_x0
xfeed_7487 0 1 tie_x0
xfeed_7486 0 1 tie_x0
xfeed_7485 0 1 tie_x0
xfeed_7484 0 1 tie_x0
xfeed_7483 0 1 tie_x0
xfeed_7482 0 1 tie_x0
xfeed_7481 0 1 tie_x0
xfeed_7480 0 1 tie_x0
xfeed_6959 0 1 tie_x0
xfeed_6958 0 1 tie_x0
xfeed_6957 0 1 tie_x0
xfeed_6956 0 1 tie_x0
xfeed_6955 0 1 tie_x0
xfeed_6954 0 1 tie_x0
xfeed_6953 0 1 tie_x0
xfeed_6952 0 1 tie_x0
xfeed_6951 0 1 tie_x0
xfeed_6950 0 1 tie_x0
xfeed_3179 0 1 tie_x0
xfeed_3178 0 1 tie_x0
xfeed_3177 0 1 tie_x0
xfeed_3176 0 1 tie_x0
xfeed_3175 0 1 tie_x0
xfeed_3174 0 1 tie_x0
xfeed_3173 0 1 tie_x0
xfeed_3172 0 1 tie_x0
xfeed_3171 0 1 tie_x0
xfeed_3170 0 1 tie_x0
xfeed_2649 0 1 tie_x0
xfeed_2648 0 1 tie_x0
xfeed_2647 0 1 tie_x0
xfeed_2646 0 1 tie_x0
xfeed_2645 0 1 tie_x0
xfeed_2644 0 1 tie_x0
xfeed_2643 0 1 tie_x0
xfeed_2642 0 1 tie_x0
xfeed_2641 0 1 tie_x0
xfeed_2640 0 1 tie_x0
xfeed_629 0 1 tie_x0
xfeed_628 0 1 tie_x0
xfeed_627 0 1 tie_x0
xfeed_626 0 1 tie_x0
xfeed_625 0 1 tie_x0
xfeed_624 0 1 tie_x0
xfeed_623 0 1 tie_x0
xfeed_622 0 1 tie_x0
xfeed_621 0 1 tie_x0
xfeed_620 0 1 tie_x0
xfeed_8109 0 1 tie_x0
xfeed_8108 0 1 tie_x0
xfeed_8107 0 1 tie_x0
xfeed_8106 0 1 tie_x0
xfeed_8105 0 1 tie_x0
xfeed_8104 0 1 tie_x0
xfeed_8103 0 1 tie_x0
xfeed_8102 0 1 tie_x0
xfeed_8101 0 1 tie_x0
xfeed_8100 0 1 tie_x0
xfeed_7499 0 1 tie_x0
xfeed_7498 0 1 tie_x0
xfeed_7497 0 1 tie_x0
xfeed_7496 0 1 tie_x0
xfeed_7495 0 1 tie_x0
xfeed_7494 0 1 tie_x0
xfeed_7493 0 1 tie_x0
xfeed_7492 0 1 tie_x0
xfeed_7491 0 1 tie_x0
xfeed_7490 0 1 tie_x0
xfeed_6969 0 1 tie_x0
xfeed_6968 0 1 tie_x0
xfeed_6967 0 1 tie_x0
xfeed_6966 0 1 tie_x0
xfeed_6965 0 1 tie_x0
xfeed_6964 0 1 tie_x0
xfeed_6963 0 1 tie_x0
xfeed_6962 0 1 tie_x0
xfeed_6961 0 1 tie_x0
xfeed_6960 0 1 tie_x0
xfeed_3189 0 1 tie_x0
xfeed_3188 0 1 tie_x0
xfeed_3187 0 1 tie_x0
xfeed_3186 0 1 tie_x0
xfeed_3185 0 1 tie_x0
xfeed_3184 0 1 tie_x0
xfeed_3183 0 1 tie_x0
xfeed_3182 0 1 tie_x0
xfeed_3181 0 1 tie_x0
xfeed_3180 0 1 tie_x0
xfeed_2659 0 1 tie_x0
xfeed_2658 0 1 tie_x0
xfeed_2657 0 1 tie_x0
xfeed_2656 0 1 tie_x0
xfeed_2655 0 1 tie_x0
xfeed_2654 0 1 tie_x0
xfeed_2653 0 1 tie_x0
xfeed_2652 0 1 tie_x0
xfeed_2651 0 1 tie_x0
xfeed_2650 0 1 tie_x0
xfeed_639 0 1 tie_x0
xfeed_638 0 1 tie_x0
xfeed_637 0 1 tie_x0
xfeed_636 0 1 tie_x0
xfeed_635 0 1 tie_x0
xfeed_634 0 1 tie_x0
xfeed_633 0 1 tie_x0
xfeed_632 0 1 tie_x0
xfeed_631 0 1 tie_x0
xfeed_630 0 1 tie_x0
xsubckt_80_na2_x1 0 1 192 197 193 na2_x1
xfeed_8116 0 1 tie_x0
xfeed_8115 0 1 tie_x0
xfeed_8114 0 1 tie_x0
xfeed_8113 0 1 tie_x0
xfeed_8112 0 1 tie_x0
xfeed_8111 0 1 tie_x0
xfeed_8110 0 1 tie_x0
xfeed_8119 0 1 tie_x0
xfeed_8118 0 1 tie_x0
xfeed_8117 0 1 tie_x0
xfeed_6979 0 1 tie_x0
xfeed_6978 0 1 tie_x0
xfeed_6977 0 1 tie_x0
xfeed_6976 0 1 tie_x0
xfeed_6975 0 1 tie_x0
xfeed_6974 0 1 tie_x0
xfeed_6973 0 1 tie_x0
xfeed_6972 0 1 tie_x0
xfeed_6971 0 1 tie_x0
xfeed_6970 0 1 tie_x0
xfeed_3199 0 1 tie_x0
xfeed_3198 0 1 tie_x0
xfeed_3197 0 1 tie_x0
xfeed_3196 0 1 tie_x0
xfeed_3195 0 1 tie_x0
xfeed_3194 0 1 tie_x0
xfeed_3193 0 1 tie_x0
xfeed_3192 0 1 tie_x0
xfeed_3191 0 1 tie_x0
xfeed_3190 0 1 tie_x0
xfeed_2669 0 1 tie_x0
xfeed_2668 0 1 tie_x0
xfeed_2667 0 1 tie_x0
xfeed_2666 0 1 tie_x0
xfeed_2665 0 1 rowend_x0
xfeed_2664 0 1 tie_x0
xfeed_2663 0 1 tie_x0
xfeed_2662 0 1 tie_x0
xfeed_2661 0 1 tie_x0
xfeed_2660 0 1 tie_x0
xfeed_646 0 1 tie_x0
xfeed_645 0 1 tie_x0
xfeed_644 0 1 tie_x0
xfeed_643 0 1 tie_x0
xfeed_642 0 1 tie_x0
xfeed_641 0 1 tie_x0
xfeed_640 0 1 tie_x0
xsubckt_62_nxr2_x1 0 1 209 82 212 nxr2_x1
xfeed_8123 0 1 tie_x0
xfeed_8122 0 1 tie_x0
xfeed_8121 0 1 tie_x0
xfeed_8120 0 1 tie_x0
xfeed_649 0 1 tie_x0
xfeed_648 0 1 tie_x0
xfeed_647 0 1 tie_x0
xsubckt_141_na3_x1 0 1 140 152 147 143 na3_x1
xfeed_8129 0 1 tie_x0
xfeed_8128 0 1 tie_x0
xfeed_8127 0 1 tie_x0
xfeed_8126 0 1 tie_x0
xfeed_8125 0 1 tie_x0
xfeed_8124 0 1 tie_x0
xfeed_6989 0 1 tie_x0
xfeed_6988 0 1 tie_x0
xfeed_6987 0 1 tie_x0
xfeed_6986 0 1 tie_x0
xfeed_6985 0 1 tie_x0
xfeed_6984 0 1 tie_x0
xfeed_6983 0 1 tie_x0
xfeed_6982 0 1 tie_x0
xfeed_6981 0 1 tie_x0
xfeed_6980 0 1 tie_x0
xfeed_2679 0 1 tie_x0
xfeed_2678 0 1 tie_x0
xfeed_2677 0 1 tie_x0
xfeed_2676 0 1 tie_x0
xfeed_2675 0 1 tie_x0
xfeed_2674 0 1 tie_x0
xfeed_2673 0 1 tie_x0
xfeed_2672 0 1 tie_x0
xfeed_2671 0 1 tie_x0
xfeed_2670 0 1 tie_x0
xfeed_653 0 1 tie_x0
xfeed_652 0 1 tie_x0
xfeed_651 0 1 tie_x0
xfeed_650 0 1 tie_x0
xfeed_8130 0 1 tie_x0
xfeed_659 0 1 tie_x0
xfeed_658 0 1 tie_x0
xfeed_657 0 1 tie_x0
xfeed_656 0 1 tie_x0
xfeed_655 0 1 tie_x0
xfeed_654 0 1 tie_x0
xsubckt_46_nao22_x1 0 1 92 117 96 94 nao22_x1
xfeed_8139 0 1 tie_x0
xfeed_8138 0 1 tie_x0
xfeed_8137 0 1 tie_x0
xfeed_8136 0 1 tie_x0
xfeed_8135 0 1 tie_x0
xfeed_8134 0 1 tie_x0
xfeed_8133 0 1 tie_x0
xfeed_8132 0 1 tie_x0
xfeed_8131 0 1 tie_x0
xfeed_7609 0 1 tie_x0
xfeed_7608 0 1 tie_x0
xfeed_7607 0 1 tie_x0
xfeed_7606 0 1 tie_x0
xfeed_7605 0 1 tie_x0
xfeed_7604 0 1 tie_x0
xfeed_7603 0 1 tie_x0
xfeed_7602 0 1 tie_x0
xfeed_7601 0 1 tie_x0
xfeed_7600 0 1 tie_x0
xfeed_6999 0 1 tie_x0
xfeed_6998 0 1 tie_x0
xfeed_6997 0 1 tie_x0
xfeed_6996 0 1 tie_x0
xfeed_6995 0 1 tie_x0
xfeed_6994 0 1 tie_x0
xfeed_6993 0 1 tie_x0
xfeed_6992 0 1 tie_x0
xfeed_6991 0 1 tie_x0
xfeed_6990 0 1 tie_x0
xfeed_2689 0 1 tie_x0
xfeed_2688 0 1 tie_x0
xfeed_2687 0 1 tie_x0
xfeed_2686 0 1 tie_x0
xfeed_2685 0 1 tie_x0
xfeed_2684 0 1 tie_x0
xfeed_2683 0 1 tie_x0
xfeed_2682 0 1 tie_x0
xfeed_2681 0 1 tie_x0
xfeed_2680 0 1 tie_x0
xfeed_660 0 1 tie_x0
xfeed_669 0 1 tie_x0
xfeed_668 0 1 tie_x0
xfeed_667 0 1 tie_x0
xfeed_666 0 1 tie_x0
xfeed_665 0 1 tie_x0
xfeed_664 0 1 tie_x0
xfeed_663 0 1 tie_x0
xfeed_662 0 1 tie_x0
xfeed_661 0 1 tie_x0
xfeed_8149 0 1 tie_x0
xfeed_8148 0 1 tie_x0
xfeed_8147 0 1 tie_x0
xfeed_8146 0 1 tie_x0
xfeed_8145 0 1 tie_x0
xfeed_8144 0 1 tie_x0
xfeed_8143 0 1 tie_x0
xfeed_8142 0 1 tie_x0
xfeed_8141 0 1 tie_x0
xfeed_8140 0 1 tie_x0
xfeed_7619 0 1 tie_x0
xfeed_7618 0 1 tie_x0
xfeed_7617 0 1 tie_x0
xfeed_7616 0 1 tie_x0
xfeed_7615 0 1 tie_x0
xfeed_7614 0 1 tie_x0
xfeed_7613 0 1 tie_x0
xfeed_7612 0 1 tie_x0
xfeed_7611 0 1 tie_x0
xfeed_7610 0 1 tie_x0
xfeed_3309 0 1 tie_x0
xfeed_3308 0 1 tie_x0
xfeed_3307 0 1 tie_x0
xfeed_3306 0 1 tie_x0
xfeed_3305 0 1 tie_x0
xfeed_3304 0 1 tie_x0
xfeed_3303 0 1 tie_x0
xfeed_3302 0 1 tie_x0
xfeed_3301 0 1 tie_x0
xfeed_3300 0 1 tie_x0
xfeed_2699 0 1 tie_x0
xfeed_2698 0 1 tie_x0
xfeed_2697 0 1 tie_x0
xfeed_2696 0 1 tie_x0
xfeed_2695 0 1 tie_x0
xfeed_2694 0 1 tie_x0
xfeed_2693 0 1 tie_x0
xfeed_2692 0 1 tie_x0
xfeed_2691 0 1 tie_x0
xfeed_2690 0 1 tie_x0
xfeed_679 0 1 tie_x0
xfeed_678 0 1 tie_x0
xfeed_677 0 1 tie_x0
xfeed_676 0 1 tie_x0
xfeed_675 0 1 tie_x0
xfeed_674 0 1 tie_x0
xfeed_673 0 1 tie_x0
xfeed_672 0 1 tie_x0
xfeed_671 0 1 tie_x0
xfeed_670 0 1 tie_x0
xsubckt_34_ao22_x2 0 1 104 107 110 112 ao22_x2
xfeed_8159 0 1 tie_x0
xfeed_8158 0 1 tie_x0
xfeed_8157 0 1 tie_x0
xfeed_8156 0 1 tie_x0
xfeed_8155 0 1 tie_x0
xfeed_8154 0 1 tie_x0
xfeed_8153 0 1 tie_x0
xfeed_8152 0 1 tie_x0
xfeed_8151 0 1 tie_x0
xfeed_8150 0 1 tie_x0
xfeed_7629 0 1 tie_x0
xfeed_7628 0 1 tie_x0
xfeed_7627 0 1 tie_x0
xfeed_7626 0 1 tie_x0
xfeed_7625 0 1 tie_x0
xfeed_7624 0 1 tie_x0
xfeed_7623 0 1 tie_x0
xfeed_7622 0 1 tie_x0
xfeed_7621 0 1 tie_x0
xfeed_7620 0 1 tie_x0
xfeed_3319 0 1 tie_x0
xfeed_3318 0 1 tie_x0
xfeed_3317 0 1 tie_x0
xfeed_3316 0 1 tie_x0
xfeed_3315 0 1 tie_x0
xfeed_3314 0 1 tie_x0
xfeed_3313 0 1 tie_x0
xfeed_3312 0 1 rowend_x0
xfeed_3311 0 1 tie_x0
xfeed_3310 0 1 tie_x0
xsubckt_123_ao22_x2 0 1 156 157 162 166 ao22_x2
xfeed_689 0 1 tie_x0
xfeed_688 0 1 tie_x0
xfeed_687 0 1 tie_x0
xfeed_686 0 1 tie_x0
xfeed_685 0 1 tie_x0
xfeed_684 0 1 tie_x0
xfeed_683 0 1 tie_x0
xfeed_682 0 1 tie_x0
xfeed_681 0 1 tie_x0
xfeed_680 0 1 tie_x0
xfeed_8169 0 1 tie_x0
xfeed_8168 0 1 tie_x0
xfeed_8167 0 1 tie_x0
xfeed_8166 0 1 tie_x0
xfeed_8165 0 1 tie_x0
xfeed_8164 0 1 tie_x0
xfeed_8163 0 1 tie_x0
xfeed_8162 0 1 tie_x0
xfeed_8161 0 1 tie_x0
xfeed_8160 0 1 tie_x0
xfeed_7639 0 1 tie_x0
xfeed_7638 0 1 tie_x0
xfeed_7637 0 1 tie_x0
xfeed_7636 0 1 tie_x0
xfeed_7635 0 1 tie_x0
xfeed_7634 0 1 tie_x0
xfeed_7633 0 1 tie_x0
xfeed_7632 0 1 tie_x0
xfeed_7631 0 1 tie_x0
xfeed_7630 0 1 tie_x0
xfeed_3329 0 1 tie_x0
xfeed_3328 0 1 tie_x0
xfeed_3327 0 1 tie_x0
xfeed_3326 0 1 tie_x0
xfeed_3325 0 1 tie_x0
xfeed_3324 0 1 tie_x0
xfeed_3323 0 1 tie_x0
xfeed_3322 0 1 tie_x0
xfeed_3321 0 1 tie_x0
xfeed_3320 0 1 tie_x0
xfeed_699 0 1 tie_x0
xfeed_698 0 1 tie_x0
xfeed_697 0 1 tie_x0
xfeed_696 0 1 tie_x0
xfeed_695 0 1 tie_x0
xfeed_694 0 1 tie_x0
xfeed_693 0 1 tie_x0
xfeed_692 0 1 tie_x0
xfeed_691 0 1 tie_x0
xfeed_690 0 1 tie_x0
xsubckt_129_o2_x2 0 1 151 76 5 o2_x2
xfeed_8179 0 1 tie_x0
xfeed_8178 0 1 tie_x0
xfeed_8177 0 1 tie_x0
xfeed_8176 0 1 tie_x0
xfeed_8175 0 1 tie_x0
xfeed_8174 0 1 tie_x0
xfeed_8173 0 1 tie_x0
xfeed_8172 0 1 tie_x0
xfeed_8171 0 1 tie_x0
xfeed_8170 0 1 tie_x0
xfeed_7649 0 1 tie_x0
xfeed_7648 0 1 tie_x0
xfeed_7647 0 1 tie_x0
xfeed_7646 0 1 tie_x0
xfeed_7645 0 1 tie_x0
xfeed_7644 0 1 tie_x0
xfeed_7643 0 1 tie_x0
xfeed_7642 0 1 tie_x0
xfeed_7641 0 1 tie_x0
xfeed_7640 0 1 tie_x0
xfeed_3339 0 1 tie_x0
xfeed_3338 0 1 tie_x0
xfeed_3337 0 1 tie_x0
xfeed_3336 0 1 tie_x0
xfeed_3335 0 1 tie_x0
xfeed_3334 0 1 tie_x0
xfeed_3333 0 1 tie_x0
xfeed_3332 0 1 tie_x0
xfeed_3331 0 1 rowend_x0
xfeed_3330 0 1 tie_x0
xfeed_2809 0 1 tie_x0
xfeed_2808 0 1 tie_x0
xfeed_2807 0 1 tie_x0
xfeed_2806 0 1 tie_x0
xfeed_2805 0 1 tie_x0
xfeed_2804 0 1 tie_x0
xfeed_2803 0 1 tie_x0
xfeed_2802 0 1 tie_x0
xfeed_2801 0 1 tie_x0
xfeed_2800 0 1 tie_x0
xfeed_8189 0 1 tie_x0
xfeed_8188 0 1 tie_x0
xfeed_8187 0 1 tie_x0
xfeed_8186 0 1 tie_x0
xfeed_8185 0 1 tie_x0
xfeed_8184 0 1 tie_x0
xfeed_8183 0 1 rowend_x0
xfeed_8182 0 1 tie_x0
xfeed_8181 0 1 tie_x0
xfeed_8180 0 1 tie_x0
xfeed_7659 0 1 tie_x0
xfeed_7658 0 1 tie_x0
xfeed_7657 0 1 tie_x0
xfeed_7656 0 1 tie_x0
xfeed_7655 0 1 tie_x0
xfeed_7654 0 1 tie_x0
xfeed_7653 0 1 tie_x0
xfeed_7652 0 1 tie_x0
xfeed_7651 0 1 tie_x0
xfeed_7650 0 1 tie_x0
xfeed_3349 0 1 tie_x0
xfeed_3348 0 1 tie_x0
xfeed_3347 0 1 tie_x0
xfeed_3346 0 1 tie_x0
xfeed_3345 0 1 tie_x0
xfeed_3344 0 1 tie_x0
xfeed_3343 0 1 tie_x0
xfeed_3342 0 1 tie_x0
xfeed_3341 0 1 tie_x0
xfeed_3340 0 1 tie_x0
xfeed_2819 0 1 tie_x0
xfeed_2818 0 1 tie_x0
xfeed_2817 0 1 tie_x0
xfeed_2816 0 1 tie_x0
xfeed_2815 0 1 tie_x0
xfeed_2814 0 1 tie_x0
xfeed_2813 0 1 tie_x0
xfeed_2812 0 1 tie_x0
xfeed_2811 0 1 rowend_x0
xfeed_2810 0 1 tie_x0
xfeed_8199 0 1 tie_x0
xfeed_8198 0 1 tie_x0
xfeed_8197 0 1 tie_x0
xfeed_8196 0 1 tie_x0
xfeed_8195 0 1 tie_x0
xfeed_8194 0 1 tie_x0
xfeed_8193 0 1 tie_x0
xfeed_8192 0 1 tie_x0
xfeed_8191 0 1 tie_x0
xfeed_8190 0 1 tie_x0
xfeed_7669 0 1 tie_x0
xfeed_7668 0 1 tie_x0
xfeed_7667 0 1 tie_x0
xfeed_7666 0 1 tie_x0
xfeed_7665 0 1 tie_x0
xfeed_7664 0 1 tie_x0
xfeed_7663 0 1 tie_x0
xfeed_7662 0 1 tie_x0
xfeed_7661 0 1 tie_x0
xfeed_7660 0 1 tie_x0
xfeed_3359 0 1 tie_x0
xfeed_3358 0 1 tie_x0
xfeed_3357 0 1 tie_x0
xfeed_3356 0 1 rowend_x0
xfeed_3355 0 1 tie_x0
xfeed_3354 0 1 tie_x0
xfeed_3353 0 1 tie_x0
xfeed_3352 0 1 tie_x0
xfeed_3351 0 1 tie_x0
xfeed_3350 0 1 tie_x0
xfeed_2829 0 1 tie_x0
xfeed_2828 0 1 tie_x0
xfeed_2827 0 1 tie_x0
xfeed_2826 0 1 tie_x0
xfeed_2825 0 1 tie_x0
xfeed_2824 0 1 tie_x0
xfeed_2823 0 1 tie_x0
xfeed_2822 0 1 tie_x0
xfeed_2821 0 1 tie_x0
xfeed_2820 0 1 tie_x0
xfeed_800 0 1 rowend_x0
xfeed_809 0 1 tie_x0
xfeed_808 0 1 tie_x0
xfeed_807 0 1 tie_x0
xfeed_806 0 1 tie_x0
xfeed_805 0 1 tie_x0
xfeed_804 0 1 tie_x0
xfeed_803 0 1 tie_x0
xfeed_802 0 1 tie_x0
xfeed_801 0 1 tie_x0
xfeed_7679 0 1 tie_x0
xfeed_7678 0 1 tie_x0
xfeed_7677 0 1 tie_x0
xfeed_7676 0 1 tie_x0
xfeed_7675 0 1 tie_x0
xfeed_7674 0 1 tie_x0
xfeed_7673 0 1 tie_x0
xfeed_7672 0 1 tie_x0
xfeed_7671 0 1 tie_x0
xfeed_7670 0 1 tie_x0
xfeed_3369 0 1 tie_x0
xfeed_3368 0 1 tie_x0
xfeed_3367 0 1 tie_x0
xfeed_3366 0 1 tie_x0
xfeed_3365 0 1 tie_x0
xfeed_3364 0 1 tie_x0
xfeed_3363 0 1 tie_x0
xfeed_3362 0 1 tie_x0
xfeed_3361 0 1 tie_x0
xfeed_3360 0 1 tie_x0
xfeed_2839 0 1 tie_x0
xfeed_2838 0 1 tie_x0
xfeed_2837 0 1 tie_x0
xfeed_2836 0 1 tie_x0
xfeed_2835 0 1 tie_x0
xfeed_2834 0 1 tie_x0
xfeed_2833 0 1 tie_x0
xfeed_2832 0 1 tie_x0
xfeed_2831 0 1 tie_x0
xfeed_2830 0 1 tie_x0
xsubckt_146_a3_x2 0 1 136 145 141 139 a3_x2
xfeed_819 0 1 tie_x0
xfeed_818 0 1 tie_x0
xfeed_817 0 1 tie_x0
xfeed_816 0 1 tie_x0
xfeed_815 0 1 tie_x0
xfeed_814 0 1 tie_x0
xfeed_813 0 1 tie_x0
xfeed_812 0 1 tie_x0
xfeed_811 0 1 tie_x0
xfeed_810 0 1 tie_x0
xsubckt_104_ao22_x2 0 1 173 177 176 179 ao22_x2
xfeed_7689 0 1 tie_x0
xfeed_7688 0 1 tie_x0
xfeed_7687 0 1 tie_x0
xfeed_7686 0 1 tie_x0
xfeed_7685 0 1 tie_x0
xfeed_7684 0 1 tie_x0
xfeed_7683 0 1 tie_x0
xfeed_7682 0 1 tie_x0
xfeed_7681 0 1 tie_x0
xfeed_7680 0 1 tie_x0
xfeed_3379 0 1 tie_x0
xfeed_3378 0 1 tie_x0
xfeed_3377 0 1 tie_x0
xfeed_3376 0 1 tie_x0
xfeed_3375 0 1 tie_x0
xfeed_3374 0 1 tie_x0
xfeed_3373 0 1 tie_x0
xfeed_3372 0 1 tie_x0
xfeed_3371 0 1 tie_x0
xfeed_3370 0 1 tie_x0
xfeed_2849 0 1 tie_x0
xfeed_2848 0 1 tie_x0
xfeed_2847 0 1 tie_x0
xfeed_2846 0 1 tie_x0
xfeed_2845 0 1 tie_x0
xfeed_2844 0 1 tie_x0
xfeed_2843 0 1 tie_x0
xfeed_2842 0 1 tie_x0
xfeed_2841 0 1 tie_x0
xfeed_2840 0 1 tie_x0
xfeed_824 0 1 tie_x0
xfeed_823 0 1 tie_x0
xfeed_822 0 1 tie_x0
xfeed_821 0 1 tie_x0
xfeed_820 0 1 tie_x0
xsubckt_161_sff1_x4 0 1 76 216 66 sff1_x4
xfeed_825 0 1 tie_x0
xfeed_826 0 1 tie_x0
xfeed_827 0 1 tie_x0
xfeed_828 0 1 tie_x0
xfeed_829 0 1 tie_x0
xfeed_8309 0 1 tie_x0
xfeed_8308 0 1 tie_x0
xfeed_8307 0 1 tie_x0
xfeed_8306 0 1 tie_x0
xfeed_8305 0 1 tie_x0
xfeed_8304 0 1 tie_x0
xfeed_8303 0 1 tie_x0
xfeed_8302 0 1 tie_x0
xfeed_8301 0 1 tie_x0
xfeed_8300 0 1 tie_x0
xfeed_7699 0 1 tie_x0
xfeed_7698 0 1 tie_x0
xfeed_7697 0 1 tie_x0
xfeed_7696 0 1 tie_x0
xfeed_7695 0 1 tie_x0
xfeed_7694 0 1 tie_x0
xfeed_7693 0 1 tie_x0
xfeed_7692 0 1 tie_x0
xfeed_7691 0 1 tie_x0
xfeed_7690 0 1 tie_x0
xfeed_3389 0 1 tie_x0
xfeed_3388 0 1 tie_x0
xfeed_3387 0 1 tie_x0
xfeed_3386 0 1 tie_x0
xfeed_3385 0 1 tie_x0
xfeed_3384 0 1 tie_x0
xfeed_3383 0 1 tie_x0
xfeed_3382 0 1 tie_x0
xfeed_3381 0 1 tie_x0
xfeed_3380 0 1 tie_x0
xfeed_2859 0 1 tie_x0
xfeed_2858 0 1 tie_x0
xfeed_2857 0 1 tie_x0
xfeed_2856 0 1 tie_x0
xfeed_2855 0 1 tie_x0
xfeed_2854 0 1 tie_x0
xfeed_2853 0 1 tie_x0
xfeed_2852 0 1 tie_x0
xfeed_2851 0 1 tie_x0
xfeed_2850 0 1 tie_x0
xsubckt_99_na2_x1 0 1 177 80 9 na2_x1
xsubckt_157_sff1_x4 0 1 80 220 34 sff1_x4
xfeed_830 0 1 tie_x0
xfeed_831 0 1 tie_x0
xfeed_832 0 1 tie_x0
xfeed_833 0 1 tie_x0
xfeed_834 0 1 tie_x0
xfeed_835 0 1 tie_x0
xfeed_836 0 1 tie_x0
xfeed_837 0 1 tie_x0
xfeed_838 0 1 tie_x0
xfeed_839 0 1 tie_x0
xfeed_8319 0 1 tie_x0
xfeed_8318 0 1 tie_x0
xfeed_8317 0 1 tie_x0
xfeed_8316 0 1 tie_x0
xfeed_8315 0 1 tie_x0
xfeed_8314 0 1 rowend_x0
xfeed_8313 0 1 tie_x0
xfeed_8312 0 1 tie_x0
xfeed_8311 0 1 tie_x0
xfeed_8310 0 1 tie_x0
xfeed_4009 0 1 tie_x0
xfeed_4008 0 1 tie_x0
xfeed_4007 0 1 tie_x0
xfeed_4006 0 1 tie_x0
xfeed_4005 0 1 rowend_x0
xfeed_4004 0 1 tie_x0
xfeed_4003 0 1 tie_x0
xfeed_4002 0 1 tie_x0
xfeed_4001 0 1 tie_x0
xfeed_4000 0 1 tie_x0
xfeed_3399 0 1 tie_x0
xfeed_3398 0 1 tie_x0
xfeed_3397 0 1 tie_x0
xfeed_3396 0 1 tie_x0
xfeed_3395 0 1 tie_x0
xfeed_3394 0 1 tie_x0
xfeed_3393 0 1 tie_x0
xfeed_3392 0 1 tie_x0
xfeed_3391 0 1 tie_x0
xfeed_3390 0 1 tie_x0
xfeed_2869 0 1 tie_x0
xfeed_2868 0 1 tie_x0
xfeed_2867 0 1 tie_x0
xfeed_2866 0 1 tie_x0
xfeed_2865 0 1 tie_x0
xfeed_2864 0 1 tie_x0
xfeed_2863 0 1 tie_x0
xfeed_2862 0 1 tie_x0
xfeed_2861 0 1 tie_x0
xfeed_2860 0 1 tie_x0
xsubckt_109_nxr2_x1 0 1 168 173 170 nxr2_x1
xfeed_840 0 1 tie_x0
xfeed_841 0 1 tie_x0
xfeed_842 0 1 tie_x0
xfeed_843 0 1 tie_x0
xfeed_844 0 1 tie_x0
xfeed_845 0 1 tie_x0
xfeed_846 0 1 tie_x0
xfeed_847 0 1 tie_x0
xfeed_848 0 1 tie_x0
xfeed_849 0 1 tie_x0
xfeed_8329 0 1 tie_x0
xfeed_8328 0 1 tie_x0
xfeed_8327 0 1 tie_x0
xfeed_8326 0 1 tie_x0
xfeed_8325 0 1 tie_x0
xfeed_8324 0 1 tie_x0
xfeed_8323 0 1 tie_x0
xfeed_8322 0 1 tie_x0
xfeed_8321 0 1 tie_x0
xfeed_8320 0 1 tie_x0
xfeed_4019 0 1 tie_x0
xfeed_4018 0 1 tie_x0
xfeed_4017 0 1 tie_x0
xfeed_4016 0 1 tie_x0
xfeed_4015 0 1 tie_x0
xfeed_4014 0 1 tie_x0
xfeed_4013 0 1 tie_x0
xfeed_4012 0 1 tie_x0
xfeed_4011 0 1 tie_x0
xfeed_4010 0 1 tie_x0
xfeed_2879 0 1 tie_x0
xfeed_2878 0 1 tie_x0
xfeed_2877 0 1 tie_x0
xfeed_2876 0 1 tie_x0
xfeed_2875 0 1 tie_x0
xfeed_2874 0 1 tie_x0
xfeed_2873 0 1 tie_x0
xfeed_2872 0 1 tie_x0
xfeed_2871 0 1 tie_x0
xfeed_2870 0 1 tie_x0
xfeed_850 0 1 tie_x0
xfeed_851 0 1 tie_x0
xfeed_852 0 1 tie_x0
xfeed_853 0 1 tie_x0
xfeed_854 0 1 tie_x0
xfeed_855 0 1 tie_x0
xfeed_856 0 1 tie_x0
xfeed_857 0 1 tie_x0
xfeed_858 0 1 tie_x0
xfeed_859 0 1 tie_x0
xfeed_8339 0 1 tie_x0
xfeed_8338 0 1 rowend_x0
xfeed_8337 0 1 tie_x0
xfeed_8336 0 1 tie_x0
xfeed_8335 0 1 tie_x0
xfeed_8334 0 1 tie_x0
xfeed_8333 0 1 tie_x0
xfeed_8332 0 1 tie_x0
xfeed_8331 0 1 tie_x0
xfeed_8330 0 1 tie_x0
xfeed_7809 0 1 tie_x0
xfeed_7808 0 1 tie_x0
xfeed_7807 0 1 tie_x0
xfeed_7806 0 1 tie_x0
xfeed_7805 0 1 tie_x0
xfeed_7804 0 1 tie_x0
xfeed_7803 0 1 tie_x0
xfeed_7802 0 1 tie_x0
xfeed_7801 0 1 tie_x0
xfeed_7800 0 1 tie_x0
xfeed_4029 0 1 tie_x0
xfeed_4028 0 1 tie_x0
xfeed_4027 0 1 tie_x0
xfeed_4026 0 1 tie_x0
xfeed_4025 0 1 tie_x0
xfeed_4024 0 1 tie_x0
xfeed_4023 0 1 tie_x0
xfeed_4022 0 1 tie_x0
xfeed_4021 0 1 tie_x0
xfeed_4020 0 1 tie_x0
xfeed_2889 0 1 tie_x0
xfeed_2888 0 1 tie_x0
xfeed_2887 0 1 tie_x0
xfeed_2886 0 1 tie_x0
xfeed_2885 0 1 tie_x0
xfeed_2884 0 1 tie_x0
xfeed_2883 0 1 tie_x0
xfeed_2882 0 1 tie_x0
xfeed_2881 0 1 tie_x0
xfeed_2880 0 1 tie_x0
xsubckt_74_ao22_x2 0 1 198 208 207 85 ao22_x2
xsubckt_112_a2_x2 0 1 166 78 7 a2_x2
xfeed_860 0 1 tie_x0
xfeed_861 0 1 tie_x0
xfeed_862 0 1 tie_x0
xfeed_863 0 1 tie_x0
xfeed_864 0 1 tie_x0
xfeed_865 0 1 tie_x0
xfeed_866 0 1 tie_x0
xfeed_867 0 1 tie_x0
xfeed_868 0 1 tie_x0
xfeed_869 0 1 tie_x0
xfeed_8349 0 1 tie_x0
xfeed_8348 0 1 tie_x0
xfeed_8347 0 1 tie_x0
xfeed_8346 0 1 tie_x0
xfeed_8345 0 1 tie_x0
xfeed_8344 0 1 tie_x0
xfeed_8343 0 1 tie_x0
xfeed_8342 0 1 tie_x0
xfeed_8341 0 1 tie_x0
xfeed_8340 0 1 tie_x0
xfeed_7819 0 1 tie_x0
xfeed_7818 0 1 tie_x0
xfeed_7817 0 1 tie_x0
xfeed_7816 0 1 tie_x0
xfeed_7815 0 1 tie_x0
xfeed_7814 0 1 tie_x0
xfeed_7813 0 1 tie_x0
xfeed_7812 0 1 tie_x0
xfeed_7811 0 1 tie_x0
xfeed_7810 0 1 tie_x0
xfeed_4039 0 1 tie_x0
xfeed_4038 0 1 tie_x0
xfeed_4037 0 1 tie_x0
xfeed_4036 0 1 tie_x0
xfeed_4035 0 1 tie_x0
xfeed_4034 0 1 tie_x0
xfeed_4033 0 1 tie_x0
xfeed_4032 0 1 tie_x0
xfeed_4031 0 1 tie_x0
xfeed_4030 0 1 tie_x0
xfeed_3509 0 1 tie_x0
xfeed_3508 0 1 tie_x0
xfeed_3507 0 1 tie_x0
xfeed_3506 0 1 tie_x0
xfeed_3505 0 1 tie_x0
xfeed_3504 0 1 tie_x0
xfeed_3503 0 1 tie_x0
xfeed_3502 0 1 tie_x0
xfeed_3501 0 1 tie_x0
xfeed_3500 0 1 tie_x0
xfeed_2899 0 1 tie_x0
xfeed_2898 0 1 tie_x0
xfeed_2897 0 1 rowend_x0
xfeed_2896 0 1 tie_x0
xfeed_2895 0 1 tie_x0
xfeed_2894 0 1 tie_x0
xfeed_2893 0 1 tie_x0
xfeed_2892 0 1 tie_x0
xfeed_2891 0 1 tie_x0
xfeed_2890 0 1 tie_x0
xsubckt_132_a2_x2 0 1 216 131 149 a2_x2
xsubckt_28_a4_x2 0 1 110 18 17 12 11 a4_x2
xfeed_870 0 1 tie_x0
xfeed_871 0 1 tie_x0
xfeed_872 0 1 tie_x0
xfeed_873 0 1 tie_x0
xfeed_874 0 1 tie_x0
xfeed_875 0 1 tie_x0
xfeed_876 0 1 tie_x0
xfeed_877 0 1 tie_x0
xfeed_878 0 1 tie_x0
xfeed_879 0 1 tie_x0
xfeed_8359 0 1 tie_x0
xfeed_8358 0 1 tie_x0
xfeed_8357 0 1 tie_x0
xfeed_8356 0 1 tie_x0
xfeed_8355 0 1 tie_x0
xfeed_8354 0 1 tie_x0
xfeed_8353 0 1 tie_x0
xfeed_8352 0 1 tie_x0
xfeed_8351 0 1 tie_x0
xfeed_8350 0 1 tie_x0
xfeed_7829 0 1 tie_x0
xfeed_7828 0 1 tie_x0
xfeed_7827 0 1 tie_x0
xfeed_7826 0 1 tie_x0
xfeed_7825 0 1 tie_x0
xfeed_7824 0 1 tie_x0
xfeed_7823 0 1 tie_x0
xfeed_7822 0 1 tie_x0
xfeed_7821 0 1 tie_x0
xfeed_7820 0 1 tie_x0
xfeed_4049 0 1 tie_x0
xfeed_4048 0 1 tie_x0
xfeed_4047 0 1 tie_x0
xfeed_4046 0 1 tie_x0
xfeed_4045 0 1 tie_x0
xfeed_4044 0 1 tie_x0
xfeed_4043 0 1 tie_x0
xfeed_4042 0 1 tie_x0
xfeed_4041 0 1 tie_x0
xfeed_4040 0 1 tie_x0
xfeed_3519 0 1 tie_x0
xfeed_3518 0 1 tie_x0
xfeed_3517 0 1 tie_x0
xfeed_3516 0 1 tie_x0
xfeed_3515 0 1 tie_x0
xfeed_3514 0 1 tie_x0
xfeed_3513 0 1 tie_x0
xfeed_3512 0 1 tie_x0
xfeed_3511 0 1 tie_x0
xfeed_3510 0 1 tie_x0
xsubckt_83_nxr2_x1 0 1 189 199 191 nxr2_x1
xfeed_880 0 1 tie_x0
xfeed_881 0 1 tie_x0
xfeed_882 0 1 tie_x0
xfeed_883 0 1 tie_x0
xfeed_884 0 1 tie_x0
xfeed_885 0 1 tie_x0
xfeed_886 0 1 tie_x0
xfeed_887 0 1 tie_x0
xfeed_888 0 1 tie_x0
xfeed_889 0 1 tie_x0
xfeed_8369 0 1 tie_x0
xfeed_8368 0 1 tie_x0
xfeed_8367 0 1 tie_x0
xfeed_8366 0 1 rowend_x0
xfeed_8365 0 1 tie_x0
xfeed_8364 0 1 tie_x0
xfeed_8363 0 1 tie_x0
xfeed_8362 0 1 tie_x0
xfeed_8361 0 1 tie_x0
xfeed_8360 0 1 tie_x0
xfeed_7839 0 1 tie_x0
xfeed_7838 0 1 tie_x0
xfeed_7837 0 1 tie_x0
xfeed_7836 0 1 tie_x0
xfeed_7835 0 1 tie_x0
xfeed_7834 0 1 tie_x0
xfeed_7833 0 1 tie_x0
xfeed_7832 0 1 tie_x0
xfeed_7831 0 1 tie_x0
xfeed_7830 0 1 tie_x0
xfeed_4059 0 1 tie_x0
xfeed_4058 0 1 tie_x0
xfeed_4057 0 1 tie_x0
xfeed_4056 0 1 tie_x0
xfeed_4055 0 1 tie_x0
xfeed_4054 0 1 tie_x0
xfeed_4053 0 1 tie_x0
xfeed_4052 0 1 tie_x0
xfeed_4051 0 1 tie_x0
xfeed_4050 0 1 tie_x0
xfeed_3529 0 1 tie_x0
xfeed_3528 0 1 tie_x0
xfeed_3527 0 1 tie_x0
xfeed_3526 0 1 tie_x0
xfeed_3525 0 1 tie_x0
xfeed_3524 0 1 tie_x0
xfeed_3523 0 1 tie_x0
xfeed_3522 0 1 tie_x0
xfeed_3521 0 1 tie_x0
xfeed_3520 0 1 tie_x0
xsubckt_79_nxr2_x1 0 1 193 196 194 nxr2_x1
xfeed_890 0 1 tie_x0
xfeed_891 0 1 tie_x0
xfeed_892 0 1 tie_x0
xfeed_893 0 1 tie_x0
xfeed_894 0 1 tie_x0
xfeed_895 0 1 tie_x0
xfeed_896 0 1 tie_x0
xfeed_897 0 1 tie_x0
xfeed_898 0 1 tie_x0
xfeed_899 0 1 tie_x0
xfeed_8379 0 1 tie_x0
xfeed_8378 0 1 tie_x0
xfeed_8377 0 1 tie_x0
xfeed_8376 0 1 tie_x0
xfeed_8375 0 1 tie_x0
xfeed_8374 0 1 tie_x0
xfeed_8373 0 1 tie_x0
xfeed_8372 0 1 tie_x0
xfeed_8371 0 1 tie_x0
xfeed_8370 0 1 tie_x0
xfeed_7849 0 1 tie_x0
xfeed_7848 0 1 tie_x0
xfeed_7847 0 1 tie_x0
xfeed_7846 0 1 tie_x0
xfeed_7845 0 1 tie_x0
xfeed_7844 0 1 tie_x0
xfeed_7843 0 1 tie_x0
xfeed_7842 0 1 tie_x0
xfeed_7841 0 1 tie_x0
xfeed_7840 0 1 tie_x0
xfeed_4069 0 1 tie_x0
xfeed_4068 0 1 tie_x0
xfeed_4067 0 1 tie_x0
xfeed_4066 0 1 tie_x0
xfeed_4065 0 1 tie_x0
xfeed_4064 0 1 tie_x0
xfeed_4063 0 1 tie_x0
xfeed_4062 0 1 tie_x0
xfeed_4061 0 1 tie_x0
xfeed_4060 0 1 tie_x0
xfeed_3539 0 1 tie_x0
xfeed_3538 0 1 tie_x0
xfeed_3537 0 1 tie_x0
xfeed_3536 0 1 tie_x0
xfeed_3535 0 1 tie_x0
xfeed_3534 0 1 tie_x0
xfeed_3533 0 1 tie_x0
xfeed_3532 0 1 tie_x0
xfeed_3531 0 1 tie_x0
xfeed_3530 0 1 tie_x0
xsubckt_93_nao22_x1 0 1 223 181 182 183 nao22_x1
xfeed_8389 0 1 tie_x0
xfeed_8388 0 1 tie_x0
xfeed_8387 0 1 tie_x0
xfeed_8386 0 1 tie_x0
xfeed_8385 0 1 tie_x0
xfeed_8384 0 1 tie_x0
xfeed_8383 0 1 tie_x0
xfeed_8382 0 1 tie_x0
xfeed_8381 0 1 tie_x0
xfeed_8380 0 1 tie_x0
xfeed_7859 0 1 tie_x0
xfeed_7858 0 1 tie_x0
xfeed_7857 0 1 tie_x0
xfeed_7856 0 1 tie_x0
xfeed_7855 0 1 tie_x0
xfeed_7854 0 1 tie_x0
xfeed_7853 0 1 tie_x0
xfeed_7852 0 1 tie_x0
xfeed_7851 0 1 tie_x0
xfeed_7850 0 1 tie_x0
xfeed_4079 0 1 tie_x0
xfeed_4078 0 1 tie_x0
xfeed_4077 0 1 tie_x0
xfeed_4076 0 1 tie_x0
xfeed_4075 0 1 tie_x0
xfeed_4074 0 1 tie_x0
xfeed_4073 0 1 tie_x0
xfeed_4072 0 1 tie_x0
xfeed_4071 0 1 tie_x0
xfeed_4070 0 1 tie_x0
xfeed_3549 0 1 tie_x0
xfeed_3548 0 1 tie_x0
xfeed_3547 0 1 tie_x0
xfeed_3546 0 1 tie_x0
xfeed_3545 0 1 tie_x0
xfeed_3544 0 1 tie_x0
xfeed_3543 0 1 tie_x0
xfeed_3542 0 1 tie_x0
xfeed_3541 0 1 tie_x0
xfeed_3540 0 1 tie_x0
xfeed_8399 0 1 tie_x0
xfeed_8398 0 1 tie_x0
xfeed_8397 0 1 tie_x0
xfeed_8396 0 1 tie_x0
xfeed_8395 0 1 tie_x0
xfeed_8394 0 1 tie_x0
xfeed_8393 0 1 tie_x0
xfeed_8392 0 1 rowend_x0
xfeed_8391 0 1 tie_x0
xfeed_8390 0 1 tie_x0
xfeed_7869 0 1 tie_x0
xfeed_7868 0 1 tie_x0
xfeed_7867 0 1 tie_x0
xfeed_7866 0 1 tie_x0
xfeed_7865 0 1 tie_x0
xfeed_7864 0 1 tie_x0
xfeed_7863 0 1 tie_x0
xfeed_7862 0 1 tie_x0
xfeed_7861 0 1 tie_x0
xfeed_7860 0 1 tie_x0
xfeed_4089 0 1 tie_x0
xfeed_4088 0 1 tie_x0
xfeed_4087 0 1 tie_x0
xfeed_4086 0 1 tie_x0
xfeed_4085 0 1 tie_x0
xfeed_4084 0 1 tie_x0
xfeed_4083 0 1 tie_x0
xfeed_4082 0 1 tie_x0
xfeed_4081 0 1 tie_x0
xfeed_4080 0 1 tie_x0
xfeed_3559 0 1 tie_x0
xfeed_3558 0 1 tie_x0
xfeed_3557 0 1 tie_x0
xfeed_3556 0 1 tie_x0
xfeed_3555 0 1 tie_x0
xfeed_3554 0 1 tie_x0
xfeed_3553 0 1 tie_x0
xfeed_3552 0 1 tie_x0
xfeed_3551 0 1 tie_x0
xfeed_3550 0 1 tie_x0
xsubckt_55_ao22_x2 0 1 84 109 107 112 ao22_x2
xfeed_7879 0 1 tie_x0
xfeed_7878 0 1 tie_x0
xfeed_7877 0 1 tie_x0
xfeed_7876 0 1 tie_x0
xfeed_7875 0 1 tie_x0
xfeed_7874 0 1 tie_x0
xfeed_7873 0 1 tie_x0
xfeed_7872 0 1 tie_x0
xfeed_7871 0 1 tie_x0
xfeed_7870 0 1 tie_x0
xfeed_4099 0 1 tie_x0
xfeed_4098 0 1 tie_x0
xfeed_4097 0 1 tie_x0
xfeed_4096 0 1 tie_x0
xfeed_4095 0 1 tie_x0
xfeed_4094 0 1 tie_x0
xfeed_4093 0 1 tie_x0
xfeed_4092 0 1 tie_x0
xfeed_4091 0 1 tie_x0
xfeed_4090 0 1 tie_x0
xfeed_3569 0 1 tie_x0
xfeed_3568 0 1 tie_x0
xfeed_3567 0 1 tie_x0
xfeed_3566 0 1 tie_x0
xfeed_3565 0 1 tie_x0
xfeed_3564 0 1 tie_x0
xfeed_3563 0 1 tie_x0
xfeed_3562 0 1 tie_x0
xfeed_3561 0 1 tie_x0
xfeed_3560 0 1 tie_x0
xfeed_7889 0 1 tie_x0
xfeed_7888 0 1 tie_x0
xfeed_7887 0 1 tie_x0
xfeed_7886 0 1 tie_x0
xfeed_7885 0 1 tie_x0
xfeed_7884 0 1 tie_x0
xfeed_7883 0 1 tie_x0
xfeed_7882 0 1 tie_x0
xfeed_7881 0 1 tie_x0
xfeed_7880 0 1 tie_x0
xfeed_3579 0 1 tie_x0
xfeed_3578 0 1 tie_x0
xfeed_3577 0 1 tie_x0
xfeed_3576 0 1 tie_x0
xfeed_3575 0 1 tie_x0
xfeed_3574 0 1 tie_x0
xfeed_3573 0 1 tie_x0
xfeed_3572 0 1 tie_x0
xfeed_3571 0 1 tie_x0
xfeed_3570 0 1 tie_x0
xfeed_8509 0 1 tie_x0
xfeed_8508 0 1 tie_x0
xfeed_8507 0 1 tie_x0
xfeed_8506 0 1 tie_x0
xfeed_8505 0 1 tie_x0
xfeed_8504 0 1 tie_x0
xfeed_8503 0 1 tie_x0
xfeed_8502 0 1 tie_x0
xfeed_8501 0 1 tie_x0
xfeed_8500 0 1 tie_x0
xfeed_7899 0 1 tie_x0
xfeed_7898 0 1 tie_x0
xfeed_7897 0 1 tie_x0
xfeed_7896 0 1 tie_x0
xfeed_7895 0 1 tie_x0
xfeed_7894 0 1 tie_x0
xfeed_7893 0 1 tie_x0
xfeed_7892 0 1 tie_x0
xfeed_7891 0 1 tie_x0
xfeed_7890 0 1 tie_x0
xfeed_3589 0 1 tie_x0
xfeed_3588 0 1 tie_x0
xfeed_3587 0 1 tie_x0
xfeed_3586 0 1 tie_x0
xfeed_3585 0 1 tie_x0
xfeed_3584 0 1 tie_x0
xfeed_3583 0 1 tie_x0
xfeed_3582 0 1 tie_x0
xfeed_3581 0 1 tie_x0
xfeed_3580 0 1 tie_x0
xfeed_8519 0 1 tie_x0
xfeed_8518 0 1 tie_x0
xfeed_8517 0 1 tie_x0
xfeed_8516 0 1 tie_x0
xfeed_8515 0 1 tie_x0
xfeed_8514 0 1 tie_x0
xfeed_8513 0 1 tie_x0
xfeed_8512 0 1 tie_x0
xfeed_8511 0 1 tie_x0
xfeed_8510 0 1 tie_x0
xfeed_4209 0 1 rowend_x0
xfeed_4208 0 1 tie_x0
xfeed_4207 0 1 tie_x0
xfeed_4206 0 1 tie_x0
xfeed_4205 0 1 tie_x0
xfeed_4204 0 1 tie_x0
xfeed_4203 0 1 tie_x0
xfeed_4202 0 1 tie_x0
xfeed_4201 0 1 tie_x0
xfeed_4200 0 1 tie_x0
xfeed_3599 0 1 tie_x0
xfeed_3598 0 1 tie_x0
xfeed_3597 0 1 tie_x0
xfeed_3596 0 1 tie_x0
xfeed_3595 0 1 tie_x0
xfeed_3594 0 1 tie_x0
xfeed_3593 0 1 tie_x0
xfeed_3592 0 1 tie_x0
xfeed_3591 0 1 tie_x0
xfeed_3590 0 1 tie_x0
xfeed_8529 0 1 tie_x0
xfeed_8528 0 1 tie_x0
xfeed_8527 0 1 tie_x0
xfeed_8526 0 1 tie_x0
xfeed_8525 0 1 tie_x0
xfeed_8524 0 1 tie_x0
xfeed_8523 0 1 tie_x0
xfeed_8522 0 1 tie_x0
xfeed_8521 0 1 tie_x0
xfeed_8520 0 1 rowend_x0
xfeed_4219 0 1 tie_x0
xfeed_4218 0 1 tie_x0
xfeed_4217 0 1 tie_x0
xfeed_4216 0 1 tie_x0
xfeed_4215 0 1 tie_x0
xfeed_4214 0 1 tie_x0
xfeed_4213 0 1 tie_x0
xfeed_4212 0 1 tie_x0
xfeed_4211 0 1 tie_x0
xfeed_4210 0 1 tie_x0
xfeed_10 0 1 tie_x0
xfeed_11 0 1 tie_x0
xfeed_12 0 1 tie_x0
xfeed_13 0 1 tie_x0
xfeed_14 0 1 tie_x0
xfeed_15 0 1 tie_x0
xfeed_16 0 1 tie_x0
xfeed_17 0 1 tie_x0
xfeed_18 0 1 tie_x0
xfeed_19 0 1 tie_x0
xfeed_8539 0 1 tie_x0
xfeed_8538 0 1 tie_x0
xfeed_8537 0 1 tie_x0
xfeed_8536 0 1 tie_x0
xfeed_8535 0 1 tie_x0
xfeed_8534 0 1 tie_x0
xfeed_8533 0 1 tie_x0
xfeed_8532 0 1 tie_x0
xfeed_8531 0 1 tie_x0
xfeed_8530 0 1 tie_x0
xfeed_4229 0 1 tie_x0
xfeed_4228 0 1 tie_x0
xfeed_4227 0 1 tie_x0
xfeed_4226 0 1 tie_x0
xfeed_4225 0 1 tie_x0
xfeed_4224 0 1 tie_x0
xfeed_4223 0 1 tie_x0
xfeed_4222 0 1 tie_x0
xfeed_4221 0 1 tie_x0
xfeed_4220 0 1 tie_x0
xfeed_20 0 1 tie_x0
xfeed_21 0 1 tie_x0
xfeed_22 0 1 tie_x0
xfeed_23 0 1 tie_x0
xfeed_24 0 1 tie_x0
xfeed_25 0 1 tie_x0
xfeed_26 0 1 tie_x0
xfeed_27 0 1 tie_x0
xfeed_28 0 1 tie_x0
xfeed_29 0 1 tie_x0
xfeed_8549 0 1 tie_x0
xfeed_8548 0 1 tie_x0
xfeed_8547 0 1 tie_x0
xfeed_8546 0 1 tie_x0
xfeed_8545 0 1 tie_x0
xfeed_8544 0 1 tie_x0
xfeed_8543 0 1 tie_x0
xfeed_8542 0 1 tie_x0
xfeed_8541 0 1 tie_x0
xfeed_8540 0 1 tie_x0
xfeed_4239 0 1 tie_x0
xfeed_4238 0 1 tie_x0
xfeed_4237 0 1 tie_x0
xfeed_4236 0 1 tie_x0
xfeed_4235 0 1 tie_x0
xfeed_4234 0 1 tie_x0
xfeed_4233 0 1 tie_x0
xfeed_4232 0 1 tie_x0
xfeed_4231 0 1 tie_x0
xfeed_4230 0 1 tie_x0
xfeed_3709 0 1 tie_x0
xfeed_3708 0 1 tie_x0
xfeed_3707 0 1 tie_x0
xfeed_3706 0 1 tie_x0
xfeed_3705 0 1 tie_x0
xfeed_3704 0 1 tie_x0
xfeed_3703 0 1 tie_x0
xfeed_3702 0 1 tie_x0
xfeed_3701 0 1 tie_x0
xfeed_3700 0 1 tie_x0
xsubckt_40_a2_x2 0 1 98 14 15 a2_x2
xsubckt_140_nao22_x1 0 1 141 144 148 153 nao22_x1
xfeed_30 0 1 tie_x0
xfeed_31 0 1 tie_x0
xfeed_32 0 1 tie_x0
xfeed_33 0 1 tie_x0
xfeed_34 0 1 tie_x0
xfeed_35 0 1 tie_x0
xfeed_36 0 1 tie_x0
xfeed_37 0 1 tie_x0
xfeed_38 0 1 tie_x0
xfeed_39 0 1 tie_x0
xfeed_8559 0 1 tie_x0
xfeed_8558 0 1 tie_x0
xfeed_8557 0 1 tie_x0
xfeed_8556 0 1 tie_x0
xfeed_8555 0 1 tie_x0
xfeed_8554 0 1 tie_x0
xfeed_8553 0 1 tie_x0
xfeed_8552 0 1 tie_x0
xfeed_8551 0 1 tie_x0
xfeed_8550 0 1 tie_x0
xfeed_4249 0 1 tie_x0
xfeed_4248 0 1 tie_x0
xfeed_4247 0 1 tie_x0
xfeed_4246 0 1 tie_x0
xfeed_4245 0 1 tie_x0
xfeed_4244 0 1 tie_x0
xfeed_4243 0 1 tie_x0
xfeed_4242 0 1 tie_x0
xfeed_4241 0 1 tie_x0
xfeed_4240 0 1 tie_x0
xfeed_3719 0 1 tie_x0
xfeed_3718 0 1 tie_x0
xfeed_3717 0 1 tie_x0
xfeed_3716 0 1 tie_x0
xfeed_3715 0 1 tie_x0
xfeed_3714 0 1 tie_x0
xfeed_3713 0 1 tie_x0
xfeed_3712 0 1 tie_x0
xfeed_3711 0 1 tie_x0
xfeed_3710 0 1 tie_x0
xfeed_40 0 1 tie_x0
xfeed_41 0 1 tie_x0
xfeed_42 0 1 tie_x0
xfeed_43 0 1 tie_x0
xfeed_44 0 1 tie_x0
xfeed_45 0 1 tie_x0
xfeed_46 0 1 tie_x0
xfeed_8569 0 1 tie_x0
xfeed_8568 0 1 rowend_x0
xfeed_8567 0 1 tie_x0
xfeed_8566 0 1 tie_x0
xfeed_8565 0 1 tie_x0
xfeed_8564 0 1 tie_x0
xfeed_8563 0 1 tie_x0
xfeed_8562 0 1 tie_x0
xfeed_8561 0 1 tie_x0
xfeed_8560 0 1 tie_x0
xfeed_4259 0 1 tie_x0
xfeed_4258 0 1 tie_x0
xfeed_4257 0 1 tie_x0
xfeed_4256 0 1 tie_x0
xfeed_4255 0 1 tie_x0
xfeed_4254 0 1 tie_x0
xfeed_4253 0 1 tie_x0
xfeed_4252 0 1 tie_x0
xfeed_4251 0 1 tie_x0
xfeed_4250 0 1 tie_x0
xfeed_3729 0 1 tie_x0
xfeed_3728 0 1 tie_x0
xfeed_3727 0 1 tie_x0
xfeed_3726 0 1 tie_x0
xfeed_3725 0 1 tie_x0
xfeed_3724 0 1 tie_x0
xfeed_3723 0 1 tie_x0
xfeed_3722 0 1 rowend_x0
xfeed_3721 0 1 tie_x0
xfeed_3720 0 1 tie_x0
xfeed_47 0 1 tie_x0
xfeed_48 0 1 tie_x0
xfeed_49 0 1 tie_x0
xfeed_50 0 1 tie_x0
xfeed_51 0 1 tie_x0
xfeed_52 0 1 tie_x0
xfeed_53 0 1 tie_x0
xfeed_8579 0 1 tie_x0
xfeed_8578 0 1 tie_x0
xfeed_8577 0 1 tie_x0
xfeed_8576 0 1 tie_x0
xfeed_8575 0 1 tie_x0
xfeed_8574 0 1 tie_x0
xfeed_8573 0 1 tie_x0
xfeed_8572 0 1 tie_x0
xfeed_8571 0 1 tie_x0
xfeed_8570 0 1 tie_x0
xfeed_4269 0 1 tie_x0
xfeed_4268 0 1 tie_x0
xfeed_4267 0 1 tie_x0
xfeed_4266 0 1 tie_x0
xfeed_4265 0 1 tie_x0
xfeed_4264 0 1 tie_x0
xfeed_4263 0 1 tie_x0
xfeed_4262 0 1 tie_x0
xfeed_4261 0 1 tie_x0
xfeed_4260 0 1 tie_x0
xfeed_3739 0 1 tie_x0
xfeed_3738 0 1 tie_x0
xfeed_3737 0 1 tie_x0
xfeed_3736 0 1 tie_x0
xfeed_3735 0 1 tie_x0
xfeed_3734 0 1 tie_x0
xfeed_3733 0 1 tie_x0
xfeed_3732 0 1 tie_x0
xfeed_3731 0 1 tie_x0
xfeed_3730 0 1 tie_x0
xfeed_54 0 1 tie_x0
xfeed_55 0 1 tie_x0
xfeed_56 0 1 tie_x0
xfeed_57 0 1 tie_x0
xfeed_58 0 1 tie_x0
xfeed_59 0 1 tie_x0
xfeed_60 0 1 tie_x0
xfeed_8589 0 1 tie_x0
xfeed_8588 0 1 tie_x0
xfeed_8587 0 1 tie_x0
xfeed_8586 0 1 tie_x0
xfeed_8585 0 1 tie_x0
xfeed_8584 0 1 tie_x0
xfeed_8583 0 1 tie_x0
xfeed_8582 0 1 tie_x0
xfeed_8581 0 1 tie_x0
xfeed_8580 0 1 tie_x0
xfeed_4279 0 1 tie_x0
xfeed_4278 0 1 tie_x0
xfeed_4277 0 1 tie_x0
xfeed_4276 0 1 tie_x0
xfeed_4275 0 1 tie_x0
xfeed_4274 0 1 tie_x0
xfeed_4273 0 1 tie_x0
xfeed_4272 0 1 tie_x0
xfeed_4271 0 1 tie_x0
xfeed_4270 0 1 tie_x0
xfeed_3749 0 1 tie_x0
xfeed_3748 0 1 tie_x0
xfeed_3747 0 1 rowend_x0
xfeed_3746 0 1 tie_x0
xfeed_3745 0 1 tie_x0
xfeed_3744 0 1 tie_x0
xfeed_3743 0 1 tie_x0
xfeed_3742 0 1 tie_x0
xfeed_3741 0 1 tie_x0
xfeed_3740 0 1 tie_x0
xsubckt_60_na4_x1 0 1 211 17 12 16 11 na4_x1
xfeed_61 0 1 tie_x0
xfeed_62 0 1 tie_x0
xfeed_63 0 1 tie_x0
xfeed_64 0 1 tie_x0
xfeed_65 0 1 tie_x0
xfeed_66 0 1 tie_x0
xfeed_67 0 1 tie_x0
xfeed_68 0 1 tie_x0
xfeed_69 0 1 tie_x0
xsubckt_95_ao22_x2 0 1 222 180 182 187 ao22_x2
xsubckt_120_a2_x2 0 1 159 77 6 a2_x2
xfeed_8599 0 1 tie_x0
xfeed_8598 0 1 tie_x0
xfeed_8597 0 1 tie_x0
xfeed_8596 0 1 tie_x0
xfeed_8595 0 1 tie_x0
xfeed_8594 0 1 tie_x0
xfeed_8593 0 1 tie_x0
xfeed_8592 0 1 tie_x0
xfeed_8591 0 1 tie_x0
xfeed_8590 0 1 tie_x0
xfeed_4289 0 1 tie_x0
xfeed_4288 0 1 tie_x0
xfeed_4287 0 1 tie_x0
xfeed_4286 0 1 tie_x0
xfeed_4285 0 1 tie_x0
xfeed_4284 0 1 tie_x0
xfeed_4283 0 1 tie_x0
xfeed_4282 0 1 tie_x0
xfeed_4281 0 1 tie_x0
xfeed_4280 0 1 tie_x0
xfeed_3759 0 1 tie_x0
xfeed_3758 0 1 tie_x0
xfeed_3757 0 1 tie_x0
xfeed_3756 0 1 tie_x0
xfeed_3755 0 1 tie_x0
xfeed_3754 0 1 tie_x0
xfeed_3753 0 1 tie_x0
xfeed_3752 0 1 tie_x0
xfeed_3751 0 1 tie_x0
xfeed_3750 0 1 tie_x0
xfeed_70 0 1 tie_x0
xfeed_71 0 1 tie_x0
xfeed_72 0 1 tie_x0
xfeed_73 0 1 tie_x0
xfeed_74 0 1 tie_x0
xfeed_75 0 1 tie_x0
xfeed_76 0 1 tie_x0
xfeed_77 0 1 tie_x0
xfeed_78 0 1 tie_x0
xfeed_79 0 1 tie_x0
xfeed_4299 0 1 tie_x0
xfeed_4298 0 1 tie_x0
xfeed_4297 0 1 tie_x0
xfeed_4296 0 1 tie_x0
xfeed_4295 0 1 tie_x0
xfeed_4294 0 1 tie_x0
xfeed_4293 0 1 tie_x0
xfeed_4292 0 1 tie_x0
xfeed_4291 0 1 tie_x0
xfeed_4290 0 1 tie_x0
xfeed_3768 0 1 tie_x0
xfeed_3767 0 1 tie_x0
xfeed_3766 0 1 tie_x0
xfeed_3765 0 1 tie_x0
xfeed_3764 0 1 tie_x0
xfeed_3763 0 1 tie_x0
xfeed_3762 0 1 tie_x0
xfeed_3761 0 1 tie_x0
xfeed_3760 0 1 tie_x0
xsubckt_163_sff1_x4 0 1 74 214 53 sff1_x4
xfeed_80 0 1 tie_x0
xfeed_81 0 1 tie_x0
xfeed_82 0 1 tie_x0
xfeed_83 0 1 tie_x0
xfeed_84 0 1 tie_x0
xfeed_85 0 1 tie_x0
xfeed_86 0 1 tie_x0
xfeed_87 0 1 tie_x0
xfeed_88 0 1 tie_x0
xfeed_89 0 1 tie_x0
xfeed_3769 0 1 tie_x0
xsubckt_77_a2_x2 0 1 195 16 11 a2_x2
xsubckt_57_a2_x2 0 1 82 12 16 a2_x2
xfeed_3775 0 1 tie_x0
xfeed_3774 0 1 tie_x0
xfeed_3773 0 1 tie_x0
xfeed_3772 0 1 rowend_x0
xfeed_3771 0 1 tie_x0
xfeed_3770 0 1 tie_x0
xsubckt_115_nxr2_x1 0 1 163 167 164 nxr2_x1
xsubckt_159_sff1_x4 0 1 78 218 21 sff1_x4
xfeed_90 0 1 tie_x0
xfeed_91 0 1 tie_x0
xfeed_92 0 1 tie_x0
xfeed_93 0 1 tie_x0
xfeed_94 0 1 tie_x0
xfeed_95 0 1 tie_x0
xfeed_96 0 1 tie_x0
xfeed_97 0 1 tie_x0
xfeed_98 0 1 tie_x0
xfeed_99 0 1 tie_x0
xfeed_3779 0 1 tie_x0
xfeed_3778 0 1 tie_x0
xfeed_3777 0 1 tie_x0
xfeed_3776 0 1 tie_x0
xfeed_8709 0 1 tie_x0
xfeed_8708 0 1 tie_x0
xfeed_8707 0 1 tie_x0
xfeed_8706 0 1 tie_x0
xfeed_8705 0 1 tie_x0
xfeed_8704 0 1 tie_x0
xfeed_8703 0 1 tie_x0
xfeed_8702 0 1 tie_x0
xfeed_8701 0 1 tie_x0
xfeed_8700 0 1 tie_x0
xfeed_3782 0 1 tie_x0
xfeed_3781 0 1 tie_x0
xfeed_3780 0 1 tie_x0
xfeed_3789 0 1 tie_x0
xfeed_3788 0 1 tie_x0
xfeed_3787 0 1 tie_x0
xfeed_3786 0 1 tie_x0
xfeed_3785 0 1 tie_x0
xfeed_3784 0 1 tie_x0
xfeed_3783 0 1 tie_x0
xfeed_8719 0 1 tie_x0
xfeed_8718 0 1 tie_x0
xfeed_8717 0 1 tie_x0
xfeed_8716 0 1 tie_x0
xfeed_8715 0 1 tie_x0
xfeed_8714 0 1 tie_x0
xfeed_8713 0 1 tie_x0
xfeed_8712 0 1 tie_x0
xfeed_8711 0 1 tie_x0
xfeed_8710 0 1 tie_x0
xfeed_4409 0 1 tie_x0
xfeed_4408 0 1 tie_x0
xfeed_4407 0 1 tie_x0
xfeed_4406 0 1 tie_x0
xfeed_4405 0 1 tie_x0
xfeed_4404 0 1 tie_x0
xfeed_4403 0 1 tie_x0
xfeed_4402 0 1 tie_x0
xfeed_4401 0 1 tie_x0
xfeed_4400 0 1 tie_x0
xfeed_3799 0 1 tie_x0
xfeed_3798 0 1 tie_x0
xfeed_3797 0 1 rowend_x0
xfeed_3796 0 1 tie_x0
xfeed_3795 0 1 tie_x0
xfeed_3794 0 1 tie_x0
xfeed_3793 0 1 tie_x0
xfeed_3792 0 1 tie_x0
xfeed_3791 0 1 tie_x0
xfeed_3790 0 1 tie_x0
xfeed_8729 0 1 tie_x0
xfeed_8728 0 1 tie_x0
xfeed_8727 0 1 tie_x0
xfeed_8726 0 1 tie_x0
xfeed_8725 0 1 tie_x0
xfeed_8724 0 1 tie_x0
xfeed_8723 0 1 rowend_x0
xfeed_8722 0 1 tie_x0
xfeed_8721 0 1 tie_x0
xfeed_8720 0 1 tie_x0
xfeed_4419 0 1 tie_x0
xfeed_4418 0 1 tie_x0
xfeed_4417 0 1 tie_x0
xfeed_4416 0 1 tie_x0
xfeed_4415 0 1 tie_x0
xfeed_4414 0 1 tie_x0
xfeed_4413 0 1 tie_x0
xfeed_4412 0 1 tie_x0
xfeed_4411 0 1 tie_x0
xfeed_4410 0 1 tie_x0
xfeed_8739 0 1 tie_x0
xfeed_8738 0 1 tie_x0
xfeed_8737 0 1 tie_x0
xfeed_8736 0 1 tie_x0
xfeed_8735 0 1 tie_x0
xfeed_8734 0 1 tie_x0
xfeed_8733 0 1 tie_x0
xfeed_8732 0 1 tie_x0
xfeed_8731 0 1 tie_x0
xfeed_8730 0 1 tie_x0
xfeed_4429 0 1 tie_x0
xfeed_4428 0 1 tie_x0
xfeed_4427 0 1 tie_x0
xfeed_4426 0 1 tie_x0
xfeed_4425 0 1 tie_x0
xfeed_4424 0 1 tie_x0
xfeed_4423 0 1 tie_x0
xfeed_4422 0 1 tie_x0
xfeed_4421 0 1 tie_x0
xfeed_4420 0 1 tie_x0
xsubckt_42_a3_x2 0 1 96 101 99 98 a3_x2
xfeed_8747 0 1 tie_x0
xfeed_8746 0 1 tie_x0
xfeed_8745 0 1 tie_x0
xfeed_8744 0 1 tie_x0
xfeed_8743 0 1 tie_x0
xfeed_8742 0 1 tie_x0
xfeed_8741 0 1 tie_x0
xfeed_8740 0 1 tie_x0
xfeed_4439 0 1 tie_x0
xfeed_4438 0 1 tie_x0
xfeed_4437 0 1 tie_x0
xfeed_4436 0 1 tie_x0
xfeed_4435 0 1 tie_x0
xfeed_4434 0 1 tie_x0
xfeed_4433 0 1 tie_x0
xfeed_4432 0 1 tie_x0
xfeed_4431 0 1 tie_x0
xfeed_4430 0 1 tie_x0
xfeed_3908 0 1 tie_x0
xfeed_3907 0 1 tie_x0
xfeed_3906 0 1 tie_x0
xfeed_3905 0 1 tie_x0
xfeed_3904 0 1 tie_x0
xfeed_3903 0 1 tie_x0
xfeed_3902 0 1 tie_x0
xfeed_3901 0 1 tie_x0
xfeed_3900 0 1 tie_x0
xsubckt_97_xr2_x4 0 1 178 81 10 xr2_x4
xfeed_8749 0 1 tie_x0
xfeed_8748 0 1 tie_x0
xfeed_3909 0 1 tie_x0
xfeed_8754 0 1 tie_x0
xfeed_8753 0 1 tie_x0
xfeed_8752 0 1 tie_x0
xfeed_8751 0 1 tie_x0
xfeed_8750 0 1 tie_x0
xfeed_4449 0 1 tie_x0
xfeed_4448 0 1 tie_x0
xfeed_4447 0 1 tie_x0
xfeed_4446 0 1 tie_x0
xfeed_4445 0 1 tie_x0
xfeed_4444 0 1 tie_x0
xfeed_4443 0 1 tie_x0
xfeed_4442 0 1 tie_x0
xfeed_4441 0 1 tie_x0
xfeed_4440 0 1 tie_x0
xfeed_3915 0 1 tie_x0
xfeed_3914 0 1 tie_x0
xfeed_3913 0 1 tie_x0
xfeed_3912 0 1 tie_x0
xfeed_3911 0 1 tie_x0
xfeed_3910 0 1 tie_x0
xfeed_8759 0 1 tie_x0
xfeed_8758 0 1 tie_x0
xfeed_8757 0 1 tie_x0
xfeed_8756 0 1 tie_x0
xfeed_8755 0 1 tie_x0
xfeed_3919 0 1 tie_x0
xfeed_3918 0 1 tie_x0
xfeed_3917 0 1 tie_x0
xfeed_3916 0 1 tie_x0
xfeed_8761 0 1 tie_x0
xfeed_8760 0 1 tie_x0
xfeed_4459 0 1 tie_x0
xfeed_4458 0 1 tie_x0
xfeed_4457 0 1 tie_x0
xfeed_4456 0 1 tie_x0
xfeed_4455 0 1 tie_x0
xfeed_4454 0 1 tie_x0
xfeed_4453 0 1 tie_x0
xfeed_4452 0 1 tie_x0
xfeed_4451 0 1 tie_x0
xfeed_4450 0 1 tie_x0
xfeed_3922 0 1 tie_x0
xfeed_3921 0 1 tie_x0
xfeed_3920 0 1 tie_x0
xfeed_8769 0 1 tie_x0
xfeed_8768 0 1 tie_x0
xfeed_8767 0 1 tie_x0
xfeed_8766 0 1 tie_x0
xfeed_8765 0 1 tie_x0
xfeed_8764 0 1 tie_x0
xfeed_8763 0 1 tie_x0
xfeed_8762 0 1 tie_x0
xfeed_3929 0 1 tie_x0
xfeed_3928 0 1 tie_x0
xfeed_3927 0 1 tie_x0
xfeed_3926 0 1 tie_x0
xfeed_3925 0 1 tie_x0
xfeed_3924 0 1 tie_x0
xfeed_3923 0 1 tie_x0
xfeed_4468 0 1 tie_x0
xfeed_4467 0 1 tie_x0
xfeed_4466 0 1 tie_x0
xfeed_4465 0 1 tie_x0
xfeed_4464 0 1 tie_x0
xfeed_4463 0 1 tie_x0
xfeed_4462 0 1 tie_x0
xfeed_4461 0 1 tie_x0
xfeed_4460 0 1 tie_x0
xsubckt_142_a3_x2 0 1 215 131 141 140 a3_x2
xfeed_8779 0 1 tie_x0
xfeed_8778 0 1 tie_x0
xfeed_8777 0 1 tie_x0
xfeed_8776 0 1 tie_x0
xfeed_8775 0 1 tie_x0
xfeed_8774 0 1 tie_x0
xfeed_8773 0 1 tie_x0
xfeed_8772 0 1 tie_x0
xfeed_8771 0 1 rowend_x0
xfeed_8770 0 1 tie_x0
xfeed_4469 0 1 tie_x0
xfeed_3939 0 1 tie_x0
xfeed_3938 0 1 tie_x0
xfeed_3937 0 1 tie_x0
xfeed_3936 0 1 tie_x0
xfeed_3935 0 1 tie_x0
xfeed_3934 0 1 tie_x0
xfeed_3933 0 1 tie_x0
xfeed_3932 0 1 tie_x0
xfeed_3931 0 1 tie_x0
xfeed_3930 0 1 tie_x0
xfeed_4475 0 1 tie_x0
xfeed_4474 0 1 tie_x0
xfeed_4473 0 1 tie_x0
xfeed_4472 0 1 tie_x0
xfeed_4471 0 1 tie_x0
xfeed_4470 0 1 tie_x0
xsubckt_84_mx2_x2 0 1 224 5 189 2 mx2_x2
xfeed_8789 0 1 tie_x0
xfeed_8788 0 1 tie_x0
xfeed_8787 0 1 tie_x0
xfeed_8786 0 1 tie_x0
xfeed_8785 0 1 tie_x0
xfeed_8784 0 1 tie_x0
xfeed_8783 0 1 tie_x0
xfeed_8782 0 1 tie_x0
xfeed_8781 0 1 tie_x0
xfeed_8780 0 1 tie_x0
xfeed_4479 0 1 tie_x0
xfeed_4478 0 1 tie_x0
xfeed_4477 0 1 tie_x0
xfeed_4476 0 1 tie_x0
xfeed_3949 0 1 tie_x0
xfeed_3948 0 1 tie_x0
xfeed_3947 0 1 tie_x0
xfeed_3946 0 1 tie_x0
xfeed_3945 0 1 tie_x0
xfeed_3944 0 1 tie_x0
xfeed_3943 0 1 tie_x0
xfeed_3942 0 1 tie_x0
xfeed_3941 0 1 tie_x0
xfeed_3940 0 1 tie_x0
xfeed_4482 0 1 tie_x0
xfeed_4481 0 1 tie_x0
xfeed_4480 0 1 tie_x0
xfeed_8795 0 1 tie_x0
xfeed_8794 0 1 tie_x0
xfeed_8793 0 1 tie_x0
xfeed_8792 0 1 tie_x0
xfeed_8791 0 1 tie_x0
xfeed_8790 0 1 tie_x0
xfeed_4489 0 1 tie_x0
xfeed_4488 0 1 tie_x0
xfeed_4487 0 1 tie_x0
xfeed_4486 0 1 tie_x0
xfeed_4485 0 1 tie_x0
xfeed_4484 0 1 tie_x0
xfeed_4483 0 1 tie_x0
xfeed_3959 0 1 tie_x0
xfeed_3958 0 1 tie_x0
xfeed_3957 0 1 tie_x0
xfeed_3956 0 1 tie_x0
xfeed_3955 0 1 tie_x0
xfeed_3954 0 1 tie_x0
xfeed_3953 0 1 rowend_x0
xfeed_3952 0 1 tie_x0
xfeed_3951 0 1 tie_x0
xfeed_3950 0 1 tie_x0
xfeed_5109 0 1 tie_x0
xfeed_5108 0 1 tie_x0
xfeed_5107 0 1 tie_x0
xfeed_5106 0 1 tie_x0
xfeed_5105 0 1 tie_x0
xfeed_5104 0 1 tie_x0
xfeed_5103 0 1 tie_x0
xfeed_5102 0 1 tie_x0
xfeed_5101 0 1 tie_x0
xfeed_5100 0 1 tie_x0
xsubckt_66_nxr2_x1 0 1 205 85 206 nxr2_x1
xsubckt_56_nao22_x1 0 1 83 109 107 112 nao22_x1
xfeed_4499 0 1 tie_x0
xfeed_4498 0 1 tie_x0
xfeed_4497 0 1 tie_x0
xfeed_4496 0 1 tie_x0
xfeed_4495 0 1 tie_x0
xfeed_4494 0 1 tie_x0
xfeed_4493 0 1 tie_x0
xfeed_4492 0 1 tie_x0
xfeed_4491 0 1 tie_x0
xfeed_4490 0 1 tie_x0
xfeed_3969 0 1 tie_x0
xfeed_3968 0 1 tie_x0
xfeed_3967 0 1 tie_x0
xfeed_3966 0 1 tie_x0
xfeed_3965 0 1 tie_x0
xfeed_3964 0 1 tie_x0
xfeed_3963 0 1 tie_x0
xfeed_3962 0 1 tie_x0
xfeed_3961 0 1 tie_x0
xfeed_3960 0 1 tie_x0
xfeed_5119 0 1 tie_x0
xfeed_5118 0 1 tie_x0
xfeed_5117 0 1 tie_x0
xfeed_5116 0 1 tie_x0
xfeed_5115 0 1 tie_x0
xfeed_5114 0 1 tie_x0
xfeed_5113 0 1 tie_x0
xfeed_5112 0 1 tie_x0
xfeed_5111 0 1 tie_x0
xfeed_5110 0 1 tie_x0
xfeed_3979 0 1 tie_x0
xfeed_3978 0 1 tie_x0
xfeed_3977 0 1 tie_x0
xfeed_3976 0 1 tie_x0
xfeed_3975 0 1 tie_x0
xfeed_3974 0 1 tie_x0
xfeed_3973 0 1 tie_x0
xfeed_3972 0 1 tie_x0
xfeed_3971 0 1 tie_x0
xfeed_3970 0 1 tie_x0
xfeed_5129 0 1 tie_x0
xfeed_5128 0 1 tie_x0
xfeed_5127 0 1 tie_x0
xfeed_5126 0 1 tie_x0
xfeed_5125 0 1 tie_x0
xfeed_5124 0 1 tie_x0
xfeed_5123 0 1 tie_x0
xfeed_5122 0 1 tie_x0
xfeed_5121 0 1 tie_x0
xfeed_5120 0 1 tie_x0
xfeed_3989 0 1 tie_x0
xfeed_3988 0 1 tie_x0
xfeed_3987 0 1 tie_x0
xfeed_3986 0 1 tie_x0
xfeed_3985 0 1 tie_x0
xfeed_3984 0 1 tie_x0
xfeed_3983 0 1 tie_x0
xfeed_3982 0 1 tie_x0
xfeed_3981 0 1 tie_x0
xfeed_3980 0 1 tie_x0
xfeed_5139 0 1 tie_x0
xfeed_5138 0 1 tie_x0
xfeed_5137 0 1 tie_x0
xfeed_5136 0 1 tie_x0
xfeed_5135 0 1 tie_x0
xfeed_5134 0 1 tie_x0
xfeed_5133 0 1 tie_x0
xfeed_5132 0 1 tie_x0
xfeed_5131 0 1 tie_x0
xfeed_5130 0 1 tie_x0
xfeed_4608 0 1 tie_x0
xfeed_4607 0 1 tie_x0
xfeed_4606 0 1 tie_x0
xfeed_4605 0 1 tie_x0
xfeed_4604 0 1 tie_x0
xfeed_4603 0 1 tie_x0
xfeed_4602 0 1 tie_x0
xfeed_4601 0 1 tie_x0
xfeed_4600 0 1 tie_x0
xfeed_4609 0 1 tie_x0
xfeed_3999 0 1 tie_x0
xfeed_3998 0 1 tie_x0
xfeed_3997 0 1 tie_x0
xfeed_3996 0 1 tie_x0
xfeed_3995 0 1 tie_x0
xfeed_3994 0 1 tie_x0
xfeed_3993 0 1 tie_x0
xfeed_3992 0 1 tie_x0
xfeed_3991 0 1 tie_x0
xfeed_3990 0 1 tie_x0
xsubckt_12_na2_x1 0 1 125 14 16 na2_x1
xsubckt_38_ao22_x2 0 1 100 114 106 104 ao22_x2
xfeed_5149 0 1 tie_x0
xfeed_5148 0 1 tie_x0
xfeed_5147 0 1 tie_x0
xfeed_5146 0 1 tie_x0
xfeed_5145 0 1 tie_x0
xfeed_5144 0 1 rowend_x0
xfeed_5143 0 1 tie_x0
xfeed_5142 0 1 tie_x0
xfeed_5141 0 1 tie_x0
xfeed_5140 0 1 tie_x0
xfeed_4615 0 1 tie_x0
xfeed_4614 0 1 tie_x0
xfeed_4613 0 1 tie_x0
xfeed_4612 0 1 tie_x0
xfeed_4611 0 1 tie_x0
xfeed_4610 0 1 tie_x0
xfeed_4619 0 1 tie_x0
xfeed_4618 0 1 tie_x0
xfeed_4617 0 1 tie_x0
xfeed_4616 0 1 tie_x0
xfeed_5159 0 1 tie_x0
xfeed_5158 0 1 tie_x0
xfeed_5157 0 1 tie_x0
xfeed_5156 0 1 tie_x0
xfeed_5155 0 1 tie_x0
xfeed_5154 0 1 tie_x0
xfeed_5153 0 1 tie_x0
xfeed_5152 0 1 tie_x0
xfeed_5151 0 1 tie_x0
xfeed_5150 0 1 tie_x0
xfeed_4622 0 1 tie_x0
xfeed_4621 0 1 tie_x0
xfeed_4620 0 1 tie_x0
xfeed_4629 0 1 tie_x0
xfeed_4628 0 1 tie_x0
xfeed_4627 0 1 tie_x0
xfeed_4626 0 1 tie_x0
xfeed_4625 0 1 tie_x0
xfeed_4624 0 1 tie_x0
xfeed_4623 0 1 tie_x0
xfeed_5168 0 1 tie_x0
xfeed_5167 0 1 tie_x0
xfeed_5166 0 1 tie_x0
xfeed_5165 0 1 tie_x0
xfeed_5164 0 1 tie_x0
xfeed_5163 0 1 tie_x0
xfeed_5162 0 1 tie_x0
xfeed_5161 0 1 tie_x0
xfeed_5160 0 1 tie_x0
xfeed_5169 0 1 tie_x0
xfeed_4639 0 1 tie_x0
xfeed_4638 0 1 tie_x0
xfeed_4637 0 1 tie_x0
xfeed_4636 0 1 tie_x0
xfeed_4635 0 1 tie_x0
xfeed_4634 0 1 tie_x0
xfeed_4633 0 1 tie_x0
xfeed_4632 0 1 tie_x0
xfeed_4631 0 1 tie_x0
xfeed_4630 0 1 tie_x0
xfeed_5175 0 1 tie_x0
xfeed_5174 0 1 tie_x0
xfeed_5173 0 1 tie_x0
xfeed_5172 0 1 tie_x0
xfeed_5171 0 1 tie_x0
xfeed_5170 0 1 rowend_x0
xfeed_5179 0 1 tie_x0
xfeed_5178 0 1 tie_x0
xfeed_5177 0 1 tie_x0
xfeed_5176 0 1 tie_x0
xfeed_4649 0 1 tie_x0
xfeed_4648 0 1 tie_x0
xfeed_4647 0 1 tie_x0
xfeed_4646 0 1 tie_x0
xfeed_4645 0 1 tie_x0
xfeed_4644 0 1 tie_x0
xfeed_4643 0 1 tie_x0
xfeed_4642 0 1 tie_x0
xfeed_4641 0 1 tie_x0
xfeed_4640 0 1 tie_x0
xsubckt_88_nao22_x1 0 1 185 211 132 133 nao22_x1
xfeed_5182 0 1 tie_x0
xfeed_5181 0 1 tie_x0
xfeed_5180 0 1 tie_x0
xfeed_5189 0 1 tie_x0
xfeed_5188 0 1 tie_x0
xfeed_5187 0 1 tie_x0
xfeed_5186 0 1 tie_x0
xfeed_5185 0 1 tie_x0
xfeed_5184 0 1 tie_x0
xfeed_5183 0 1 tie_x0
xfeed_4659 0 1 tie_x0
xfeed_4658 0 1 tie_x0
xfeed_4657 0 1 tie_x0
xfeed_4656 0 1 tie_x0
xfeed_4655 0 1 tie_x0
xfeed_4654 0 1 tie_x0
xfeed_4653 0 1 tie_x0
xfeed_4652 0 1 tie_x0
xfeed_4651 0 1 tie_x0
xfeed_4650 0 1 tie_x0
xsubckt_71_nao22_x1 0 1 200 131 91 203 nao22_x1
xsubckt_125_a2_x2 0 1 217 131 155 a2_x2
xfeed_5199 0 1 tie_x0
xfeed_5198 0 1 tie_x0
xfeed_5197 0 1 tie_x0
xfeed_5196 0 1 tie_x0
xfeed_5195 0 1 rowend_x0
xfeed_5194 0 1 tie_x0
xfeed_5193 0 1 tie_x0
xfeed_5192 0 1 tie_x0
xfeed_5191 0 1 tie_x0
xfeed_5190 0 1 tie_x0
xfeed_4669 0 1 tie_x0
xfeed_4668 0 1 tie_x0
xfeed_4667 0 1 tie_x0
xfeed_4666 0 1 tie_x0
xfeed_4665 0 1 tie_x0
xfeed_4664 0 1 tie_x0
xfeed_4663 0 1 tie_x0
xfeed_4662 0 1 tie_x0
xfeed_4661 0 1 tie_x0
xfeed_4660 0 1 tie_x0
xfeed_4679 0 1 tie_x0
xfeed_4678 0 1 tie_x0
xfeed_4677 0 1 tie_x0
xfeed_4676 0 1 tie_x0
xfeed_4675 0 1 tie_x0
xfeed_4674 0 1 tie_x0
xfeed_4673 0 1 tie_x0
xfeed_4672 0 1 tie_x0
xfeed_4671 0 1 tie_x0
xfeed_4670 0 1 tie_x0
xfeed_4689 0 1 tie_x0
xfeed_4688 0 1 tie_x0
xfeed_4687 0 1 tie_x0
xfeed_4686 0 1 tie_x0
xfeed_4685 0 1 tie_x0
xfeed_4684 0 1 tie_x0
xfeed_4683 0 1 tie_x0
xfeed_4682 0 1 tie_x0
xfeed_4681 0 1 tie_x0
xfeed_4680 0 1 tie_x0
xsubckt_105_na2_x1 0 1 172 79 8 na2_x1
xfeed_5308 0 1 tie_x0
xfeed_5307 0 1 tie_x0
xfeed_5306 0 1 tie_x0
xfeed_5305 0 1 tie_x0
xfeed_5304 0 1 tie_x0
xfeed_5303 0 1 tie_x0
xfeed_5302 0 1 tie_x0
xfeed_5301 0 1 tie_x0
xfeed_5300 0 1 tie_x0
xfeed_5309 0 1 tie_x0
xfeed_4699 0 1 rowend_x0
xfeed_4698 0 1 tie_x0
xfeed_4697 0 1 tie_x0
xfeed_4696 0 1 tie_x0
xfeed_4695 0 1 tie_x0
xfeed_4694 0 1 tie_x0
xfeed_4693 0 1 tie_x0
xfeed_4692 0 1 tie_x0
xfeed_4691 0 1 tie_x0
xfeed_4690 0 1 tie_x0
xfeed_5315 0 1 tie_x0
xfeed_5314 0 1 tie_x0
xfeed_5313 0 1 tie_x0
xfeed_5312 0 1 tie_x0
xfeed_5311 0 1 tie_x0
xfeed_5310 0 1 tie_x0
xfeed_1000 0 1 tie_x0
xfeed_1001 0 1 tie_x0
xfeed_1002 0 1 tie_x0
xfeed_1003 0 1 tie_x0
xfeed_1004 0 1 tie_x0
xfeed_1005 0 1 tie_x0
xfeed_1006 0 1 tie_x0
xfeed_1007 0 1 tie_x0
xfeed_1008 0 1 tie_x0
xfeed_1009 0 1 tie_x0
xfeed_5319 0 1 tie_x0
xfeed_5318 0 1 tie_x0
xfeed_5317 0 1 tie_x0
xfeed_5316 0 1 tie_x0
xfeed_5322 0 1 tie_x0
xfeed_5321 0 1 tie_x0
xfeed_5320 0 1 tie_x0
xfeed_1010 0 1 tie_x0
xfeed_1011 0 1 tie_x0
xfeed_1012 0 1 tie_x0
xfeed_1013 0 1 tie_x0
xfeed_1014 0 1 tie_x0
xfeed_1015 0 1 tie_x0
xfeed_1016 0 1 tie_x0
xfeed_1017 0 1 tie_x0
xfeed_1018 0 1 tie_x0
xfeed_1019 0 1 tie_x0
xfeed_5329 0 1 tie_x0
xfeed_5328 0 1 tie_x0
xfeed_5327 0 1 tie_x0
xfeed_5326 0 1 tie_x0
xfeed_5325 0 1 tie_x0
xfeed_5324 0 1 tie_x0
xfeed_5323 0 1 tie_x0
xfeed_1020 0 1 tie_x0
xfeed_1021 0 1 tie_x0
xfeed_1022 0 1 tie_x0
xfeed_1023 0 1 tie_x0
xfeed_1024 0 1 tie_x0
xfeed_1025 0 1 tie_x0
xfeed_1026 0 1 tie_x0
xfeed_1027 0 1 tie_x0
xfeed_1028 0 1 tie_x0
xfeed_1029 0 1 tie_x0
xfeed_5339 0 1 tie_x0
xfeed_5338 0 1 tie_x0
xfeed_5337 0 1 tie_x0
xfeed_5336 0 1 tie_x0
xfeed_5335 0 1 tie_x0
xfeed_5334 0 1 tie_x0
xfeed_5333 0 1 tie_x0
xfeed_5332 0 1 rowend_x0
xfeed_5331 0 1 tie_x0
xfeed_5330 0 1 tie_x0
xfeed_4809 0 1 tie_x0
xfeed_4808 0 1 tie_x0
xfeed_4807 0 1 tie_x0
xfeed_4806 0 1 tie_x0
xfeed_4805 0 1 tie_x0
xfeed_4804 0 1 tie_x0
xfeed_4803 0 1 tie_x0
xfeed_4802 0 1 tie_x0
xfeed_4801 0 1 tie_x0
xfeed_4800 0 1 rowend_x0
xsubckt_47_a3_x2 0 1 91 118 95 93 a3_x2
xsubckt_150_sff1_x4 0 1 8 227 24 sff1_x4
xfeed_1030 0 1 tie_x0
xfeed_1031 0 1 tie_x0
xfeed_1032 0 1 tie_x0
xfeed_1033 0 1 tie_x0
xfeed_1034 0 1 tie_x0
xfeed_1035 0 1 tie_x0
xfeed_1036 0 1 tie_x0
xfeed_5349 0 1 tie_x0
xfeed_5348 0 1 tie_x0
xfeed_5347 0 1 tie_x0
xfeed_5346 0 1 tie_x0
xfeed_5345 0 1 tie_x0
xfeed_5344 0 1 tie_x0
xfeed_5343 0 1 tie_x0
xfeed_5342 0 1 tie_x0
xfeed_5341 0 1 tie_x0
xfeed_5340 0 1 tie_x0
xfeed_4819 0 1 tie_x0
xfeed_4818 0 1 tie_x0
xfeed_4817 0 1 tie_x0
xfeed_4816 0 1 tie_x0
xfeed_4815 0 1 tie_x0
xfeed_4814 0 1 tie_x0
xfeed_4813 0 1 tie_x0
xfeed_4812 0 1 tie_x0
xfeed_4811 0 1 tie_x0
xfeed_4810 0 1 tie_x0
xsubckt_102_nxr2_x1 0 1 174 179 175 nxr2_x1
xfeed_1037 0 1 tie_x0
xfeed_1038 0 1 tie_x0
xfeed_1039 0 1 tie_x0
xfeed_1040 0 1 tie_x0
xfeed_1041 0 1 tie_x0
xfeed_1042 0 1 tie_x0
xfeed_1043 0 1 tie_x0
xfeed_5359 0 1 tie_x0
xfeed_5358 0 1 tie_x0
xfeed_5357 0 1 tie_x0
xfeed_5356 0 1 tie_x0
xfeed_5355 0 1 tie_x0
xfeed_5354 0 1 tie_x0
xfeed_5353 0 1 rowend_x0
xfeed_5352 0 1 tie_x0
xfeed_5351 0 1 tie_x0
xfeed_5350 0 1 tie_x0
xfeed_4829 0 1 tie_x0
xfeed_4828 0 1 tie_x0
xfeed_4827 0 1 tie_x0
xfeed_4826 0 1 rowend_x0
xfeed_4825 0 1 tie_x0
xfeed_4824 0 1 tie_x0
xfeed_4823 0 1 tie_x0
xfeed_4822 0 1 tie_x0
xfeed_4821 0 1 tie_x0
xfeed_4820 0 1 tie_x0
xfeed_1044 0 1 tie_x0
xfeed_1045 0 1 tie_x0
xfeed_1046 0 1 tie_x0
xfeed_1047 0 1 tie_x0
xfeed_1048 0 1 tie_x0
xfeed_1049 0 1 tie_x0
xfeed_1050 0 1 tie_x0
xfeed_5369 0 1 tie_x0
xfeed_5368 0 1 tie_x0
xfeed_5367 0 1 tie_x0
xfeed_5366 0 1 tie_x0
xfeed_5365 0 1 tie_x0
xfeed_5364 0 1 tie_x0
xfeed_5363 0 1 tie_x0
xfeed_5362 0 1 tie_x0
xfeed_5361 0 1 tie_x0
xfeed_5360 0 1 tie_x0
xfeed_4839 0 1 tie_x0
xfeed_4838 0 1 tie_x0
xfeed_4837 0 1 tie_x0
xfeed_4836 0 1 tie_x0
xfeed_4835 0 1 tie_x0
xfeed_4834 0 1 tie_x0
xfeed_4833 0 1 tie_x0
xfeed_4832 0 1 tie_x0
xfeed_4831 0 1 tie_x0
xfeed_4830 0 1 tie_x0
xfeed_1051 0 1 tie_x0
xfeed_1052 0 1 tie_x0
xfeed_1053 0 1 tie_x0
xfeed_1054 0 1 tie_x0
xfeed_1055 0 1 tie_x0
xfeed_1056 0 1 tie_x0
xfeed_1057 0 1 tie_x0
xfeed_1058 0 1 tie_x0
xfeed_1059 0 1 tie_x0
xfeed_5379 0 1 tie_x0
xfeed_5378 0 1 tie_x0
xfeed_5377 0 1 tie_x0
xfeed_5376 0 1 tie_x0
xfeed_5375 0 1 tie_x0
xfeed_5374 0 1 tie_x0
xfeed_5373 0 1 tie_x0
xfeed_5372 0 1 tie_x0
xfeed_5371 0 1 tie_x0
xfeed_5370 0 1 tie_x0
xfeed_4849 0 1 tie_x0
xfeed_4848 0 1 tie_x0
xfeed_4847 0 1 tie_x0
xfeed_4846 0 1 tie_x0
xfeed_4845 0 1 tie_x0
xfeed_4844 0 1 tie_x0
xfeed_4843 0 1 tie_x0
xfeed_4842 0 1 tie_x0
xfeed_4841 0 1 tie_x0
xfeed_4840 0 1 tie_x0
xsubckt_75_nao22_x1 0 1 197 208 207 85 nao22_x1
xfeed_1060 0 1 tie_x0
xfeed_1061 0 1 tie_x0
xfeed_1062 0 1 tie_x0
xfeed_1063 0 1 tie_x0
xfeed_1064 0 1 tie_x0
xfeed_1065 0 1 tie_x0
xfeed_1066 0 1 tie_x0
xfeed_1067 0 1 tie_x0
xfeed_1068 0 1 tie_x0
xfeed_1069 0 1 tie_x0
xfeed_5389 0 1 tie_x0
xfeed_5388 0 1 tie_x0
xfeed_5387 0 1 tie_x0
xfeed_5386 0 1 tie_x0
xfeed_5385 0 1 tie_x0
xfeed_5384 0 1 tie_x0
xfeed_5383 0 1 tie_x0
xfeed_5382 0 1 tie_x0
xfeed_5381 0 1 tie_x0
xfeed_5380 0 1 tie_x0
xfeed_4859 0 1 tie_x0
xfeed_4858 0 1 tie_x0
xfeed_4857 0 1 tie_x0
xfeed_4856 0 1 tie_x0
xfeed_4855 0 1 tie_x0
xfeed_4854 0 1 tie_x0
xfeed_4853 0 1 tie_x0
xfeed_4852 0 1 tie_x0
xfeed_4851 0 1 tie_x0
xfeed_4850 0 1 tie_x0
xfeed_1070 0 1 tie_x0
xfeed_1071 0 1 tie_x0
xfeed_1072 0 1 tie_x0
xfeed_1073 0 1 tie_x0
xfeed_1074 0 1 tie_x0
xfeed_1075 0 1 tie_x0
xfeed_1076 0 1 tie_x0
xfeed_1077 0 1 tie_x0
xfeed_1078 0 1 tie_x0
xfeed_1079 0 1 rowend_x0
xfeed_6008 0 1 tie_x0
xfeed_6007 0 1 tie_x0
xfeed_6006 0 1 tie_x0
xfeed_6005 0 1 tie_x0
xfeed_6004 0 1 tie_x0
xfeed_6003 0 1 tie_x0
xfeed_6002 0 1 tie_x0
xfeed_6001 0 1 tie_x0
xfeed_6000 0 1 tie_x0
xfeed_6009 0 1 tie_x0
xfeed_5399 0 1 tie_x0
xfeed_5398 0 1 tie_x0
xfeed_5397 0 1 tie_x0
xfeed_5396 0 1 tie_x0
xfeed_5395 0 1 tie_x0
xfeed_5394 0 1 tie_x0
xfeed_5393 0 1 tie_x0
xfeed_5392 0 1 tie_x0
xfeed_5391 0 1 tie_x0
xfeed_5390 0 1 tie_x0
xfeed_4869 0 1 tie_x0
xfeed_4868 0 1 tie_x0
xfeed_4867 0 1 tie_x0
xfeed_4866 0 1 tie_x0
xfeed_4865 0 1 tie_x0
xfeed_4864 0 1 tie_x0
xfeed_4863 0 1 tie_x0
xfeed_4862 0 1 tie_x0
xfeed_4861 0 1 tie_x0
xfeed_4860 0 1 tie_x0
xfeed_1080 0 1 tie_x0
xfeed_1081 0 1 tie_x0
xfeed_1082 0 1 tie_x0
xfeed_1083 0 1 tie_x0
xfeed_1084 0 1 tie_x0
xfeed_1085 0 1 tie_x0
xfeed_1086 0 1 tie_x0
xfeed_1087 0 1 tie_x0
xfeed_1088 0 1 tie_x0
xfeed_1089 0 1 tie_x0
xfeed_6015 0 1 tie_x0
xfeed_6014 0 1 tie_x0
xfeed_6013 0 1 tie_x0
xfeed_6012 0 1 tie_x0
xfeed_6011 0 1 tie_x0
xfeed_6010 0 1 tie_x0
xfeed_6019 0 1 tie_x0
xfeed_6018 0 1 tie_x0
xfeed_6017 0 1 tie_x0
xfeed_6016 0 1 tie_x0
xfeed_4879 0 1 tie_x0
xfeed_4878 0 1 tie_x0
xfeed_4877 0 1 tie_x0
xfeed_4876 0 1 tie_x0
xfeed_4875 0 1 tie_x0
xfeed_4874 0 1 tie_x0
xfeed_4873 0 1 tie_x0
xfeed_4872 0 1 tie_x0
xfeed_4871 0 1 tie_x0
xfeed_4870 0 1 tie_x0
xsubckt_68_nxr2_x1 0 1 203 87 205 nxr2_x1
xfeed_1090 0 1 tie_x0
xfeed_1091 0 1 tie_x0
xfeed_1092 0 1 tie_x0
xfeed_1093 0 1 tie_x0
xfeed_1094 0 1 tie_x0
xfeed_1095 0 1 tie_x0
xfeed_1096 0 1 tie_x0
xfeed_1097 0 1 tie_x0
xfeed_1098 0 1 tie_x0
xfeed_1099 0 1 tie_x0
xfeed_6022 0 1 tie_x0
xfeed_6021 0 1 tie_x0
xfeed_6020 0 1 tie_x0
xfeed_6029 0 1 tie_x0
xfeed_6028 0 1 tie_x0
xfeed_6027 0 1 tie_x0
xfeed_6026 0 1 tie_x0
xfeed_6025 0 1 tie_x0
xfeed_6024 0 1 tie_x0
xfeed_6023 0 1 tie_x0
xfeed_4889 0 1 tie_x0
xfeed_4888 0 1 tie_x0
xfeed_4887 0 1 tie_x0
xfeed_4886 0 1 tie_x0
xfeed_4885 0 1 tie_x0
xfeed_4884 0 1 tie_x0
xfeed_4883 0 1 tie_x0
xfeed_4882 0 1 tie_x0
xfeed_4881 0 1 tie_x0
xfeed_4880 0 1 tie_x0
xsubckt_9_oa2a22_x2 0 1 127 18 13 17 14 oa2a22_x2
xfeed_6039 0 1 tie_x0
xfeed_6038 0 1 tie_x0
xfeed_6037 0 1 tie_x0
xfeed_6036 0 1 tie_x0
xfeed_6035 0 1 tie_x0
xfeed_6034 0 1 tie_x0
xfeed_6033 0 1 tie_x0
xfeed_6032 0 1 tie_x0
xfeed_6031 0 1 tie_x0
xfeed_6030 0 1 tie_x0
xfeed_5509 0 1 tie_x0
xfeed_5508 0 1 tie_x0
xfeed_5507 0 1 tie_x0
xfeed_5506 0 1 tie_x0
xfeed_5505 0 1 tie_x0
xfeed_5504 0 1 tie_x0
xfeed_5503 0 1 tie_x0
xfeed_5502 0 1 tie_x0
xfeed_5501 0 1 tie_x0
xfeed_5500 0 1 tie_x0
xfeed_4899 0 1 tie_x0
xfeed_4898 0 1 tie_x0
xfeed_4897 0 1 tie_x0
xfeed_4896 0 1 tie_x0
xfeed_4895 0 1 tie_x0
xfeed_4894 0 1 tie_x0
xfeed_4893 0 1 tie_x0
xfeed_4892 0 1 tie_x0
xfeed_4891 0 1 tie_x0
xfeed_4890 0 1 tie_x0
xsubckt_44_ao22_x2 0 1 94 97 100 102 ao22_x2
xfeed_6049 0 1 tie_x0
xfeed_6048 0 1 tie_x0
xfeed_6047 0 1 tie_x0
xfeed_6046 0 1 tie_x0
xfeed_6045 0 1 tie_x0
xfeed_6044 0 1 tie_x0
xfeed_6043 0 1 tie_x0
xfeed_6042 0 1 tie_x0
xfeed_6041 0 1 tie_x0
xfeed_6040 0 1 tie_x0
xfeed_5519 0 1 tie_x0
xfeed_5518 0 1 tie_x0
xfeed_5517 0 1 tie_x0
xfeed_5516 0 1 tie_x0
xfeed_5515 0 1 tie_x0
xfeed_5514 0 1 tie_x0
xfeed_5513 0 1 tie_x0
xfeed_5512 0 1 tie_x0
xfeed_5511 0 1 tie_x0
xfeed_5510 0 1 tie_x0
xsubckt_133_ao22_x2 0 1 148 151 156 159 ao22_x2
xfeed_1200 0 1 tie_x0
xfeed_1201 0 1 tie_x0
xfeed_1202 0 1 tie_x0
xfeed_1203 0 1 tie_x0
xfeed_1204 0 1 tie_x0
xfeed_1205 0 1 tie_x0
xfeed_1206 0 1 tie_x0
xfeed_1207 0 1 tie_x0
xfeed_1208 0 1 tie_x0
xfeed_1209 0 1 tie_x0
xfeed_6059 0 1 tie_x0
xfeed_6058 0 1 tie_x0
xfeed_6057 0 1 tie_x0
xfeed_6056 0 1 tie_x0
xfeed_6055 0 1 tie_x0
xfeed_6054 0 1 tie_x0
xfeed_6053 0 1 tie_x0
xfeed_6052 0 1 tie_x0
xfeed_6051 0 1 tie_x0
xfeed_6050 0 1 tie_x0
xfeed_5529 0 1 tie_x0
xfeed_5528 0 1 tie_x0
xfeed_5527 0 1 tie_x0
xfeed_5526 0 1 tie_x0
xfeed_5525 0 1 tie_x0
xfeed_5524 0 1 tie_x0
xfeed_5523 0 1 tie_x0
xfeed_5522 0 1 tie_x0
xfeed_5521 0 1 tie_x0
xfeed_5520 0 1 tie_x0
xfeed_1210 0 1 tie_x0
xfeed_1211 0 1 tie_x0
xfeed_1212 0 1 tie_x0
xfeed_1213 0 1 tie_x0
xfeed_1214 0 1 tie_x0
xfeed_1215 0 1 tie_x0
xfeed_1216 0 1 tie_x0
xfeed_1217 0 1 tie_x0
xfeed_1218 0 1 tie_x0
xfeed_1219 0 1 tie_x0
xfeed_6069 0 1 tie_x0
xfeed_6068 0 1 tie_x0
xfeed_6067 0 1 tie_x0
xfeed_6066 0 1 tie_x0
xfeed_6065 0 1 tie_x0
xfeed_6064 0 1 tie_x0
xfeed_6063 0 1 tie_x0
xfeed_6062 0 1 tie_x0
xfeed_6061 0 1 tie_x0
xfeed_6060 0 1 tie_x0
xfeed_5539 0 1 tie_x0
xfeed_5538 0 1 tie_x0
xfeed_5537 0 1 tie_x0
xfeed_5536 0 1 tie_x0
xfeed_5535 0 1 tie_x0
xfeed_5534 0 1 tie_x0
xfeed_5533 0 1 tie_x0
xfeed_5532 0 1 tie_x0
xfeed_5531 0 1 tie_x0
xfeed_5530 0 1 tie_x0
xfeed_1220 0 1 tie_x0
xfeed_1221 0 1 tie_x0
xfeed_1222 0 1 tie_x0
xfeed_1223 0 1 tie_x0
xfeed_1224 0 1 tie_x0
xfeed_1225 0 1 tie_x0
xfeed_1226 0 1 tie_x0
xfeed_1227 0 1 tie_x0
xfeed_1228 0 1 tie_x0
xfeed_1229 0 1 tie_x0
xfeed_6079 0 1 tie_x0
xfeed_6078 0 1 tie_x0
xfeed_6077 0 1 tie_x0
xfeed_6076 0 1 tie_x0
xfeed_6075 0 1 tie_x0
xfeed_6074 0 1 tie_x0
xfeed_6073 0 1 tie_x0
xfeed_6072 0 1 tie_x0
xfeed_6071 0 1 tie_x0
xfeed_6070 0 1 tie_x0
xfeed_5549 0 1 tie_x0
xfeed_5548 0 1 tie_x0
xfeed_5547 0 1 tie_x0
xfeed_5546 0 1 tie_x0
xfeed_5545 0 1 tie_x0
xfeed_5544 0 1 tie_x0
xfeed_5543 0 1 tie_x0
xfeed_5542 0 1 tie_x0
xfeed_5541 0 1 tie_x0
xfeed_5540 0 1 tie_x0
xsubckt_138_nxr2_x1 0 1 143 75 4 nxr2_x1
xfeed_1230 0 1 tie_x0
xfeed_1231 0 1 tie_x0
xfeed_1232 0 1 tie_x0
xfeed_1233 0 1 tie_x0
xfeed_1234 0 1 tie_x0
xfeed_1235 0 1 tie_x0
xfeed_1236 0 1 tie_x0
xfeed_1237 0 1 tie_x0
xfeed_1238 0 1 tie_x0
xfeed_1239 0 1 tie_x0
xfeed_6089 0 1 tie_x0
xfeed_6088 0 1 tie_x0
xfeed_6087 0 1 tie_x0
xfeed_6086 0 1 tie_x0
xfeed_6085 0 1 tie_x0
xfeed_6084 0 1 tie_x0
xfeed_6083 0 1 tie_x0
xfeed_6082 0 1 tie_x0
xfeed_6081 0 1 tie_x0
xfeed_6080 0 1 tie_x0
xfeed_5559 0 1 tie_x0
xfeed_5558 0 1 tie_x0
xfeed_5557 0 1 tie_x0
xfeed_5556 0 1 tie_x0
xfeed_5555 0 1 tie_x0
xfeed_5554 0 1 rowend_x0
xfeed_5553 0 1 tie_x0
xfeed_5552 0 1 tie_x0
xfeed_5551 0 1 tie_x0
xfeed_5550 0 1 tie_x0
xfeed_1240 0 1 tie_x0
xfeed_1241 0 1 tie_x0
xfeed_1242 0 1 tie_x0
xfeed_1243 0 1 tie_x0
xfeed_1244 0 1 tie_x0
xfeed_1245 0 1 tie_x0
xfeed_1246 0 1 tie_x0
xfeed_1247 0 1 tie_x0
xfeed_1248 0 1 tie_x0
xfeed_1249 0 1 tie_x0
xfeed_6099 0 1 tie_x0
xfeed_6098 0 1 tie_x0
xfeed_6097 0 1 tie_x0
xfeed_6096 0 1 tie_x0
xfeed_6095 0 1 tie_x0
xfeed_6094 0 1 tie_x0
xfeed_6093 0 1 tie_x0
xfeed_6092 0 1 tie_x0
xfeed_6091 0 1 tie_x0
xfeed_6090 0 1 tie_x0
xfeed_5569 0 1 tie_x0
xfeed_5568 0 1 tie_x0
xfeed_5567 0 1 tie_x0
xfeed_5566 0 1 tie_x0
xfeed_5565 0 1 tie_x0
xfeed_5564 0 1 tie_x0
xfeed_5563 0 1 tie_x0
xfeed_5562 0 1 tie_x0
xfeed_5561 0 1 tie_x0
xfeed_5560 0 1 tie_x0
xfeed_1250 0 1 tie_x0
xfeed_1251 0 1 tie_x0
xfeed_1252 0 1 tie_x0
xfeed_1253 0 1 tie_x0
xfeed_1254 0 1 tie_x0
xfeed_1255 0 1 tie_x0
xfeed_1256 0 1 tie_x0
xfeed_1257 0 1 tie_x0
xfeed_1258 0 1 tie_x0
xfeed_1259 0 1 tie_x0
xfeed_5579 0 1 tie_x0
xfeed_5578 0 1 tie_x0
xfeed_5577 0 1 tie_x0
xfeed_5576 0 1 tie_x0
xfeed_5575 0 1 tie_x0
xfeed_5574 0 1 tie_x0
xfeed_5573 0 1 tie_x0
xfeed_5572 0 1 tie_x0
xfeed_5571 0 1 tie_x0
xfeed_5570 0 1 tie_x0
xfeed_1260 0 1 tie_x0
xfeed_1261 0 1 tie_x0
xfeed_1262 0 1 tie_x0
xfeed_1263 0 1 tie_x0
xfeed_1264 0 1 tie_x0
xfeed_1265 0 1 tie_x0
xfeed_1266 0 1 tie_x0
xfeed_1267 0 1 rowend_x0
xfeed_1268 0 1 tie_x0
xfeed_1269 0 1 tie_x0
xfeed_5589 0 1 tie_x0
xfeed_5588 0 1 tie_x0
xfeed_5587 0 1 tie_x0
xfeed_5586 0 1 tie_x0
xfeed_5585 0 1 tie_x0
xfeed_5584 0 1 tie_x0
xfeed_5583 0 1 tie_x0
xfeed_5582 0 1 tie_x0
xfeed_5581 0 1 tie_x0
xfeed_5580 0 1 tie_x0
xfeed_1270 0 1 tie_x0
xfeed_1271 0 1 tie_x0
xfeed_1272 0 1 tie_x0
xfeed_1273 0 1 tie_x0
xfeed_1274 0 1 tie_x0
xfeed_1275 0 1 tie_x0
xfeed_1276 0 1 tie_x0
xfeed_1277 0 1 tie_x0
xfeed_1278 0 1 tie_x0
xfeed_1279 0 1 tie_x0
xfeed_6209 0 1 tie_x0
xfeed_6208 0 1 tie_x0
xfeed_6207 0 1 tie_x0
xfeed_6206 0 1 tie_x0
xfeed_6205 0 1 tie_x0
xfeed_6204 0 1 tie_x0
xfeed_6203 0 1 tie_x0
xfeed_6202 0 1 tie_x0
xfeed_6201 0 1 tie_x0
xfeed_6200 0 1 tie_x0
xfeed_5599 0 1 tie_x0
xfeed_5598 0 1 tie_x0
xfeed_5597 0 1 tie_x0
xfeed_5596 0 1 tie_x0
xfeed_5595 0 1 tie_x0
xfeed_5594 0 1 tie_x0
xfeed_5593 0 1 tie_x0
xfeed_5592 0 1 tie_x0
xfeed_5591 0 1 tie_x0
xfeed_5590 0 1 tie_x0
xfeed_1280 0 1 tie_x0
xfeed_1281 0 1 tie_x0
xfeed_1282 0 1 tie_x0
xfeed_1283 0 1 tie_x0
xfeed_1284 0 1 tie_x0
xfeed_1285 0 1 tie_x0
xfeed_1286 0 1 tie_x0
xfeed_1287 0 1 rowend_x0
xfeed_1288 0 1 tie_x0
xfeed_1289 0 1 tie_x0
xsubckt_121_na2_x1 0 1 158 77 6 na2_x1
xfeed_6219 0 1 tie_x0
xfeed_6218 0 1 tie_x0
xfeed_6217 0 1 rowend_x0
xfeed_6216 0 1 tie_x0
xfeed_6215 0 1 tie_x0
xfeed_6214 0 1 tie_x0
xfeed_6213 0 1 tie_x0
xfeed_6212 0 1 tie_x0
xfeed_6211 0 1 tie_x0
xfeed_6210 0 1 tie_x0
xfeed_1290 0 1 tie_x0
xfeed_1291 0 1 tie_x0
xfeed_1292 0 1 tie_x0
xfeed_1293 0 1 tie_x0
xfeed_1294 0 1 tie_x0
xfeed_1295 0 1 tie_x0
xfeed_1296 0 1 tie_x0
xfeed_1297 0 1 tie_x0
xfeed_1298 0 1 tie_x0
xfeed_1299 0 1 tie_x0
xfeed_6229 0 1 tie_x0
xfeed_6228 0 1 tie_x0
xfeed_6227 0 1 tie_x0
xfeed_6226 0 1 tie_x0
xfeed_6225 0 1 tie_x0
xfeed_6224 0 1 tie_x0
xfeed_6223 0 1 tie_x0
xfeed_6222 0 1 tie_x0
xfeed_6221 0 1 tie_x0
xfeed_6220 0 1 tie_x0
xfeed_6239 0 1 tie_x0
xfeed_6238 0 1 tie_x0
xfeed_6237 0 1 tie_x0
xfeed_6236 0 1 tie_x0
xfeed_6235 0 1 tie_x0
xfeed_6234 0 1 tie_x0
xfeed_6233 0 1 tie_x0
xfeed_6232 0 1 tie_x0
xfeed_6231 0 1 tie_x0
xfeed_6230 0 1 tie_x0
xfeed_5709 0 1 rowend_x0
xfeed_5708 0 1 tie_x0
xfeed_5707 0 1 tie_x0
xfeed_5706 0 1 tie_x0
xfeed_5705 0 1 tie_x0
xfeed_5704 0 1 tie_x0
xfeed_5703 0 1 tie_x0
xfeed_5702 0 1 tie_x0
xfeed_5701 0 1 tie_x0
xfeed_5700 0 1 tie_x0
xsubckt_41_na2_x1 0 1 97 14 15 na2_x1
xfeed_6249 0 1 tie_x0
xfeed_6248 0 1 tie_x0
xfeed_6247 0 1 tie_x0
xfeed_6246 0 1 tie_x0
xfeed_6245 0 1 tie_x0
xfeed_6244 0 1 tie_x0
xfeed_6243 0 1 tie_x0
xfeed_6242 0 1 tie_x0
xfeed_6241 0 1 tie_x0
xfeed_6240 0 1 tie_x0
xfeed_5719 0 1 tie_x0
xfeed_5718 0 1 tie_x0
xfeed_5717 0 1 tie_x0
xfeed_5716 0 1 tie_x0
xfeed_5715 0 1 tie_x0
xfeed_5714 0 1 tie_x0
xfeed_5713 0 1 tie_x0
xfeed_5712 0 1 tie_x0
xfeed_5711 0 1 tie_x0
xfeed_5710 0 1 tie_x0
xfeed_1400 0 1 tie_x0
xfeed_1401 0 1 tie_x0
xfeed_1402 0 1 tie_x0
xfeed_1403 0 1 tie_x0
xfeed_1404 0 1 tie_x0
xfeed_1405 0 1 tie_x0
xfeed_1406 0 1 tie_x0
xfeed_1407 0 1 tie_x0
xfeed_1408 0 1 tie_x0
xfeed_1409 0 1 tie_x0
xsubckt_152_sff1_x4 0 1 6 225 40 sff1_x4
xfeed_6259 0 1 tie_x0
xfeed_6258 0 1 tie_x0
xfeed_6257 0 1 tie_x0
xfeed_6256 0 1 tie_x0
xfeed_6255 0 1 tie_x0
xfeed_6254 0 1 tie_x0
xfeed_6253 0 1 tie_x0
xfeed_6252 0 1 tie_x0
xfeed_6251 0 1 tie_x0
xfeed_6250 0 1 tie_x0
xfeed_5729 0 1 tie_x0
xfeed_5728 0 1 tie_x0
xfeed_5727 0 1 tie_x0
xfeed_5726 0 1 tie_x0
xfeed_5725 0 1 tie_x0
xfeed_5724 0 1 tie_x0
xfeed_5723 0 1 tie_x0
xfeed_5722 0 1 tie_x0
xfeed_5721 0 1 tie_x0
xfeed_5720 0 1 tie_x0
xfeed_1410 0 1 tie_x0
xfeed_1411 0 1 tie_x0
xfeed_1412 0 1 tie_x0
xfeed_1413 0 1 tie_x0
xfeed_1414 0 1 tie_x0
xfeed_1415 0 1 tie_x0
xfeed_1416 0 1 tie_x0
xfeed_1417 0 1 tie_x0
xfeed_1418 0 1 tie_x0
xfeed_1419 0 1 tie_x0
xsubckt_101_xr2_x4 0 1 175 80 9 xr2_x4
xsubckt_148_sff1_x4 0 1 10 229 40 sff1_x4
xfeed_6269 0 1 tie_x0
xfeed_6268 0 1 tie_x0
xfeed_6267 0 1 tie_x0
xfeed_6266 0 1 tie_x0
xfeed_6265 0 1 tie_x0
xfeed_6264 0 1 tie_x0
xfeed_6263 0 1 tie_x0
xfeed_6262 0 1 tie_x0
xfeed_6261 0 1 tie_x0
xfeed_6260 0 1 tie_x0
xfeed_5739 0 1 tie_x0
xfeed_5738 0 1 tie_x0
xfeed_5737 0 1 tie_x0
xfeed_5736 0 1 tie_x0
xfeed_5735 0 1 tie_x0
xfeed_5734 0 1 tie_x0
xfeed_5733 0 1 tie_x0
xfeed_5732 0 1 tie_x0
xfeed_5731 0 1 tie_x0
xfeed_5730 0 1 tie_x0
xsubckt_107_xr2_x4 0 1 170 79 8 xr2_x4
xfeed_1420 0 1 tie_x0
xfeed_1421 0 1 tie_x0
xfeed_1422 0 1 tie_x0
xfeed_1423 0 1 tie_x0
xfeed_1424 0 1 tie_x0
xfeed_1425 0 1 tie_x0
xfeed_1426 0 1 tie_x0
xfeed_1427 0 1 tie_x0
xfeed_1428 0 1 tie_x0
xfeed_1429 0 1 tie_x0
xfeed_6279 0 1 tie_x0
xfeed_6278 0 1 tie_x0
xfeed_6277 0 1 tie_x0
xfeed_6276 0 1 tie_x0
xfeed_6275 0 1 tie_x0
xfeed_6274 0 1 tie_x0
xfeed_6273 0 1 tie_x0
xfeed_6272 0 1 tie_x0
xfeed_6271 0 1 tie_x0
xfeed_6270 0 1 tie_x0
xfeed_5749 0 1 tie_x0
xfeed_5748 0 1 tie_x0
xfeed_5747 0 1 tie_x0
xfeed_5746 0 1 tie_x0
xfeed_5745 0 1 tie_x0
xfeed_5744 0 1 tie_x0
xfeed_5743 0 1 tie_x0
xfeed_5742 0 1 tie_x0
xfeed_5741 0 1 tie_x0
xfeed_5740 0 1 tie_x0
xfeed_1430 0 1 tie_x0
xfeed_1431 0 1 tie_x0
xfeed_1432 0 1 tie_x0
xfeed_1433 0 1 tie_x0
xfeed_1434 0 1 tie_x0
xfeed_1435 0 1 tie_x0
xfeed_1436 0 1 tie_x0
xfeed_1437 0 1 tie_x0
xfeed_1438 0 1 tie_x0
xfeed_1439 0 1 tie_x0
xsubckt_26_noa2a22_x1 0 1 112 17 12 11 18 noa2a22_x1
xfeed_6289 0 1 tie_x0
xfeed_6288 0 1 tie_x0
xfeed_6287 0 1 tie_x0
xfeed_6286 0 1 tie_x0
xfeed_6285 0 1 tie_x0
xfeed_6284 0 1 tie_x0
xfeed_6283 0 1 tie_x0
xfeed_6282 0 1 tie_x0
xfeed_6281 0 1 tie_x0
xfeed_6280 0 1 tie_x0
xfeed_5759 0 1 tie_x0
xfeed_5758 0 1 tie_x0
xfeed_5757 0 1 tie_x0
xfeed_5756 0 1 rowend_x0
xfeed_5755 0 1 tie_x0
xfeed_5754 0 1 tie_x0
xfeed_5753 0 1 tie_x0
xfeed_5752 0 1 tie_x0
xfeed_5751 0 1 tie_x0
xfeed_5750 0 1 tie_x0
xfeed_1440 0 1 tie_x0
xfeed_1441 0 1 tie_x0
xfeed_1442 0 1 tie_x0
xfeed_1443 0 1 tie_x0
xfeed_1444 0 1 tie_x0
xfeed_1445 0 1 tie_x0
xfeed_1446 0 1 tie_x0
xfeed_1447 0 1 tie_x0
xfeed_1448 0 1 tie_x0
xfeed_1449 0 1 tie_x0
xfeed_6299 0 1 tie_x0
xfeed_6298 0 1 tie_x0
xfeed_6297 0 1 tie_x0
xfeed_6296 0 1 tie_x0
xfeed_6295 0 1 tie_x0
xfeed_6294 0 1 tie_x0
xfeed_6293 0 1 tie_x0
xfeed_6292 0 1 tie_x0
xfeed_6291 0 1 tie_x0
xfeed_6290 0 1 tie_x0
xfeed_5769 0 1 tie_x0
xfeed_5768 0 1 tie_x0
xfeed_5767 0 1 tie_x0
xfeed_5766 0 1 tie_x0
xfeed_5765 0 1 tie_x0
xfeed_5764 0 1 tie_x0
xfeed_5763 0 1 tie_x0
xfeed_5762 0 1 tie_x0
xfeed_5761 0 1 tie_x0
xfeed_5760 0 1 tie_x0
xfeed_1450 0 1 tie_x0
xfeed_1451 0 1 tie_x0
xfeed_1452 0 1 tie_x0
xfeed_1453 0 1 tie_x0
xfeed_1454 0 1 tie_x0
xfeed_1455 0 1 tie_x0
xfeed_1456 0 1 tie_x0
xfeed_1457 0 1 tie_x0
xfeed_1458 0 1 tie_x0
xfeed_1459 0 1 tie_x0
xfeed_5779 0 1 tie_x0
xfeed_5778 0 1 tie_x0
xfeed_5777 0 1 tie_x0
xfeed_5776 0 1 tie_x0
xfeed_5775 0 1 tie_x0
xfeed_5774 0 1 tie_x0
xfeed_5773 0 1 tie_x0
xfeed_5772 0 1 tie_x0
xfeed_5771 0 1 tie_x0
xfeed_5770 0 1 tie_x0
xsubckt_6_mx2_x2 0 1 229 10 130 2 mx2_x2
xfeed_1460 0 1 tie_x0
xfeed_1461 0 1 tie_x0
xfeed_1462 0 1 tie_x0
xfeed_1463 0 1 tie_x0
xfeed_1464 0 1 tie_x0
xfeed_1465 0 1 tie_x0
xfeed_1466 0 1 tie_x0
xfeed_1467 0 1 tie_x0
xfeed_1468 0 1 tie_x0
xfeed_1469 0 1 tie_x0
xfeed_5789 0 1 tie_x0
xfeed_5788 0 1 tie_x0
xfeed_5787 0 1 tie_x0
xfeed_5786 0 1 tie_x0
xfeed_5785 0 1 tie_x0
xfeed_5784 0 1 tie_x0
xfeed_5783 0 1 rowend_x0
xfeed_5782 0 1 tie_x0
xfeed_5781 0 1 tie_x0
xfeed_5780 0 1 tie_x0
xsubckt_78_a2_x2 0 1 194 211 195 a2_x2
xsubckt_98_a2_x2 0 1 221 131 178 a2_x2
xfeed_1470 0 1 tie_x0
xfeed_1471 0 1 tie_x0
xfeed_1472 0 1 tie_x0
xfeed_1473 0 1 tie_x0
xfeed_1474 0 1 tie_x0
xfeed_1475 0 1 tie_x0
xfeed_1476 0 1 tie_x0
xfeed_1477 0 1 tie_x0
xfeed_1478 0 1 tie_x0
xfeed_1479 0 1 tie_x0
xsubckt_16_noa2a22_x1 0 1 121 13 17 12 18 noa2a22_x1
xfeed_6409 0 1 tie_x0
xfeed_6408 0 1 tie_x0
xfeed_6407 0 1 tie_x0
xfeed_6406 0 1 tie_x0
xfeed_6405 0 1 tie_x0
xfeed_6404 0 1 tie_x0
xfeed_6403 0 1 tie_x0
xfeed_6402 0 1 tie_x0
xfeed_6401 0 1 tie_x0
xfeed_6400 0 1 rowend_x0
xfeed_5799 0 1 tie_x0
xfeed_5798 0 1 tie_x0
xfeed_5797 0 1 tie_x0
xfeed_5796 0 1 tie_x0
xfeed_5795 0 1 tie_x0
xfeed_5794 0 1 tie_x0
xfeed_5793 0 1 tie_x0
xfeed_5792 0 1 tie_x0
xfeed_5791 0 1 tie_x0
xfeed_5790 0 1 tie_x0
xsubckt_136_na2_x1 0 1 145 75 4 na2_x1
xfeed_1480 0 1 tie_x0
xfeed_1481 0 1 tie_x0
xfeed_1482 0 1 tie_x0
xfeed_1483 0 1 tie_x0
xfeed_1484 0 1 tie_x0
xfeed_1485 0 1 tie_x0
xfeed_1486 0 1 tie_x0
xfeed_1487 0 1 tie_x0
xfeed_1488 0 1 tie_x0
xfeed_1489 0 1 tie_x0
xfeed_6419 0 1 tie_x0
xfeed_6418 0 1 tie_x0
xfeed_6417 0 1 tie_x0
xfeed_6416 0 1 tie_x0
xfeed_6415 0 1 tie_x0
xfeed_6414 0 1 tie_x0
xfeed_6413 0 1 tie_x0
xfeed_6412 0 1 tie_x0
xfeed_6411 0 1 tie_x0
xfeed_6410 0 1 tie_x0
xfeed_2109 0 1 tie_x0
xfeed_2108 0 1 tie_x0
xfeed_2107 0 1 tie_x0
xfeed_2106 0 1 tie_x0
xfeed_2105 0 1 tie_x0
xfeed_1490 0 1 tie_x0
xfeed_1491 0 1 tie_x0
xfeed_1492 0 1 tie_x0
xfeed_1493 0 1 tie_x0
xfeed_1494 0 1 tie_x0
xfeed_1495 0 1 tie_x0
xfeed_1496 0 1 tie_x0
xfeed_1497 0 1 tie_x0
xfeed_1498 0 1 tie_x0
xfeed_1499 0 1 tie_x0
xfeed_2100 0 1 tie_x0
xfeed_2101 0 1 tie_x0
xfeed_2102 0 1 tie_x0
xfeed_2103 0 1 tie_x0
xfeed_2104 0 1 tie_x0
xfeed_6429 0 1 tie_x0
xfeed_6428 0 1 tie_x0
xfeed_6427 0 1 rowend_x0
xfeed_6426 0 1 tie_x0
xfeed_6425 0 1 tie_x0
xfeed_6424 0 1 tie_x0
xfeed_6423 0 1 tie_x0
xfeed_6422 0 1 tie_x0
xfeed_6421 0 1 tie_x0
xfeed_6420 0 1 tie_x0
xfeed_2119 0 1 tie_x0
xfeed_2118 0 1 tie_x0
xfeed_2117 0 1 tie_x0
xfeed_2116 0 1 tie_x0
xfeed_2115 0 1 tie_x0
xfeed_2114 0 1 tie_x0
xfeed_2113 0 1 tie_x0
xfeed_2112 0 1 tie_x0
xfeed_2111 0 1 tie_x0
xfeed_2110 0 1 tie_x0
xfeed_6439 0 1 tie_x0
xfeed_6438 0 1 tie_x0
xfeed_6437 0 1 tie_x0
xfeed_6436 0 1 tie_x0
xfeed_6435 0 1 tie_x0
xfeed_6434 0 1 tie_x0
xfeed_6433 0 1 tie_x0
xfeed_6432 0 1 tie_x0
xfeed_6431 0 1 tie_x0
xfeed_6430 0 1 tie_x0
xfeed_5909 0 1 tie_x0
xfeed_5908 0 1 tie_x0
xfeed_5907 0 1 tie_x0
xfeed_5906 0 1 tie_x0
xfeed_5905 0 1 tie_x0
xfeed_5904 0 1 tie_x0
xfeed_5903 0 1 tie_x0
xfeed_5902 0 1 tie_x0
xfeed_5901 0 1 tie_x0
xfeed_5900 0 1 tie_x0
xfeed_2129 0 1 tie_x0
xfeed_2128 0 1 tie_x0
xfeed_2127 0 1 tie_x0
xfeed_2126 0 1 rowend_x0
xfeed_2125 0 1 tie_x0
xfeed_2124 0 1 tie_x0
xfeed_2123 0 1 tie_x0
xfeed_2122 0 1 tie_x0
xfeed_2121 0 1 tie_x0
xfeed_2120 0 1 tie_x0
xsubckt_54_na2_x1 0 1 85 13 15 na2_x1
xsubckt_58_na2_x1 0 1 213 12 16 na2_x1
xfeed_100 0 1 tie_x0
xfeed_101 0 1 tie_x0
xfeed_102 0 1 tie_x0
xfeed_103 0 1 tie_x0
xfeed_104 0 1 tie_x0
xfeed_105 0 1 tie_x0
xfeed_106 0 1 tie_x0
xfeed_107 0 1 tie_x0
xfeed_108 0 1 tie_x0
xfeed_109 0 1 tie_x0
xfeed_6449 0 1 tie_x0
xfeed_6448 0 1 tie_x0
xfeed_6447 0 1 tie_x0
xfeed_6446 0 1 tie_x0
xfeed_6445 0 1 tie_x0
xfeed_6444 0 1 tie_x0
xfeed_6443 0 1 tie_x0
xfeed_6442 0 1 tie_x0
xfeed_6441 0 1 tie_x0
xfeed_6440 0 1 tie_x0
xfeed_5919 0 1 tie_x0
xfeed_5918 0 1 tie_x0
xfeed_5917 0 1 tie_x0
xfeed_5916 0 1 tie_x0
xfeed_5915 0 1 tie_x0
xfeed_5914 0 1 tie_x0
xfeed_5913 0 1 tie_x0
xfeed_5912 0 1 tie_x0
xfeed_5911 0 1 tie_x0
xfeed_5910 0 1 tie_x0
xfeed_2139 0 1 tie_x0
xfeed_2138 0 1 tie_x0
xfeed_2137 0 1 tie_x0
xfeed_2136 0 1 tie_x0
xfeed_2135 0 1 tie_x0
xfeed_2134 0 1 tie_x0
xfeed_2133 0 1 tie_x0
xfeed_2132 0 1 tie_x0
xfeed_2131 0 1 tie_x0
xfeed_2130 0 1 tie_x0
xfeed_1600 0 1 tie_x0
xfeed_1601 0 1 tie_x0
xfeed_1602 0 1 tie_x0
xfeed_1603 0 1 tie_x0
xfeed_1604 0 1 tie_x0
xfeed_1605 0 1 tie_x0
xfeed_1606 0 1 tie_x0
xfeed_1607 0 1 tie_x0
xfeed_1608 0 1 tie_x0
xfeed_1609 0 1 tie_x0
xfeed_110 0 1 tie_x0
xfeed_111 0 1 tie_x0
xfeed_112 0 1 tie_x0
xfeed_113 0 1 tie_x0
xfeed_114 0 1 tie_x0
xfeed_115 0 1 tie_x0
xfeed_116 0 1 tie_x0
xfeed_117 0 1 tie_x0
xfeed_118 0 1 tie_x0
xfeed_119 0 1 tie_x0
xfeed_6459 0 1 tie_x0
xfeed_6458 0 1 tie_x0
xfeed_6457 0 1 tie_x0
xfeed_6456 0 1 tie_x0
xfeed_6455 0 1 tie_x0
xfeed_6454 0 1 tie_x0
xfeed_6453 0 1 tie_x0
xfeed_6452 0 1 tie_x0
xfeed_6451 0 1 tie_x0
xfeed_6450 0 1 tie_x0
xfeed_5929 0 1 tie_x0
xfeed_5928 0 1 tie_x0
xfeed_5927 0 1 tie_x0
xfeed_5926 0 1 tie_x0
xfeed_5925 0 1 tie_x0
xfeed_5924 0 1 tie_x0
xfeed_5923 0 1 tie_x0
xfeed_5922 0 1 tie_x0
xfeed_5921 0 1 tie_x0
xfeed_5920 0 1 tie_x0
xfeed_2149 0 1 tie_x0
xfeed_2148 0 1 tie_x0
xfeed_2147 0 1 tie_x0
xfeed_2146 0 1 tie_x0
xfeed_2145 0 1 tie_x0
xfeed_2144 0 1 tie_x0
xfeed_2143 0 1 tie_x0
xfeed_2142 0 1 tie_x0
xfeed_2141 0 1 tie_x0
xfeed_2140 0 1 tie_x0
xsubckt_114_xr2_x4 0 1 164 78 7 xr2_x4
xsubckt_144_nxr2_x1 0 1 138 74 3 nxr2_x1
xfeed_1610 0 1 tie_x0
xfeed_1611 0 1 tie_x0
xfeed_1612 0 1 tie_x0
xfeed_1613 0 1 tie_x0
xfeed_1614 0 1 tie_x0
xfeed_1615 0 1 tie_x0
xfeed_1616 0 1 tie_x0
xfeed_1617 0 1 tie_x0
xfeed_1618 0 1 tie_x0
xfeed_1619 0 1 tie_x0
xfeed_120 0 1 tie_x0
xfeed_121 0 1 tie_x0
xfeed_122 0 1 tie_x0
xfeed_123 0 1 tie_x0
xfeed_124 0 1 tie_x0
xfeed_125 0 1 tie_x0
xfeed_126 0 1 tie_x0
xfeed_127 0 1 tie_x0
xfeed_128 0 1 tie_x0
xfeed_129 0 1 tie_x0
xfeed_6469 0 1 tie_x0
xfeed_6468 0 1 tie_x0
xfeed_6467 0 1 tie_x0
xfeed_6466 0 1 tie_x0
xfeed_6465 0 1 tie_x0
xfeed_6464 0 1 tie_x0
xfeed_6463 0 1 tie_x0
xfeed_6462 0 1 tie_x0
xfeed_6461 0 1 tie_x0
xfeed_6460 0 1 tie_x0
xfeed_5939 0 1 tie_x0
xfeed_5938 0 1 tie_x0
xfeed_5937 0 1 tie_x0
xfeed_5936 0 1 tie_x0
xfeed_5935 0 1 tie_x0
xfeed_5934 0 1 tie_x0
xfeed_5933 0 1 tie_x0
xfeed_5932 0 1 tie_x0
xfeed_5931 0 1 tie_x0
xfeed_5930 0 1 tie_x0
xfeed_2159 0 1 tie_x0
xfeed_2158 0 1 tie_x0
xfeed_2157 0 1 tie_x0
xfeed_2156 0 1 tie_x0
xfeed_2155 0 1 tie_x0
xfeed_2154 0 1 tie_x0
xfeed_2153 0 1 tie_x0
xfeed_2152 0 1 tie_x0
xfeed_2151 0 1 tie_x0
xfeed_2150 0 1 tie_x0
xfeed_1620 0 1 tie_x0
xfeed_1621 0 1 tie_x0
xfeed_1622 0 1 tie_x0
xfeed_1623 0 1 tie_x0
xfeed_1624 0 1 tie_x0
xfeed_1625 0 1 tie_x0
xfeed_1626 0 1 tie_x0
xfeed_1627 0 1 tie_x0
xfeed_1628 0 1 tie_x0
xfeed_1629 0 1 tie_x0
xfeed_130 0 1 rowend_x0
xfeed_131 0 1 tie_x0
xfeed_132 0 1 tie_x0
xfeed_133 0 1 tie_x0
xfeed_134 0 1 tie_x0
xfeed_135 0 1 tie_x0
xfeed_136 0 1 tie_x0
xfeed_137 0 1 tie_x0
xfeed_138 0 1 tie_x0
xfeed_139 0 1 tie_x0
xfeed_6479 0 1 tie_x0
xfeed_6478 0 1 rowend_x0
xfeed_6477 0 1 tie_x0
xfeed_6476 0 1 tie_x0
xfeed_6475 0 1 tie_x0
xfeed_6474 0 1 tie_x0
xfeed_6473 0 1 tie_x0
xfeed_6472 0 1 tie_x0
xfeed_6471 0 1 tie_x0
xfeed_6470 0 1 tie_x0
xfeed_5946 0 1 tie_x0
xfeed_5945 0 1 tie_x0
xfeed_5944 0 1 tie_x0
xfeed_5943 0 1 tie_x0
xfeed_5942 0 1 tie_x0
xfeed_5941 0 1 tie_x0
xfeed_5940 0 1 tie_x0
xfeed_2169 0 1 tie_x0
xfeed_2168 0 1 tie_x0
xfeed_2167 0 1 tie_x0
xfeed_2166 0 1 tie_x0
xfeed_2165 0 1 tie_x0
xfeed_2164 0 1 tie_x0
xfeed_2163 0 1 tie_x0
xfeed_2162 0 1 tie_x0
xfeed_2161 0 1 tie_x0
xfeed_2160 0 1 tie_x0
xfeed_1630 0 1 tie_x0
xfeed_1631 0 1 tie_x0
xfeed_1632 0 1 tie_x0
xfeed_1633 0 1 tie_x0
xfeed_1634 0 1 tie_x0
xfeed_1635 0 1 tie_x0
xfeed_1636 0 1 tie_x0
xfeed_1637 0 1 tie_x0
xfeed_1638 0 1 tie_x0
xfeed_1639 0 1 tie_x0
xfeed_5949 0 1 tie_x0
xfeed_5948 0 1 tie_x0
xfeed_5947 0 1 tie_x0
xfeed_140 0 1 tie_x0
xfeed_141 0 1 tie_x0
xfeed_142 0 1 tie_x0
xfeed_143 0 1 tie_x0
xfeed_144 0 1 tie_x0
xfeed_145 0 1 tie_x0
xfeed_146 0 1 tie_x0
xfeed_147 0 1 tie_x0
xfeed_148 0 1 tie_x0
xfeed_149 0 1 tie_x0
xfeed_6489 0 1 tie_x0
xfeed_6488 0 1 tie_x0
xfeed_6487 0 1 tie_x0
xfeed_6486 0 1 tie_x0
xfeed_6485 0 1 tie_x0
xfeed_6484 0 1 tie_x0
xfeed_6483 0 1 tie_x0
xfeed_6482 0 1 tie_x0
xfeed_6481 0 1 tie_x0
xfeed_6480 0 1 tie_x0
xfeed_5953 0 1 tie_x0
xfeed_5952 0 1 tie_x0
xfeed_5951 0 1 tie_x0
xfeed_5950 0 1 tie_x0
xfeed_2179 0 1 tie_x0
xfeed_2178 0 1 tie_x0
xfeed_2177 0 1 tie_x0
xfeed_2176 0 1 tie_x0
xfeed_2175 0 1 tie_x0
xfeed_2174 0 1 tie_x0
xfeed_2173 0 1 tie_x0
xfeed_2172 0 1 tie_x0
xfeed_2171 0 1 tie_x0
xfeed_2170 0 1 tie_x0
xsubckt_33_na3_x1 0 1 105 111 109 108 na3_x1
xsubckt_37_na3_x1 0 1 101 113 105 103 na3_x1
xfeed_1640 0 1 tie_x0
xfeed_1641 0 1 tie_x0
xfeed_1642 0 1 tie_x0
xfeed_1643 0 1 tie_x0
xfeed_1644 0 1 tie_x0
xfeed_1645 0 1 tie_x0
xfeed_1646 0 1 tie_x0
xfeed_1647 0 1 tie_x0
xfeed_1648 0 1 tie_x0
xfeed_1649 0 1 tie_x0
xfeed_5959 0 1 tie_x0
xfeed_5958 0 1 tie_x0
xfeed_5957 0 1 tie_x0
xfeed_5956 0 1 tie_x0
xfeed_5955 0 1 tie_x0
xfeed_5954 0 1 tie_x0
xfeed_150 0 1 tie_x0
xfeed_151 0 1 tie_x0
xfeed_152 0 1 tie_x0
xfeed_153 0 1 tie_x0
xfeed_154 0 1 tie_x0
xfeed_155 0 1 tie_x0
xfeed_156 0 1 tie_x0
xfeed_157 0 1 tie_x0
xfeed_158 0 1 tie_x0
xfeed_159 0 1 tie_x0
xfeed_7109 0 1 tie_x0
xfeed_7108 0 1 tie_x0
xfeed_7107 0 1 tie_x0
xfeed_7106 0 1 tie_x0
xfeed_7105 0 1 tie_x0
xfeed_7104 0 1 tie_x0
xfeed_7103 0 1 tie_x0
xfeed_7102 0 1 tie_x0
xfeed_7101 0 1 tie_x0
xfeed_7100 0 1 tie_x0
xfeed_6499 0 1 tie_x0
xfeed_6498 0 1 tie_x0
xfeed_6497 0 1 tie_x0
xfeed_6496 0 1 tie_x0
xfeed_6495 0 1 tie_x0
xfeed_6494 0 1 tie_x0
xfeed_6493 0 1 tie_x0
xfeed_6492 0 1 tie_x0
xfeed_6491 0 1 tie_x0
xfeed_6490 0 1 tie_x0
xfeed_5960 0 1 tie_x0
xfeed_2189 0 1 tie_x0
xfeed_2188 0 1 tie_x0
xfeed_2187 0 1 tie_x0
xfeed_2186 0 1 tie_x0
xfeed_2185 0 1 tie_x0
xfeed_2184 0 1 tie_x0
xfeed_2183 0 1 tie_x0
xfeed_2182 0 1 tie_x0
xfeed_2181 0 1 tie_x0
xfeed_2180 0 1 tie_x0
xsubckt_8_na4_x1 0 1 128 18 14 13 17 na4_x1
xfeed_1650 0 1 tie_x0
xfeed_1651 0 1 tie_x0
xfeed_1652 0 1 tie_x0
xfeed_1653 0 1 tie_x0
xfeed_1654 0 1 tie_x0
xfeed_1655 0 1 tie_x0
xfeed_1656 0 1 tie_x0
xfeed_1657 0 1 tie_x0
xfeed_1658 0 1 tie_x0
xfeed_1659 0 1 tie_x0
xfeed_5969 0 1 tie_x0
xfeed_5968 0 1 tie_x0
xfeed_5967 0 1 tie_x0
xfeed_5966 0 1 tie_x0
xfeed_5965 0 1 tie_x0
xfeed_5964 0 1 tie_x0
xfeed_5963 0 1 tie_x0
xfeed_5962 0 1 tie_x0
xfeed_5961 0 1 rowend_x0
xfeed_160 0 1 tie_x0
xfeed_161 0 1 tie_x0
xfeed_162 0 1 tie_x0
xfeed_163 0 1 tie_x0
xfeed_164 0 1 tie_x0
xfeed_165 0 1 tie_x0
xfeed_166 0 1 tie_x0
xfeed_167 0 1 tie_x0
xfeed_168 0 1 tie_x0
xfeed_169 0 1 tie_x0
xfeed_7119 0 1 tie_x0
xfeed_7118 0 1 tie_x0
xfeed_7117 0 1 tie_x0
xfeed_7116 0 1 tie_x0
xfeed_7115 0 1 tie_x0
xfeed_7114 0 1 tie_x0
xfeed_7113 0 1 tie_x0
xfeed_7112 0 1 tie_x0
xfeed_7111 0 1 tie_x0
xfeed_7110 0 1 tie_x0
xfeed_2199 0 1 tie_x0
xfeed_2198 0 1 tie_x0
xfeed_2197 0 1 tie_x0
xfeed_2196 0 1 tie_x0
xfeed_2195 0 1 tie_x0
xfeed_2194 0 1 tie_x0
xfeed_2193 0 1 tie_x0
xfeed_2192 0 1 tie_x0
xfeed_2191 0 1 tie_x0
xfeed_2190 0 1 tie_x0
xsubckt_53_nao22_x1 0 1 86 101 100 97 nao22_x1
xspare_feed_200 0 1 rowend_x0
xspare_feed_201 0 1 tie_x0
xspare_feed_202 0 1 rowend_x0
xspare_feed_203 0 1 rowend_x0
xspare_feed_204 0 1 tie_x0
xspare_feed_205 0 1 rowend_x0
xspare_feed_206 0 1 tie_x0
xspare_feed_207 0 1 rowend_x0
xspare_feed_208 0 1 rowend_x0
xspare_feed_209 0 1 tie_x0
xfeed_1660 0 1 tie_x0
xfeed_1661 0 1 tie_x0
xfeed_1662 0 1 tie_x0
xfeed_1663 0 1 tie_x0
xfeed_1664 0 1 tie_x0
xfeed_1665 0 1 tie_x0
xfeed_1666 0 1 tie_x0
xfeed_1667 0 1 tie_x0
xfeed_5979 0 1 tie_x0
xfeed_5978 0 1 tie_x0
xfeed_5977 0 1 tie_x0
xfeed_5976 0 1 tie_x0
xfeed_5975 0 1 tie_x0
xfeed_5974 0 1 tie_x0
xfeed_5973 0 1 tie_x0
xfeed_5972 0 1 tie_x0
xfeed_5971 0 1 tie_x0
xfeed_5970 0 1 tie_x0
xsubckt_7_a4_x2 0 1 129 18 14 13 17 a4_x2
xfeed_170 0 1 tie_x0
xfeed_171 0 1 tie_x0
xfeed_172 0 1 tie_x0
xfeed_173 0 1 tie_x0
xfeed_174 0 1 tie_x0
xfeed_175 0 1 tie_x0
xfeed_176 0 1 tie_x0
xfeed_177 0 1 tie_x0
xfeed_178 0 1 tie_x0
xfeed_179 0 1 tie_x0
xfeed_1668 0 1 tie_x0
xfeed_1669 0 1 tie_x0
xfeed_7129 0 1 tie_x0
xfeed_7128 0 1 tie_x0
xfeed_7127 0 1 tie_x0
xfeed_7126 0 1 tie_x0
xfeed_7125 0 1 tie_x0
xfeed_7124 0 1 tie_x0
xfeed_7123 0 1 tie_x0
xfeed_7122 0 1 tie_x0
xfeed_7121 0 1 tie_x0
xfeed_7120 0 1 tie_x0
xspare_feed_210 0 1 rowend_x0
xspare_feed_211 0 1 tie_x0
xspare_feed_212 0 1 rowend_x0
xspare_feed_213 0 1 rowend_x0
xspare_feed_214 0 1 tie_x0
xspare_feed_215 0 1 rowend_x0
xspare_feed_216 0 1 tie_x0
xspare_feed_217 0 1 rowend_x0
xspare_feed_218 0 1 rowend_x0
xspare_feed_219 0 1 tie_x0
xfeed_1670 0 1 tie_x0
xfeed_1671 0 1 tie_x0
xfeed_1672 0 1 tie_x0
xfeed_1673 0 1 tie_x0
xfeed_1674 0 1 tie_x0
xfeed_5989 0 1 tie_x0
xfeed_5988 0 1 tie_x0
xfeed_5987 0 1 tie_x0
xfeed_5986 0 1 rowend_x0
xfeed_5985 0 1 tie_x0
xfeed_5984 0 1 tie_x0
xfeed_5983 0 1 tie_x0
xfeed_5982 0 1 tie_x0
xfeed_5981 0 1 tie_x0
xfeed_5980 0 1 tie_x0
xfeed_189 0 1 tie_x0
xfeed_188 0 1 tie_x0
xfeed_187 0 1 tie_x0
xfeed_186 0 1 tie_x0
xfeed_185 0 1 tie_x0
xfeed_180 0 1 tie_x0
xfeed_181 0 1 tie_x0
xfeed_182 0 1 tie_x0
xfeed_183 0 1 tie_x0
xfeed_184 0 1 tie_x0
xfeed_1675 0 1 tie_x0
xfeed_1676 0 1 rowend_x0
xfeed_1677 0 1 tie_x0
xfeed_1678 0 1 tie_x0
xfeed_1679 0 1 tie_x0
xfeed_7139 0 1 tie_x0
xfeed_7138 0 1 tie_x0
xfeed_7137 0 1 tie_x0
xfeed_7136 0 1 tie_x0
xfeed_7135 0 1 tie_x0
xfeed_7134 0 1 tie_x0
xfeed_7133 0 1 tie_x0
xfeed_7132 0 1 tie_x0
xfeed_7131 0 1 tie_x0
xfeed_7130 0 1 tie_x0
xfeed_6609 0 1 tie_x0
xfeed_6608 0 1 tie_x0
xfeed_6607 0 1 tie_x0
xfeed_6606 0 1 tie_x0
xfeed_6605 0 1 tie_x0
xfeed_6604 0 1 tie_x0
xfeed_6603 0 1 tie_x0
xfeed_6602 0 1 tie_x0
xfeed_6601 0 1 tie_x0
xfeed_6600 0 1 tie_x0
xspare_feed_220 0 1 rowend_x0
xspare_feed_221 0 1 tie_x0
xspare_feed_222 0 1 rowend_x0
xspare_feed_223 0 1 rowend_x0
xspare_feed_224 0 1 tie_x0
xspare_feed_225 0 1 rowend_x0
xspare_feed_226 0 1 tie_x0
xspare_feed_227 0 1 rowend_x0
xspare_feed_228 0 1 rowend_x0
xspare_feed_229 0 1 tie_x0
xfeed_1680 0 1 tie_x0
xfeed_1681 0 1 tie_x0
xfeed_5999 0 1 tie_x0
xfeed_5998 0 1 tie_x0
xfeed_5997 0 1 tie_x0
xfeed_5996 0 1 tie_x0
xfeed_5995 0 1 tie_x0
xfeed_5994 0 1 tie_x0
xfeed_5993 0 1 tie_x0
xfeed_5992 0 1 tie_x0
xfeed_5991 0 1 tie_x0
xfeed_5990 0 1 tie_x0
xfeed_199 0 1 tie_x0
xfeed_198 0 1 tie_x0
xfeed_197 0 1 tie_x0
xfeed_196 0 1 tie_x0
xfeed_195 0 1 tie_x0
xfeed_194 0 1 tie_x0
xfeed_193 0 1 tie_x0
xfeed_192 0 1 tie_x0
xfeed_191 0 1 tie_x0
xfeed_190 0 1 tie_x0
xfeed_1682 0 1 tie_x0
xfeed_1683 0 1 tie_x0
xfeed_1684 0 1 tie_x0
xfeed_1685 0 1 tie_x0
xfeed_1686 0 1 tie_x0
xfeed_1687 0 1 tie_x0
xfeed_1688 0 1 tie_x0
xfeed_1689 0 1 tie_x0
xfeed_7149 0 1 tie_x0
xfeed_7148 0 1 tie_x0
xfeed_7147 0 1 tie_x0
xfeed_7146 0 1 rowend_x0
xfeed_7145 0 1 tie_x0
xfeed_7144 0 1 tie_x0
xfeed_7143 0 1 tie_x0
xfeed_7142 0 1 tie_x0
xfeed_7141 0 1 tie_x0
xfeed_7140 0 1 tie_x0
xfeed_6619 0 1 tie_x0
xfeed_6618 0 1 tie_x0
xfeed_6617 0 1 tie_x0
xfeed_6616 0 1 tie_x0
xfeed_6615 0 1 tie_x0
xfeed_6614 0 1 tie_x0
xfeed_6613 0 1 tie_x0
xfeed_6612 0 1 tie_x0
xfeed_6611 0 1 tie_x0
xfeed_6610 0 1 tie_x0
xfeed_2309 0 1 tie_x0
xfeed_2308 0 1 tie_x0
xfeed_2307 0 1 tie_x0
xfeed_2306 0 1 tie_x0
xfeed_2305 0 1 tie_x0
xfeed_2304 0 1 tie_x0
xfeed_2303 0 1 tie_x0
xfeed_2302 0 1 tie_x0
xfeed_2301 0 1 tie_x0
xfeed_2300 0 1 tie_x0
xspare_feed_230 0 1 rowend_x0
xspare_feed_231 0 1 tie_x0
xspare_feed_232 0 1 rowend_x0
xspare_feed_233 0 1 rowend_x0
xspare_feed_234 0 1 tie_x0
xspare_feed_235 0 1 rowend_x0
xspare_feed_236 0 1 tie_x0
xspare_feed_237 0 1 rowend_x0
xspare_feed_238 0 1 rowend_x0
xsubckt_25_nao22_x1 0 1 113 122 121 125 nao22_x1
xfeed_1690 0 1 tie_x0
xfeed_1691 0 1 tie_x0
xfeed_1692 0 1 tie_x0
xfeed_1693 0 1 tie_x0
xfeed_1694 0 1 tie_x0
xfeed_1695 0 1 tie_x0
xfeed_1696 0 1 rowend_x0
xfeed_1697 0 1 tie_x0
xfeed_1698 0 1 tie_x0
xfeed_1699 0 1 tie_x0
xfeed_7159 0 1 tie_x0
xfeed_7158 0 1 tie_x0
xfeed_7157 0 1 tie_x0
xfeed_7156 0 1 tie_x0
xfeed_7155 0 1 tie_x0
xfeed_7154 0 1 tie_x0
xfeed_7153 0 1 tie_x0
xfeed_7152 0 1 tie_x0
xfeed_7151 0 1 tie_x0
xfeed_7150 0 1 tie_x0
xfeed_6629 0 1 tie_x0
xfeed_6628 0 1 tie_x0
xfeed_6627 0 1 tie_x0
xfeed_6626 0 1 tie_x0
xfeed_6625 0 1 tie_x0
xfeed_6624 0 1 tie_x0
xfeed_6623 0 1 tie_x0
xfeed_6622 0 1 tie_x0
xfeed_6621 0 1 tie_x0
xfeed_6620 0 1 tie_x0
xfeed_2319 0 1 tie_x0
xfeed_2318 0 1 tie_x0
xfeed_2317 0 1 tie_x0
xfeed_2316 0 1 tie_x0
xfeed_2315 0 1 tie_x0
xfeed_2314 0 1 tie_x0
xfeed_2313 0 1 tie_x0
xfeed_2312 0 1 tie_x0
xfeed_2311 0 1 tie_x0
xfeed_2310 0 1 tie_x0
xsubckt_67_na2_x1 0 1 204 86 205 na2_x1
xsubckt_63_na2_x1 0 1 208 83 210 na2_x1
xfeed_7169 0 1 tie_x0
xfeed_7168 0 1 tie_x0
xfeed_7167 0 1 tie_x0
xfeed_7166 0 1 tie_x0
xfeed_7165 0 1 tie_x0
xfeed_7164 0 1 tie_x0
xfeed_7163 0 1 tie_x0
xfeed_7162 0 1 tie_x0
xfeed_7161 0 1 tie_x0
xfeed_7160 0 1 tie_x0
xfeed_6639 0 1 tie_x0
xfeed_6638 0 1 tie_x0
xfeed_6637 0 1 tie_x0
xfeed_6636 0 1 tie_x0
xfeed_6635 0 1 tie_x0
xfeed_6634 0 1 tie_x0
xfeed_6633 0 1 tie_x0
xfeed_6632 0 1 tie_x0
xfeed_6631 0 1 tie_x0
xfeed_6630 0 1 tie_x0
xfeed_2329 0 1 tie_x0
xfeed_2328 0 1 tie_x0
xfeed_2327 0 1 tie_x0
xfeed_2326 0 1 tie_x0
xfeed_2325 0 1 tie_x0
xfeed_2324 0 1 tie_x0
xfeed_2323 0 1 tie_x0
xfeed_2322 0 1 tie_x0
xfeed_2321 0 1 rowend_x0
xfeed_2320 0 1 tie_x0
xsubckt_21_nxr2_x1 0 1 116 128 119 nxr2_x1
xsubckt_154_sff1_x4 0 1 4 223 56 sff1_x4
xfeed_309 0 1 tie_x0
xfeed_308 0 1 tie_x0
xfeed_307 0 1 tie_x0
xfeed_306 0 1 tie_x0
xfeed_305 0 1 tie_x0
xfeed_304 0 1 tie_x0
xfeed_303 0 1 tie_x0
xfeed_302 0 1 tie_x0
xfeed_301 0 1 tie_x0
xfeed_300 0 1 tie_x0
xfeed_7179 0 1 tie_x0
xfeed_7178 0 1 tie_x0
xfeed_7177 0 1 tie_x0
xfeed_7176 0 1 tie_x0
xfeed_7175 0 1 tie_x0
xfeed_7174 0 1 tie_x0
xfeed_7173 0 1 tie_x0
xfeed_7172 0 1 tie_x0
xfeed_7171 0 1 tie_x0
xfeed_7170 0 1 tie_x0
xfeed_6646 0 1 tie_x0
xfeed_6645 0 1 tie_x0
xfeed_6644 0 1 tie_x0
xfeed_6643 0 1 tie_x0
xfeed_6642 0 1 tie_x0
xfeed_6641 0 1 tie_x0
xfeed_6640 0 1 tie_x0
xfeed_2339 0 1 tie_x0
xfeed_2338 0 1 tie_x0
xfeed_2337 0 1 tie_x0
xfeed_2336 0 1 tie_x0
xfeed_2335 0 1 tie_x0
xfeed_2334 0 1 tie_x0
xfeed_2333 0 1 tie_x0
xfeed_2332 0 1 tie_x0
xfeed_2331 0 1 tie_x0
xfeed_2330 0 1 tie_x0
xsubckt_17_nxr2_x1 0 1 120 124 123 nxr2_x1
xfeed_1800 0 1 tie_x0
xfeed_1801 0 1 tie_x0
xfeed_1802 0 1 tie_x0
xfeed_1803 0 1 tie_x0
xfeed_1804 0 1 tie_x0
xfeed_1805 0 1 tie_x0
xfeed_1806 0 1 tie_x0
xfeed_1807 0 1 tie_x0
xfeed_6649 0 1 tie_x0
xfeed_6648 0 1 tie_x0
xfeed_6647 0 1 tie_x0
xfeed_319 0 1 tie_x0
xfeed_318 0 1 tie_x0
xfeed_317 0 1 tie_x0
xfeed_316 0 1 tie_x0
xfeed_315 0 1 tie_x0
xfeed_314 0 1 tie_x0
xfeed_313 0 1 tie_x0
xfeed_312 0 1 tie_x0
xfeed_311 0 1 tie_x0
xfeed_310 0 1 tie_x0
xfeed_1808 0 1 tie_x0
xfeed_1809 0 1 tie_x0
xfeed_7189 0 1 tie_x0
xfeed_7188 0 1 tie_x0
xfeed_7187 0 1 rowend_x0
xfeed_7186 0 1 tie_x0
xfeed_7185 0 1 tie_x0
xfeed_7184 0 1 tie_x0
xfeed_7183 0 1 tie_x0
xfeed_7182 0 1 tie_x0
xfeed_7181 0 1 tie_x0
xfeed_7180 0 1 tie_x0
xfeed_6653 0 1 tie_x0
xfeed_6652 0 1 tie_x0
xfeed_6651 0 1 tie_x0
xfeed_6650 0 1 tie_x0
xfeed_2349 0 1 tie_x0
xfeed_2348 0 1 rowend_x0
xfeed_2347 0 1 tie_x0
xfeed_2346 0 1 tie_x0
xfeed_2345 0 1 tie_x0
xfeed_2344 0 1 tie_x0
xfeed_2343 0 1 tie_x0
xfeed_2342 0 1 tie_x0
xfeed_2341 0 1 tie_x0
xfeed_2340 0 1 tie_x0
xfeed_1810 0 1 tie_x0
xfeed_1811 0 1 tie_x0
xfeed_1812 0 1 tie_x0
xfeed_1813 0 1 tie_x0
xfeed_1814 0 1 tie_x0
xfeed_6659 0 1 tie_x0
xfeed_6658 0 1 tie_x0
xfeed_6657 0 1 tie_x0
xfeed_6656 0 1 tie_x0
xfeed_6655 0 1 tie_x0
xfeed_6654 0 1 tie_x0
xfeed_329 0 1 tie_x0
xfeed_328 0 1 tie_x0
xfeed_327 0 1 tie_x0
xfeed_326 0 1 tie_x0
xfeed_325 0 1 tie_x0
xfeed_324 0 1 tie_x0
xfeed_323 0 1 tie_x0
xfeed_322 0 1 tie_x0
xfeed_321 0 1 tie_x0
xfeed_320 0 1 tie_x0
xfeed_1815 0 1 tie_x0
xfeed_1816 0 1 tie_x0
xfeed_1817 0 1 tie_x0
xfeed_1818 0 1 tie_x0
xfeed_1819 0 1 tie_x0
xfeed_7199 0 1 tie_x0
xfeed_7198 0 1 tie_x0
xfeed_7197 0 1 tie_x0
xfeed_7196 0 1 tie_x0
xfeed_7195 0 1 tie_x0
xfeed_7194 0 1 tie_x0
xfeed_7193 0 1 tie_x0
xfeed_7192 0 1 tie_x0
xfeed_7191 0 1 tie_x0
xfeed_7190 0 1 tie_x0
xfeed_6660 0 1 tie_x0
xfeed_2359 0 1 tie_x0
xfeed_2358 0 1 tie_x0
xfeed_2357 0 1 tie_x0
xfeed_2356 0 1 tie_x0
xfeed_2355 0 1 tie_x0
xfeed_2354 0 1 tie_x0
xfeed_2353 0 1 tie_x0
xfeed_2352 0 1 tie_x0
xfeed_2351 0 1 tie_x0
xfeed_2350 0 1 tie_x0
xfeed_1820 0 1 tie_x0
xfeed_1821 0 1 tie_x0
xfeed_6669 0 1 tie_x0
xfeed_6668 0 1 tie_x0
xfeed_6667 0 1 tie_x0
xfeed_6666 0 1 tie_x0
xfeed_6665 0 1 rowend_x0
xfeed_6664 0 1 tie_x0
xfeed_6663 0 1 tie_x0
xfeed_6662 0 1 tie_x0
xfeed_6661 0 1 tie_x0
xfeed_339 0 1 tie_x0
xfeed_338 0 1 tie_x0
xfeed_337 0 1 tie_x0
xfeed_336 0 1 tie_x0
xfeed_335 0 1 tie_x0
xfeed_334 0 1 tie_x0
xfeed_333 0 1 tie_x0
xfeed_332 0 1 rowend_x0
xfeed_331 0 1 tie_x0
xfeed_330 0 1 tie_x0
xfeed_1822 0 1 tie_x0
xfeed_1823 0 1 tie_x0
xfeed_1824 0 1 tie_x0
xfeed_1825 0 1 tie_x0
xfeed_1826 0 1 tie_x0
xfeed_1827 0 1 tie_x0
xfeed_1828 0 1 tie_x0
xfeed_1829 0 1 tie_x0
xfeed_2367 0 1 tie_x0
xfeed_2366 0 1 tie_x0
xfeed_2365 0 1 tie_x0
xfeed_2364 0 1 tie_x0
xfeed_2363 0 1 tie_x0
xfeed_2362 0 1 tie_x0
xfeed_2361 0 1 tie_x0
xfeed_2360 0 1 tie_x0
xfeed_6679 0 1 tie_x0
xfeed_6678 0 1 tie_x0
xfeed_6677 0 1 tie_x0
xfeed_6676 0 1 tie_x0
xfeed_6675 0 1 tie_x0
xfeed_6674 0 1 tie_x0
xfeed_6673 0 1 tie_x0
xfeed_6672 0 1 tie_x0
xfeed_6671 0 1 tie_x0
xfeed_6670 0 1 tie_x0
xfeed_2369 0 1 tie_x0
xfeed_2368 0 1 tie_x0
xfeed_349 0 1 tie_x0
xfeed_348 0 1 tie_x0
xfeed_347 0 1 tie_x0
xfeed_346 0 1 tie_x0
xfeed_345 0 1 tie_x0
xfeed_344 0 1 tie_x0
xfeed_343 0 1 tie_x0
xfeed_342 0 1 tie_x0
xfeed_341 0 1 tie_x0
xfeed_340 0 1 tie_x0
xsubckt_48_na3_x1 0 1 90 118 95 93 na3_x1
xfeed_1830 0 1 tie_x0
xfeed_1831 0 1 tie_x0
xfeed_1832 0 1 tie_x0
xfeed_1833 0 1 tie_x0
xfeed_1834 0 1 tie_x0
xfeed_1835 0 1 tie_x0
xfeed_1836 0 1 tie_x0
xfeed_1837 0 1 tie_x0
xfeed_1838 0 1 tie_x0
xfeed_1839 0 1 tie_x0
xfeed_2374 0 1 tie_x0
xfeed_2373 0 1 tie_x0
xfeed_2372 0 1 tie_x0
xfeed_2371 0 1 tie_x0
xfeed_2370 0 1 tie_x0
xfeed_6689 0 1 tie_x0
xfeed_6688 0 1 tie_x0
xfeed_6687 0 1 tie_x0
xfeed_6686 0 1 tie_x0
xfeed_6685 0 1 rowend_x0
xfeed_6684 0 1 tie_x0
xfeed_6683 0 1 tie_x0
xfeed_6682 0 1 tie_x0
xfeed_6681 0 1 tie_x0
xfeed_6680 0 1 tie_x0
xfeed_2379 0 1 tie_x0
xfeed_2378 0 1 tie_x0
xfeed_2377 0 1 tie_x0
xfeed_2376 0 1 tie_x0
xfeed_2375 0 1 tie_x0
xfeed_359 0 1 tie_x0
xfeed_358 0 1 tie_x0
xfeed_357 0 1 rowend_x0
xfeed_356 0 1 tie_x0
xfeed_355 0 1 tie_x0
xfeed_354 0 1 tie_x0
xfeed_353 0 1 tie_x0
xfeed_352 0 1 tie_x0
xfeed_351 0 1 tie_x0
xfeed_350 0 1 tie_x0
xfeed_1840 0 1 tie_x0
xfeed_1841 0 1 tie_x0
xfeed_1842 0 1 tie_x0
xfeed_1843 0 1 tie_x0
xfeed_1844 0 1 tie_x0
xfeed_1845 0 1 tie_x0
xfeed_1846 0 1 tie_x0
xfeed_1847 0 1 tie_x0
xfeed_1848 0 1 tie_x0
xfeed_1849 0 1 tie_x0
xfeed_7309 0 1 tie_x0
xfeed_7308 0 1 tie_x0
xfeed_7307 0 1 tie_x0
xfeed_7306 0 1 tie_x0
xfeed_7305 0 1 tie_x0
xfeed_7304 0 1 tie_x0
xfeed_7303 0 1 tie_x0
xfeed_7302 0 1 tie_x0
xfeed_7301 0 1 tie_x0
xfeed_7300 0 1 tie_x0
xfeed_2381 0 1 tie_x0
xfeed_2380 0 1 tie_x0
xfeed_6699 0 1 tie_x0
xfeed_6698 0 1 tie_x0
xfeed_6697 0 1 tie_x0
xfeed_6696 0 1 tie_x0
xfeed_6695 0 1 tie_x0
xfeed_6694 0 1 tie_x0
xfeed_6693 0 1 tie_x0
xfeed_6692 0 1 tie_x0
xfeed_6691 0 1 tie_x0
xfeed_6690 0 1 tie_x0
xfeed_2389 0 1 tie_x0
xfeed_2388 0 1 tie_x0
xfeed_2387 0 1 tie_x0
xfeed_2386 0 1 tie_x0
xfeed_2385 0 1 tie_x0
xfeed_2384 0 1 tie_x0
xfeed_2383 0 1 tie_x0
xfeed_2382 0 1 tie_x0
xfeed_369 0 1 tie_x0
xfeed_368 0 1 tie_x0
xfeed_367 0 1 tie_x0
xfeed_366 0 1 tie_x0
xfeed_365 0 1 tie_x0
xfeed_364 0 1 tie_x0
xfeed_363 0 1 tie_x0
xfeed_362 0 1 tie_x0
xfeed_361 0 1 tie_x0
xfeed_360 0 1 tie_x0
xfeed_1850 0 1 tie_x0
xfeed_1851 0 1 tie_x0
xfeed_1852 0 1 tie_x0
xfeed_1853 0 1 tie_x0
xfeed_1854 0 1 tie_x0
xfeed_1855 0 1 tie_x0
xfeed_1856 0 1 tie_x0
xfeed_1857 0 1 tie_x0
xfeed_1858 0 1 tie_x0
xfeed_1859 0 1 tie_x0
xfeed_7319 0 1 tie_x0
xfeed_7318 0 1 tie_x0
xfeed_7317 0 1 rowend_x0
xfeed_7316 0 1 tie_x0
xfeed_7315 0 1 tie_x0
xfeed_7314 0 1 tie_x0
xfeed_7313 0 1 tie_x0
xfeed_7312 0 1 tie_x0
xfeed_7311 0 1 tie_x0
xfeed_7310 0 1 tie_x0
xfeed_3009 0 1 tie_x0
xfeed_3008 0 1 tie_x0
xfeed_3007 0 1 tie_x0
xfeed_3006 0 1 tie_x0
xfeed_3005 0 1 tie_x0
xfeed_3004 0 1 tie_x0
xfeed_3003 0 1 tie_x0
xfeed_3002 0 1 tie_x0
xfeed_3001 0 1 tie_x0
xfeed_3000 0 1 tie_x0
xfeed_2399 0 1 tie_x0
xfeed_2398 0 1 tie_x0
xfeed_2397 0 1 tie_x0
xfeed_2396 0 1 rowend_x0
xfeed_2395 0 1 tie_x0
xfeed_2394 0 1 tie_x0
xfeed_2393 0 1 tie_x0
xfeed_2392 0 1 tie_x0
xfeed_2391 0 1 tie_x0
xfeed_2390 0 1 tie_x0
xfeed_379 0 1 tie_x0
xfeed_378 0 1 tie_x0
xfeed_377 0 1 tie_x0
xfeed_376 0 1 tie_x0
xfeed_375 0 1 tie_x0
xfeed_374 0 1 tie_x0
xfeed_373 0 1 tie_x0
xfeed_372 0 1 tie_x0
xfeed_371 0 1 tie_x0
xfeed_370 0 1 tie_x0
xfeed_1860 0 1 tie_x0
xfeed_1861 0 1 tie_x0
xfeed_1862 0 1 tie_x0
xfeed_1863 0 1 tie_x0
xfeed_1864 0 1 tie_x0
xfeed_1865 0 1 tie_x0
xfeed_1866 0 1 tie_x0
xfeed_1867 0 1 tie_x0
xfeed_1868 0 1 tie_x0
xfeed_1869 0 1 tie_x0
xfeed_7329 0 1 tie_x0
xfeed_7328 0 1 tie_x0
xfeed_7327 0 1 tie_x0
xfeed_7326 0 1 tie_x0
xfeed_7325 0 1 tie_x0
xfeed_7324 0 1 tie_x0
xfeed_7323 0 1 tie_x0
xfeed_7322 0 1 tie_x0
xfeed_7321 0 1 tie_x0
xfeed_7320 0 1 tie_x0
xfeed_3019 0 1 tie_x0
xfeed_3018 0 1 tie_x0
xfeed_3017 0 1 tie_x0
xfeed_3016 0 1 tie_x0
xfeed_3015 0 1 tie_x0
xfeed_3014 0 1 tie_x0
xfeed_3013 0 1 tie_x0
xfeed_3012 0 1 tie_x0
xfeed_3011 0 1 tie_x0
xfeed_3010 0 1 tie_x0
xfeed_389 0 1 tie_x0
xfeed_388 0 1 tie_x0
xfeed_387 0 1 tie_x0
xfeed_386 0 1 tie_x0
xfeed_385 0 1 tie_x0
xfeed_384 0 1 tie_x0
xfeed_383 0 1 tie_x0
xfeed_382 0 1 tie_x0
xfeed_381 0 1 tie_x0
xfeed_380 0 1 rowend_x0
xfeed_1870 0 1 tie_x0
xfeed_1871 0 1 tie_x0
xfeed_1872 0 1 tie_x0
xfeed_1873 0 1 tie_x0
xfeed_1874 0 1 tie_x0
xfeed_1875 0 1 tie_x0
xfeed_1876 0 1 rowend_x0
xfeed_1877 0 1 tie_x0
xfeed_1878 0 1 tie_x0
xfeed_1879 0 1 tie_x0
xfeed_7339 0 1 tie_x0
xfeed_7338 0 1 tie_x0
xfeed_7337 0 1 rowend_x0
xfeed_7336 0 1 tie_x0
xfeed_7335 0 1 tie_x0
xfeed_7334 0 1 tie_x0
xfeed_7333 0 1 tie_x0
xfeed_7332 0 1 tie_x0
xfeed_7331 0 1 tie_x0
xfeed_7330 0 1 tie_x0
xfeed_6800 0 1 tie_x0
xfeed_3029 0 1 tie_x0
xfeed_3028 0 1 tie_x0
xfeed_3027 0 1 tie_x0
xfeed_3026 0 1 tie_x0
xfeed_3025 0 1 tie_x0
xfeed_3024 0 1 tie_x0
xfeed_3023 0 1 tie_x0
xfeed_3022 0 1 tie_x0
xfeed_3021 0 1 rowend_x0
xfeed_3020 0 1 tie_x0
xsubckt_52_ao22_x2 0 1 87 101 100 97 ao22_x2
xfeed_6809 0 1 tie_x0
xfeed_6808 0 1 tie_x0
xfeed_6807 0 1 tie_x0
xfeed_6806 0 1 tie_x0
xfeed_6805 0 1 tie_x0
xfeed_6804 0 1 tie_x0
xfeed_6803 0 1 tie_x0
xfeed_6802 0 1 tie_x0
xfeed_6801 0 1 tie_x0
xfeed_399 0 1 tie_x0
xfeed_398 0 1 tie_x0
xfeed_397 0 1 tie_x0
xfeed_396 0 1 tie_x0
xfeed_395 0 1 tie_x0
xfeed_394 0 1 tie_x0
xfeed_393 0 1 tie_x0
xfeed_392 0 1 tie_x0
xfeed_391 0 1 tie_x0
xfeed_390 0 1 tie_x0
xsubckt_29_na4_x1 0 1 109 18 17 12 11 na4_x1
xfeed_1880 0 1 tie_x0
xfeed_1881 0 1 tie_x0
xfeed_1882 0 1 tie_x0
xfeed_1883 0 1 tie_x0
xfeed_1884 0 1 tie_x0
xfeed_1885 0 1 tie_x0
xfeed_1886 0 1 tie_x0
xfeed_1887 0 1 tie_x0
xfeed_1888 0 1 tie_x0
xfeed_1889 0 1 tie_x0
xfeed_7346 0 1 tie_x0
xfeed_7345 0 1 tie_x0
xfeed_7344 0 1 tie_x0
xfeed_7343 0 1 tie_x0
xfeed_7342 0 1 tie_x0
xfeed_7341 0 1 tie_x0
xfeed_7340 0 1 tie_x0
xfeed_3039 0 1 tie_x0
xfeed_3038 0 1 tie_x0
xfeed_3037 0 1 tie_x0
xfeed_3036 0 1 tie_x0
xfeed_3035 0 1 tie_x0
xfeed_3034 0 1 tie_x0
xfeed_3033 0 1 tie_x0
xfeed_3032 0 1 tie_x0
xfeed_3031 0 1 tie_x0
xfeed_3030 0 1 tie_x0
xfeed_2507 0 1 tie_x0
xfeed_2506 0 1 tie_x0
xfeed_2505 0 1 tie_x0
xfeed_2504 0 1 tie_x0
xfeed_2503 0 1 tie_x0
xfeed_2502 0 1 tie_x0
xfeed_2501 0 1 tie_x0
xfeed_2500 0 1 tie_x0
xfeed_7349 0 1 tie_x0
xfeed_7348 0 1 tie_x0
xfeed_7347 0 1 tie_x0
xfeed_6819 0 1 tie_x0
xfeed_6818 0 1 tie_x0
xfeed_6817 0 1 tie_x0
xfeed_6816 0 1 tie_x0
xfeed_6815 0 1 tie_x0
xfeed_6814 0 1 tie_x0
xfeed_6813 0 1 tie_x0
xfeed_6812 0 1 tie_x0
xfeed_6811 0 1 tie_x0
xfeed_6810 0 1 tie_x0
xfeed_2509 0 1 tie_x0
xfeed_2508 0 1 tie_x0
xfeed_1890 0 1 tie_x0
xfeed_1891 0 1 tie_x0
xfeed_1892 0 1 tie_x0
xfeed_1893 0 1 tie_x0
xfeed_1894 0 1 tie_x0
xfeed_1895 0 1 tie_x0
xfeed_1896 0 1 tie_x0
xfeed_1897 0 1 tie_x0
xfeed_1898 0 1 tie_x0
xfeed_1899 0 1 tie_x0
xfeed_7353 0 1 tie_x0
xfeed_7352 0 1 tie_x0
xfeed_7351 0 1 tie_x0
xfeed_7350 0 1 tie_x0
xfeed_3049 0 1 tie_x0
xfeed_3048 0 1 tie_x0
xfeed_3047 0 1 tie_x0
xfeed_3046 0 1 tie_x0
xfeed_3045 0 1 tie_x0
xfeed_3044 0 1 tie_x0
xfeed_3043 0 1 tie_x0
xfeed_3042 0 1 tie_x0
xfeed_3041 0 1 tie_x0
xfeed_3040 0 1 tie_x0
xfeed_2514 0 1 tie_x0
xfeed_2513 0 1 tie_x0
xfeed_2512 0 1 tie_x0
xfeed_2511 0 1 tie_x0
xfeed_2510 0 1 tie_x0
xsubckt_76_na2_x1 0 1 196 12 15 na2_x1
xsubckt_61_nxr2_x1 0 1 210 213 212 nxr2_x1
xfeed_7359 0 1 tie_x0
xfeed_7358 0 1 tie_x0
xfeed_7357 0 1 tie_x0
xfeed_7356 0 1 tie_x0
xfeed_7355 0 1 tie_x0
xfeed_7354 0 1 tie_x0
xfeed_6829 0 1 tie_x0
xfeed_6828 0 1 tie_x0
xfeed_6827 0 1 tie_x0
xfeed_6826 0 1 tie_x0
xfeed_6825 0 1 tie_x0
xfeed_6824 0 1 tie_x0
xfeed_6823 0 1 tie_x0
xfeed_6822 0 1 tie_x0
xfeed_6821 0 1 tie_x0
xfeed_6820 0 1 tie_x0
xfeed_2519 0 1 tie_x0
xfeed_2518 0 1 tie_x0
xfeed_2517 0 1 tie_x0
xfeed_2516 0 1 tie_x0
xfeed_2515 0 1 tie_x0
xfeed_7360 0 1 tie_x0
xfeed_3059 0 1 tie_x0
xfeed_3058 0 1 tie_x0
xfeed_3057 0 1 tie_x0
xfeed_3056 0 1 tie_x0
xfeed_3055 0 1 tie_x0
xfeed_3054 0 1 tie_x0
xfeed_3053 0 1 tie_x0
xfeed_3052 0 1 tie_x0
xfeed_3051 0 1 tie_x0
xfeed_3050 0 1 tie_x0
xfeed_2521 0 1 tie_x0
xfeed_2520 0 1 tie_x0
xfeed_7369 0 1 tie_x0
xfeed_7368 0 1 tie_x0
xfeed_7367 0 1 tie_x0
xfeed_7366 0 1 tie_x0
xfeed_7365 0 1 tie_x0
xfeed_7364 0 1 tie_x0
xfeed_7363 0 1 tie_x0
xfeed_7362 0 1 tie_x0
xfeed_7361 0 1 tie_x0
xfeed_6839 0 1 tie_x0
xfeed_6838 0 1 tie_x0
xfeed_6837 0 1 tie_x0
xfeed_6836 0 1 tie_x0
xfeed_6835 0 1 tie_x0
xfeed_6834 0 1 tie_x0
xfeed_6833 0 1 tie_x0
xfeed_6832 0 1 tie_x0
xfeed_6831 0 1 tie_x0
xfeed_6830 0 1 tie_x0
xfeed_2529 0 1 tie_x0
xfeed_2528 0 1 tie_x0
xfeed_2527 0 1 tie_x0
xfeed_2526 0 1 tie_x0
xfeed_2525 0 1 tie_x0
xfeed_2524 0 1 tie_x0
xfeed_2523 0 1 rowend_x0
xfeed_2522 0 1 tie_x0
xfeed_509 0 1 tie_x0
xfeed_508 0 1 tie_x0
xfeed_507 0 1 tie_x0
xfeed_506 0 1 tie_x0
xfeed_505 0 1 tie_x0
xfeed_504 0 1 tie_x0
xfeed_503 0 1 tie_x0
xfeed_502 0 1 tie_x0
xfeed_501 0 1 tie_x0
xfeed_500 0 1 tie_x0
xsubckt_130_xr2_x4 0 1 150 76 5 xr2_x4
xfeed_3067 0 1 tie_x0
xfeed_3066 0 1 tie_x0
xfeed_3065 0 1 tie_x0
xfeed_3064 0 1 tie_x0
xfeed_3063 0 1 tie_x0
xfeed_3062 0 1 tie_x0
xfeed_3061 0 1 tie_x0
xfeed_3060 0 1 tie_x0
xfeed_7379 0 1 tie_x0
xfeed_7378 0 1 tie_x0
xfeed_7377 0 1 tie_x0
xfeed_7376 0 1 tie_x0
xfeed_7375 0 1 tie_x0
xfeed_7374 0 1 tie_x0
xfeed_7373 0 1 tie_x0
xfeed_7372 0 1 tie_x0
xfeed_7371 0 1 tie_x0
xfeed_7370 0 1 tie_x0
xfeed_6849 0 1 tie_x0
xfeed_6848 0 1 tie_x0
xfeed_6847 0 1 tie_x0
xfeed_6846 0 1 tie_x0
xfeed_6845 0 1 tie_x0
xfeed_6844 0 1 tie_x0
xfeed_6843 0 1 tie_x0
xfeed_6842 0 1 tie_x0
xfeed_6841 0 1 tie_x0
xfeed_6840 0 1 tie_x0
xfeed_3069 0 1 tie_x0
xfeed_3068 0 1 tie_x0
xfeed_2539 0 1 tie_x0
xfeed_2538 0 1 tie_x0
xfeed_2537 0 1 tie_x0
xfeed_2536 0 1 tie_x0
xfeed_2535 0 1 tie_x0
xfeed_2534 0 1 tie_x0
xfeed_2533 0 1 tie_x0
xfeed_2532 0 1 tie_x0
xfeed_2531 0 1 tie_x0
xfeed_2530 0 1 tie_x0
xfeed_519 0 1 tie_x0
xfeed_518 0 1 tie_x0
xfeed_517 0 1 tie_x0
xfeed_516 0 1 tie_x0
xfeed_515 0 1 tie_x0
xfeed_514 0 1 tie_x0
xfeed_513 0 1 tie_x0
xfeed_512 0 1 tie_x0
xfeed_511 0 1 tie_x0
xfeed_510 0 1 tie_x0
xfeed_3074 0 1 tie_x0
xfeed_3073 0 1 tie_x0
xfeed_3072 0 1 tie_x0
xfeed_3071 0 1 tie_x0
xfeed_3070 0 1 tie_x0
xfeed_7389 0 1 tie_x0
xfeed_7388 0 1 tie_x0
xfeed_7387 0 1 tie_x0
xfeed_7386 0 1 rowend_x0
xfeed_7385 0 1 tie_x0
xfeed_7384 0 1 tie_x0
xfeed_7383 0 1 tie_x0
xfeed_7382 0 1 tie_x0
xfeed_7381 0 1 tie_x0
xfeed_7380 0 1 tie_x0
xfeed_6859 0 1 tie_x0
xfeed_6858 0 1 tie_x0
xfeed_6857 0 1 tie_x0
xfeed_6856 0 1 tie_x0
xfeed_6855 0 1 tie_x0
xfeed_6854 0 1 tie_x0
xfeed_6853 0 1 tie_x0
xfeed_6852 0 1 tie_x0
xfeed_6851 0 1 tie_x0
xfeed_6850 0 1 tie_x0
xfeed_3079 0 1 tie_x0
xfeed_3078 0 1 tie_x0
xfeed_3077 0 1 tie_x0
xfeed_3076 0 1 tie_x0
xfeed_3075 0 1 tie_x0
xfeed_2549 0 1 tie_x0
xfeed_2548 0 1 tie_x0
xfeed_2547 0 1 rowend_x0
xfeed_2546 0 1 tie_x0
xfeed_2545 0 1 tie_x0
xfeed_2544 0 1 tie_x0
xfeed_2543 0 1 tie_x0
xfeed_2542 0 1 tie_x0
xfeed_2541 0 1 tie_x0
xfeed_2540 0 1 tie_x0
xfeed_529 0 1 tie_x0
xfeed_528 0 1 tie_x0
xfeed_527 0 1 tie_x0
xfeed_526 0 1 tie_x0
xfeed_525 0 1 tie_x0
xfeed_524 0 1 tie_x0
xfeed_523 0 1 tie_x0
xfeed_522 0 1 tie_x0
xfeed_521 0 1 tie_x0
xfeed_520 0 1 tie_x0
xfeed_8009 0 1 tie_x0
xfeed_8008 0 1 tie_x0
xfeed_8007 0 1 tie_x0
xfeed_8006 0 1 tie_x0
xfeed_8005 0 1 tie_x0
xfeed_8004 0 1 tie_x0
xfeed_8003 0 1 tie_x0
xfeed_8002 0 1 tie_x0
xfeed_8001 0 1 tie_x0
xfeed_8000 0 1 tie_x0
xfeed_3081 0 1 tie_x0
xfeed_3080 0 1 tie_x0
xsubckt_72_nao22_x1 0 1 225 88 201 200 nao22_x1
xsubckt_1_inv_x1 0 1 134 7 inv_x1
xsubckt_3_inv_x1 0 1 132 15 inv_x1
xfeed_7399 0 1 tie_x0
xfeed_7398 0 1 tie_x0
xfeed_7397 0 1 tie_x0
xfeed_7396 0 1 tie_x0
xfeed_7395 0 1 tie_x0
xfeed_7394 0 1 tie_x0
xfeed_7393 0 1 tie_x0
xfeed_7392 0 1 tie_x0
xfeed_7391 0 1 tie_x0
xfeed_7390 0 1 tie_x0
xfeed_6869 0 1 tie_x0
xfeed_6868 0 1 tie_x0
xfeed_6867 0 1 tie_x0
xfeed_6866 0 1 tie_x0
xfeed_6865 0 1 tie_x0
xfeed_6864 0 1 tie_x0
xfeed_6863 0 1 tie_x0
xfeed_6862 0 1 tie_x0
xfeed_6861 0 1 tie_x0
xfeed_6860 0 1 tie_x0
xfeed_3089 0 1 tie_x0
xfeed_3088 0 1 tie_x0
xfeed_3087 0 1 tie_x0
xfeed_3086 0 1 tie_x0
xfeed_3085 0 1 tie_x0
xfeed_3084 0 1 tie_x0
xfeed_3083 0 1 tie_x0
xfeed_3082 0 1 tie_x0
xfeed_2559 0 1 tie_x0
xfeed_2558 0 1 tie_x0
xfeed_2557 0 1 tie_x0
xfeed_2556 0 1 tie_x0
xfeed_2555 0 1 tie_x0
xfeed_2554 0 1 tie_x0
xfeed_2553 0 1 tie_x0
xfeed_2552 0 1 tie_x0
xfeed_2551 0 1 tie_x0
xfeed_2550 0 1 tie_x0
xfeed_539 0 1 tie_x0
xfeed_538 0 1 tie_x0
xfeed_537 0 1 tie_x0
xfeed_536 0 1 tie_x0
xfeed_535 0 1 tie_x0
xfeed_534 0 1 tie_x0
xfeed_533 0 1 tie_x0
xfeed_532 0 1 tie_x0
xfeed_531 0 1 tie_x0
xfeed_530 0 1 tie_x0
xfeed_8019 0 1 tie_x0
xfeed_8018 0 1 tie_x0
xfeed_8017 0 1 tie_x0
xfeed_8016 0 1 tie_x0
xfeed_8015 0 1 tie_x0
xfeed_8014 0 1 tie_x0
xfeed_8013 0 1 tie_x0
xfeed_8012 0 1 tie_x0
xfeed_8011 0 1 tie_x0
xfeed_8010 0 1 tie_x0
xfeed_6879 0 1 tie_x0
xfeed_6878 0 1 tie_x0
xfeed_6877 0 1 tie_x0
xfeed_6876 0 1 tie_x0
xfeed_6875 0 1 tie_x0
xfeed_6874 0 1 tie_x0
xfeed_6873 0 1 tie_x0
xfeed_6872 0 1 tie_x0
xfeed_6871 0 1 tie_x0
xfeed_6870 0 1 tie_x0
xfeed_3099 0 1 tie_x0
xfeed_3098 0 1 tie_x0
xfeed_3097 0 1 tie_x0
xfeed_3096 0 1 tie_x0
xfeed_3095 0 1 tie_x0
xfeed_3094 0 1 tie_x0
xfeed_3093 0 1 tie_x0
xfeed_3092 0 1 tie_x0
xfeed_3091 0 1 tie_x0
xfeed_3090 0 1 tie_x0
xfeed_2569 0 1 tie_x0
xfeed_2568 0 1 tie_x0
xfeed_2567 0 1 tie_x0
xfeed_2566 0 1 tie_x0
xfeed_2565 0 1 tie_x0
xfeed_2564 0 1 tie_x0
xfeed_2563 0 1 tie_x0
xfeed_2562 0 1 tie_x0
xfeed_2561 0 1 tie_x0
xfeed_2560 0 1 tie_x0
xfeed_549 0 1 tie_x0
xfeed_548 0 1 tie_x0
xfeed_547 0 1 tie_x0
xfeed_546 0 1 tie_x0
xfeed_545 0 1 tie_x0
xfeed_544 0 1 tie_x0
xfeed_543 0 1 tie_x0
xfeed_542 0 1 tie_x0
xfeed_541 0 1 tie_x0
xfeed_540 0 1 tie_x0
xsubckt_14_a2_x2 0 1 123 18 12 a2_x2
xfeed_8029 0 1 tie_x0
xfeed_8028 0 1 tie_x0
xfeed_8027 0 1 tie_x0
xfeed_8026 0 1 tie_x0
xfeed_8025 0 1 tie_x0
xfeed_8024 0 1 tie_x0
xfeed_8023 0 1 tie_x0
xfeed_8022 0 1 tie_x0
xfeed_8021 0 1 tie_x0
xfeed_8020 0 1 tie_x0
xsubckt_131_nxr2_x1 0 1 149 154 150 nxr2_x1
xfeed_6889 0 1 tie_x0
xfeed_6888 0 1 tie_x0
xfeed_6887 0 1 tie_x0
xfeed_6886 0 1 tie_x0
xfeed_6885 0 1 tie_x0
xfeed_6884 0 1 tie_x0
xfeed_6883 0 1 tie_x0
xfeed_6882 0 1 tie_x0
xfeed_6881 0 1 tie_x0
xfeed_6880 0 1 tie_x0
xfeed_2579 0 1 tie_x0
xfeed_2578 0 1 tie_x0
xfeed_2577 0 1 tie_x0
xfeed_2576 0 1 tie_x0
xfeed_2575 0 1 tie_x0
xfeed_2574 0 1 tie_x0
xfeed_2573 0 1 tie_x0
xfeed_2572 0 1 tie_x0
xfeed_2571 0 1 tie_x0
xfeed_2570 0 1 tie_x0
xfeed_559 0 1 tie_x0
xfeed_558 0 1 tie_x0
xfeed_557 0 1 tie_x0
xfeed_556 0 1 tie_x0
xfeed_555 0 1 tie_x0
xfeed_554 0 1 tie_x0
xfeed_553 0 1 tie_x0
xfeed_552 0 1 tie_x0
xfeed_551 0 1 tie_x0
xfeed_550 0 1 tie_x0
xfeed_8039 0 1 tie_x0
xfeed_8038 0 1 tie_x0
xfeed_8037 0 1 tie_x0
xfeed_8036 0 1 tie_x0
xfeed_8035 0 1 tie_x0
xfeed_8034 0 1 tie_x0
xfeed_8033 0 1 tie_x0
xfeed_8032 0 1 tie_x0
xfeed_8031 0 1 tie_x0
xfeed_8030 0 1 tie_x0
xfeed_7500 0 1 tie_x0
xfeed_7509 0 1 tie_x0
xfeed_7508 0 1 tie_x0
xfeed_7507 0 1 tie_x0
xfeed_7506 0 1 tie_x0
xfeed_7505 0 1 tie_x0
xfeed_7504 0 1 tie_x0
xfeed_7503 0 1 tie_x0
xfeed_7502 0 1 tie_x0
xfeed_7501 0 1 tie_x0
xfeed_6899 0 1 tie_x0
xfeed_6898 0 1 tie_x0
xfeed_6897 0 1 tie_x0
xfeed_6896 0 1 tie_x0
xfeed_6895 0 1 tie_x0
xfeed_6894 0 1 tie_x0
xfeed_6893 0 1 tie_x0
xfeed_6892 0 1 tie_x0
xfeed_6891 0 1 tie_x0
xfeed_6890 0 1 tie_x0
xfeed_2589 0 1 tie_x0
xfeed_2588 0 1 tie_x0
xfeed_2587 0 1 tie_x0
xfeed_2586 0 1 tie_x0
xfeed_2585 0 1 tie_x0
xfeed_2584 0 1 tie_x0
xfeed_2583 0 1 tie_x0
xfeed_2582 0 1 tie_x0
xfeed_2581 0 1 tie_x0
xfeed_2580 0 1 tie_x0
xfeed_569 0 1 tie_x0
xfeed_568 0 1 tie_x0
xfeed_567 0 1 rowend_x0
xfeed_566 0 1 tie_x0
xfeed_565 0 1 tie_x0
xfeed_564 0 1 tie_x0
xfeed_563 0 1 tie_x0
xfeed_562 0 1 tie_x0
xfeed_561 0 1 tie_x0
xfeed_560 0 1 tie_x0
xfeed_8046 0 1 tie_x0
xfeed_8045 0 1 tie_x0
xfeed_8044 0 1 tie_x0
xfeed_8043 0 1 tie_x0
xfeed_8042 0 1 tie_x0
xfeed_8041 0 1 tie_x0
xfeed_8040 0 1 tie_x0
xfeed_3207 0 1 tie_x0
xfeed_3206 0 1 tie_x0
xfeed_3205 0 1 tie_x0
xfeed_3204 0 1 tie_x0
xfeed_3203 0 1 tie_x0
xfeed_3202 0 1 tie_x0
xfeed_3201 0 1 tie_x0
xfeed_3200 0 1 tie_x0
xfeed_8049 0 1 tie_x0
xfeed_8048 0 1 tie_x0
xfeed_8047 0 1 tie_x0
xfeed_7519 0 1 tie_x0
xfeed_7518 0 1 tie_x0
xfeed_7517 0 1 tie_x0
xfeed_7516 0 1 tie_x0
xfeed_7515 0 1 tie_x0
xfeed_7514 0 1 tie_x0
xfeed_7513 0 1 tie_x0
xfeed_7512 0 1 tie_x0
xfeed_7511 0 1 tie_x0
xfeed_7510 0 1 tie_x0
xfeed_3209 0 1 tie_x0
xfeed_3208 0 1 tie_x0
xfeed_2599 0 1 tie_x0
xfeed_2598 0 1 tie_x0
xfeed_2597 0 1 tie_x0
xfeed_2596 0 1 tie_x0
xfeed_2595 0 1 tie_x0
xfeed_2594 0 1 tie_x0
xfeed_2593 0 1 tie_x0
xfeed_2592 0 1 tie_x0
xfeed_2591 0 1 tie_x0
xfeed_2590 0 1 tie_x0
xfeed_576 0 1 tie_x0
xfeed_575 0 1 tie_x0
xfeed_574 0 1 tie_x0
xfeed_573 0 1 tie_x0
xfeed_572 0 1 tie_x0
xfeed_571 0 1 tie_x0
xfeed_570 0 1 tie_x0
xfeed_8053 0 1 tie_x0
xfeed_8052 0 1 tie_x0
xfeed_8051 0 1 tie_x0
xfeed_8050 0 1 tie_x0
xfeed_3214 0 1 tie_x0
xfeed_3213 0 1 tie_x0
xfeed_3212 0 1 tie_x0
xfeed_3211 0 1 tie_x0
xfeed_3210 0 1 tie_x0
xfeed_579 0 1 tie_x0
xfeed_578 0 1 tie_x0
xfeed_577 0 1 tie_x0
xfeed_8059 0 1 tie_x0
xfeed_8058 0 1 tie_x0
xfeed_8057 0 1 tie_x0
xfeed_8056 0 1 tie_x0
xfeed_8055 0 1 tie_x0
xfeed_8054 0 1 tie_x0
xfeed_7529 0 1 tie_x0
xfeed_7528 0 1 tie_x0
xfeed_7527 0 1 tie_x0
xfeed_7526 0 1 tie_x0
xfeed_7525 0 1 tie_x0
xfeed_7524 0 1 tie_x0
xfeed_7523 0 1 tie_x0
xfeed_7522 0 1 tie_x0
xfeed_7521 0 1 tie_x0
xfeed_7520 0 1 tie_x0
xfeed_3219 0 1 tie_x0
xfeed_3218 0 1 tie_x0
xfeed_3217 0 1 tie_x0
xfeed_3216 0 1 tie_x0
xfeed_3215 0 1 tie_x0
xfeed_583 0 1 tie_x0
xfeed_582 0 1 tie_x0
xfeed_581 0 1 tie_x0
xfeed_580 0 1 tie_x0
xfeed_8060 0 1 tie_x0
xfeed_3221 0 1 tie_x0
xfeed_3220 0 1 tie_x0
xfeed_589 0 1 tie_x0
xfeed_588 0 1 tie_x0
xfeed_587 0 1 tie_x0
xfeed_586 0 1 tie_x0
xfeed_585 0 1 tie_x0
xfeed_584 0 1 tie_x0
xfeed_8069 0 1 tie_x0
xfeed_8068 0 1 tie_x0
xfeed_8067 0 1 tie_x0
xfeed_8066 0 1 tie_x0
xfeed_8065 0 1 tie_x0
xfeed_8064 0 1 tie_x0
xfeed_8063 0 1 tie_x0
xfeed_8062 0 1 tie_x0
xfeed_8061 0 1 tie_x0
xfeed_7539 0 1 tie_x0
xfeed_7538 0 1 tie_x0
xfeed_7537 0 1 tie_x0
xfeed_7536 0 1 tie_x0
xfeed_7535 0 1 tie_x0
xfeed_7534 0 1 tie_x0
xfeed_7533 0 1 tie_x0
xfeed_7532 0 1 tie_x0
xfeed_7531 0 1 tie_x0
xfeed_7530 0 1 tie_x0
xfeed_3229 0 1 tie_x0
xfeed_3228 0 1 tie_x0
xfeed_3227 0 1 tie_x0
xfeed_3226 0 1 tie_x0
xfeed_3225 0 1 tie_x0
xfeed_3224 0 1 tie_x0
xfeed_3223 0 1 tie_x0
xfeed_3222 0 1 tie_x0
xfeed_590 0 1 tie_x0
xfeed_599 0 1 tie_x0
xfeed_598 0 1 tie_x0
xfeed_597 0 1 tie_x0
xfeed_596 0 1 tie_x0
xfeed_595 0 1 tie_x0
xfeed_594 0 1 tie_x0
xfeed_593 0 1 tie_x0
xfeed_592 0 1 tie_x0
xfeed_591 0 1 tie_x0
xsubckt_160_sff1_x4 0 1 77 217 40 sff1_x4
xfeed_8079 0 1 tie_x0
xfeed_8078 0 1 tie_x0
xfeed_8077 0 1 tie_x0
xfeed_8076 0 1 tie_x0
xfeed_8075 0 1 tie_x0
xfeed_8074 0 1 tie_x0
xfeed_8073 0 1 tie_x0
xfeed_8072 0 1 tie_x0
xfeed_8071 0 1 tie_x0
xfeed_8070 0 1 tie_x0
xfeed_7549 0 1 tie_x0
xfeed_7548 0 1 tie_x0
xfeed_7547 0 1 tie_x0
xfeed_7546 0 1 tie_x0
xfeed_7545 0 1 tie_x0
xfeed_7544 0 1 tie_x0
xfeed_7543 0 1 tie_x0
xfeed_7542 0 1 tie_x0
xfeed_7541 0 1 tie_x0
xfeed_7540 0 1 tie_x0
xfeed_3239 0 1 tie_x0
xfeed_3238 0 1 tie_x0
xfeed_3237 0 1 tie_x0
xfeed_3236 0 1 tie_x0
xfeed_3235 0 1 tie_x0
xfeed_3234 0 1 tie_x0
xfeed_3233 0 1 tie_x0
xfeed_3232 0 1 tie_x0
xfeed_3231 0 1 tie_x0
xfeed_3230 0 1 tie_x0
xfeed_2709 0 1 tie_x0
xfeed_2708 0 1 tie_x0
xfeed_2707 0 1 tie_x0
xfeed_2706 0 1 tie_x0
xfeed_2705 0 1 tie_x0
xfeed_2704 0 1 tie_x0
xfeed_2703 0 1 tie_x0
xfeed_2702 0 1 tie_x0
xfeed_2701 0 1 tie_x0
xfeed_2700 0 1 tie_x0
xsubckt_89_na2_x1 0 1 184 186 185 na2_x1
xsubckt_156_sff1_x4 0 1 81 221 34 sff1_x4
xfeed_8089 0 1 tie_x0
xfeed_8088 0 1 tie_x0
xfeed_8087 0 1 tie_x0
xfeed_8086 0 1 tie_x0
xfeed_8085 0 1 tie_x0
xfeed_8084 0 1 tie_x0
xfeed_8083 0 1 tie_x0
xfeed_8082 0 1 tie_x0
xfeed_8081 0 1 tie_x0
xfeed_8080 0 1 tie_x0
xfeed_7559 0 1 tie_x0
xfeed_7558 0 1 tie_x0
xfeed_7557 0 1 tie_x0
xfeed_7556 0 1 tie_x0
xfeed_7555 0 1 tie_x0
xfeed_7554 0 1 tie_x0
xfeed_7553 0 1 tie_x0
xfeed_7552 0 1 tie_x0
xfeed_7551 0 1 tie_x0
xfeed_7550 0 1 tie_x0
xfeed_3249 0 1 tie_x0
xfeed_3248 0 1 tie_x0
xfeed_3247 0 1 tie_x0
xfeed_3246 0 1 tie_x0
xfeed_3245 0 1 tie_x0
xfeed_3244 0 1 tie_x0
xfeed_3243 0 1 tie_x0
xfeed_3242 0 1 tie_x0
xfeed_3241 0 1 tie_x0
xfeed_3240 0 1 tie_x0
xfeed_2719 0 1 tie_x0
xfeed_2718 0 1 tie_x0
xfeed_2717 0 1 tie_x0
xfeed_2716 0 1 tie_x0
xfeed_2715 0 1 tie_x0
xfeed_2714 0 1 tie_x0
xfeed_2713 0 1 tie_x0
xfeed_2712 0 1 tie_x0
xfeed_2711 0 1 rowend_x0
xfeed_2710 0 1 tie_x0
xsubckt_108_nxr2_x1 0 1 169 79 8 nxr2_x1
xsubckt_143_xr2_x4 0 1 139 74 3 xr2_x4
xfeed_8099 0 1 tie_x0
xfeed_8098 0 1 tie_x0
xfeed_8097 0 1 tie_x0
xfeed_8096 0 1 tie_x0
xfeed_8095 0 1 tie_x0
xfeed_8094 0 1 tie_x0
xfeed_8093 0 1 tie_x0
xfeed_8092 0 1 tie_x0
xfeed_8091 0 1 tie_x0
xfeed_8090 0 1 tie_x0
xfeed_7569 0 1 tie_x0
xfeed_7568 0 1 rowend_x0
xfeed_7567 0 1 tie_x0
xfeed_7566 0 1 tie_x0
xfeed_7565 0 1 tie_x0
xfeed_7564 0 1 tie_x0
xfeed_7563 0 1 tie_x0
xfeed_7562 0 1 tie_x0
xfeed_7561 0 1 tie_x0
xfeed_7560 0 1 tie_x0
xfeed_3259 0 1 tie_x0
xfeed_3258 0 1 tie_x0
xfeed_3257 0 1 tie_x0
xfeed_3256 0 1 tie_x0
xfeed_3255 0 1 tie_x0
xfeed_3254 0 1 tie_x0
xfeed_3253 0 1 tie_x0
xfeed_3252 0 1 tie_x0
xfeed_3251 0 1 tie_x0
xfeed_3250 0 1 tie_x0
xfeed_2729 0 1 tie_x0
xfeed_2728 0 1 tie_x0
xfeed_2727 0 1 tie_x0
xfeed_2726 0 1 tie_x0
xfeed_2725 0 1 tie_x0
xfeed_2724 0 1 tie_x0
xfeed_2723 0 1 tie_x0
xfeed_2722 0 1 tie_x0
xfeed_2721 0 1 tie_x0
xfeed_2720 0 1 tie_x0
xfeed_709 0 1 tie_x0
xfeed_708 0 1 tie_x0
xfeed_707 0 1 tie_x0
xfeed_706 0 1 tie_x0
xfeed_705 0 1 tie_x0
xfeed_704 0 1 tie_x0
xfeed_703 0 1 tie_x0
xfeed_702 0 1 tie_x0
xfeed_701 0 1 tie_x0
xfeed_700 0 1 tie_x0
xfeed_7579 0 1 tie_x0
xfeed_7578 0 1 tie_x0
xfeed_7577 0 1 tie_x0
xfeed_7576 0 1 tie_x0
xfeed_7575 0 1 tie_x0
xfeed_7574 0 1 tie_x0
xfeed_7573 0 1 tie_x0
xfeed_7572 0 1 tie_x0
xfeed_7571 0 1 tie_x0
xfeed_7570 0 1 tie_x0
xfeed_3269 0 1 tie_x0
xfeed_3268 0 1 tie_x0
xfeed_3267 0 1 tie_x0
xfeed_3266 0 1 tie_x0
xfeed_3265 0 1 tie_x0
xfeed_3264 0 1 tie_x0
xfeed_3263 0 1 tie_x0
xfeed_3262 0 1 tie_x0
xfeed_3261 0 1 tie_x0
xfeed_3260 0 1 tie_x0
xfeed_2739 0 1 tie_x0
xfeed_2738 0 1 tie_x0
xfeed_2737 0 1 rowend_x0
xfeed_2736 0 1 tie_x0
xfeed_2735 0 1 tie_x0
xfeed_2734 0 1 tie_x0
xfeed_2733 0 1 tie_x0
xfeed_2732 0 1 tie_x0
xfeed_2731 0 1 tie_x0
xfeed_2730 0 1 tie_x0
xfeed_716 0 1 tie_x0
xfeed_715 0 1 tie_x0
xfeed_714 0 1 tie_x0
xfeed_713 0 1 tie_x0
xfeed_712 0 1 tie_x0
xfeed_711 0 1 tie_x0
xfeed_710 0 1 tie_x0
xsubckt_73_ao22_x2 0 1 199 204 202 90 ao22_x2
xfeed_719 0 1 tie_x0
xfeed_718 0 1 tie_x0
xfeed_717 0 1 tie_x0
xfeed_7589 0 1 tie_x0
xfeed_7588 0 1 tie_x0
xfeed_7587 0 1 tie_x0
xfeed_7586 0 1 tie_x0
xfeed_7585 0 1 tie_x0
xfeed_7584 0 1 tie_x0
xfeed_7583 0 1 tie_x0
xfeed_7582 0 1 tie_x0
xfeed_7581 0 1 tie_x0
xfeed_7580 0 1 tie_x0
xfeed_3279 0 1 tie_x0
xfeed_3278 0 1 tie_x0
xfeed_3277 0 1 tie_x0
xfeed_3276 0 1 tie_x0
xfeed_3275 0 1 tie_x0
xfeed_3274 0 1 tie_x0
xfeed_3273 0 1 tie_x0
xfeed_3272 0 1 tie_x0
xfeed_3271 0 1 tie_x0
xfeed_3270 0 1 tie_x0
xfeed_2749 0 1 tie_x0
xfeed_2748 0 1 tie_x0
xfeed_2747 0 1 tie_x0
xfeed_2746 0 1 tie_x0
xfeed_2745 0 1 tie_x0
xfeed_2744 0 1 tie_x0
xfeed_2743 0 1 tie_x0
xfeed_2742 0 1 tie_x0
xfeed_2741 0 1 tie_x0
xfeed_2740 0 1 tie_x0
xfeed_723 0 1 tie_x0
xfeed_722 0 1 tie_x0
xfeed_721 0 1 tie_x0
xfeed_720 0 1 tie_x0
xfeed_8200 0 1 tie_x0
xfeed_729 0 1 tie_x0
xfeed_728 0 1 tie_x0
xfeed_727 0 1 tie_x0
xfeed_726 0 1 tie_x0
xfeed_725 0 1 tie_x0
xfeed_724 0 1 rowend_x0
xfeed_8209 0 1 tie_x0
xfeed_8208 0 1 tie_x0
xfeed_8207 0 1 tie_x0
xfeed_8206 0 1 tie_x0
xfeed_8205 0 1 tie_x0
xfeed_8204 0 1 tie_x0
xfeed_8203 0 1 tie_x0
xfeed_8202 0 1 tie_x0
xfeed_8201 0 1 tie_x0
xfeed_7599 0 1 tie_x0
xfeed_7598 0 1 tie_x0
xfeed_7597 0 1 tie_x0
xfeed_7596 0 1 tie_x0
xfeed_7595 0 1 tie_x0
xfeed_7594 0 1 tie_x0
xfeed_7593 0 1 tie_x0
xfeed_7592 0 1 tie_x0
xfeed_7591 0 1 tie_x0
xfeed_7590 0 1 tie_x0
xfeed_3289 0 1 tie_x0
xfeed_3288 0 1 rowend_x0
xfeed_3287 0 1 tie_x0
xfeed_3286 0 1 tie_x0
xfeed_3285 0 1 tie_x0
xfeed_3284 0 1 tie_x0
xfeed_3283 0 1 tie_x0
xfeed_3282 0 1 tie_x0
xfeed_3281 0 1 tie_x0
xfeed_3280 0 1 tie_x0
xfeed_2759 0 1 tie_x0
xfeed_2758 0 1 tie_x0
xfeed_2757 0 1 tie_x0
xfeed_2756 0 1 tie_x0
xfeed_2755 0 1 tie_x0
xfeed_2754 0 1 tie_x0
xfeed_2753 0 1 tie_x0
xfeed_2752 0 1 tie_x0
xfeed_2751 0 1 tie_x0
xfeed_2750 0 1 tie_x0
xfeed_730 0 1 tie_x0
xsubckt_36_a3_x2 0 1 102 113 105 103 a3_x2
xfeed_739 0 1 tie_x0
xfeed_738 0 1 tie_x0
xfeed_737 0 1 tie_x0
xfeed_736 0 1 tie_x0
xfeed_735 0 1 tie_x0
xfeed_734 0 1 tie_x0
xfeed_733 0 1 tie_x0
xfeed_732 0 1 tie_x0
xfeed_731 0 1 tie_x0
xsubckt_82_nxr2_x1 0 1 190 197 193 nxr2_x1
xfeed_8219 0 1 tie_x0
xfeed_8218 0 1 tie_x0
xfeed_8217 0 1 tie_x0
xfeed_8216 0 1 tie_x0
xfeed_8215 0 1 tie_x0
xfeed_8214 0 1 tie_x0
xfeed_8213 0 1 tie_x0
xfeed_8212 0 1 tie_x0
xfeed_8211 0 1 tie_x0
xfeed_8210 0 1 tie_x0
xfeed_3299 0 1 tie_x0
xfeed_3298 0 1 tie_x0
xfeed_3297 0 1 tie_x0
xfeed_3296 0 1 tie_x0
xfeed_3295 0 1 tie_x0
xfeed_3294 0 1 tie_x0
xfeed_3293 0 1 tie_x0
xfeed_3292 0 1 tie_x0
xfeed_3291 0 1 tie_x0
xfeed_3290 0 1 tie_x0
xfeed_2769 0 1 tie_x0
xfeed_2768 0 1 tie_x0
xfeed_2767 0 1 tie_x0
xfeed_2766 0 1 tie_x0
xfeed_2765 0 1 tie_x0
xfeed_2764 0 1 tie_x0
xfeed_2763 0 1 tie_x0
xfeed_2762 0 1 tie_x0
xfeed_2761 0 1 tie_x0
xfeed_2760 0 1 tie_x0
xfeed_749 0 1 tie_x0
xfeed_748 0 1 tie_x0
xfeed_747 0 1 tie_x0
xfeed_746 0 1 tie_x0
xfeed_745 0 1 tie_x0
xfeed_744 0 1 tie_x0
xfeed_743 0 1 tie_x0
xfeed_742 0 1 tie_x0
xfeed_741 0 1 tie_x0
xfeed_740 0 1 tie_x0
xfeed_8229 0 1 tie_x0
xfeed_8228 0 1 tie_x0
xfeed_8227 0 1 tie_x0
xfeed_8226 0 1 tie_x0
xfeed_8225 0 1 tie_x0
xfeed_8224 0 1 tie_x0
xfeed_8223 0 1 tie_x0
xfeed_8222 0 1 tie_x0
xfeed_8221 0 1 tie_x0
xfeed_8220 0 1 tie_x0
xfeed_2779 0 1 tie_x0
xfeed_2778 0 1 tie_x0
xfeed_2777 0 1 tie_x0
xfeed_2776 0 1 tie_x0
xfeed_2775 0 1 tie_x0
xfeed_2774 0 1 tie_x0
xfeed_2773 0 1 tie_x0
xfeed_2772 0 1 tie_x0
xfeed_2771 0 1 tie_x0
xfeed_2770 0 1 tie_x0
xfeed_759 0 1 tie_x0
xfeed_758 0 1 tie_x0
xfeed_757 0 1 tie_x0
xfeed_756 0 1 tie_x0
xfeed_755 0 1 tie_x0
xfeed_754 0 1 tie_x0
xfeed_753 0 1 tie_x0
xfeed_752 0 1 tie_x0
xfeed_751 0 1 tie_x0
xfeed_750 0 1 tie_x0
xfeed_8239 0 1 tie_x0
xfeed_8238 0 1 tie_x0
xfeed_8237 0 1 tie_x0
xfeed_8236 0 1 tie_x0
xfeed_8235 0 1 tie_x0
xfeed_8234 0 1 tie_x0
xfeed_8233 0 1 tie_x0
xfeed_8232 0 1 tie_x0
xfeed_8231 0 1 tie_x0
xfeed_8230 0 1 tie_x0
xfeed_7709 0 1 tie_x0
xfeed_7708 0 1 tie_x0
xfeed_7707 0 1 tie_x0
xfeed_7706 0 1 tie_x0
xfeed_7705 0 1 tie_x0
xfeed_7704 0 1 tie_x0
xfeed_7703 0 1 tie_x0
xfeed_7702 0 1 tie_x0
xfeed_7701 0 1 tie_x0
xfeed_7700 0 1 tie_x0
xfeed_2789 0 1 tie_x0
xfeed_2788 0 1 tie_x0
xfeed_2787 0 1 tie_x0
xfeed_2786 0 1 tie_x0
xfeed_2785 0 1 tie_x0
xfeed_2784 0 1 tie_x0
xfeed_2783 0 1 tie_x0
xfeed_2782 0 1 tie_x0
xfeed_2781 0 1 tie_x0
xfeed_2780 0 1 tie_x0
xfeed_769 0 1 tie_x0
xfeed_768 0 1 tie_x0
xfeed_767 0 1 tie_x0
xfeed_766 0 1 tie_x0
xfeed_765 0 1 tie_x0
xfeed_764 0 1 tie_x0
xfeed_763 0 1 tie_x0
xfeed_762 0 1 tie_x0
xfeed_761 0 1 tie_x0
xfeed_760 0 1 tie_x0
xfeed_8249 0 1 tie_x0
xfeed_8248 0 1 tie_x0
xfeed_8247 0 1 tie_x0
xfeed_8246 0 1 tie_x0
xfeed_8245 0 1 tie_x0
xfeed_8244 0 1 tie_x0
xfeed_8243 0 1 tie_x0
xfeed_8242 0 1 tie_x0
xfeed_8241 0 1 tie_x0
xfeed_8240 0 1 tie_x0
xfeed_7719 0 1 tie_x0
xfeed_7718 0 1 tie_x0
xfeed_7717 0 1 tie_x0
xfeed_7716 0 1 tie_x0
xfeed_7715 0 1 tie_x0
xfeed_7714 0 1 tie_x0
xfeed_7713 0 1 tie_x0
xfeed_7712 0 1 tie_x0
xfeed_7711 0 1 tie_x0
xfeed_7710 0 1 tie_x0
xfeed_3409 0 1 tie_x0
xfeed_3408 0 1 tie_x0
xfeed_3407 0 1 tie_x0
xfeed_3406 0 1 tie_x0
xfeed_3405 0 1 tie_x0
xfeed_3404 0 1 tie_x0
xfeed_3403 0 1 tie_x0
xfeed_3402 0 1 tie_x0
xfeed_3401 0 1 tie_x0
xfeed_3400 0 1 tie_x0
xfeed_2799 0 1 tie_x0
xfeed_2798 0 1 tie_x0
xfeed_2797 0 1 tie_x0
xfeed_2796 0 1 tie_x0
xfeed_2795 0 1 tie_x0
xfeed_2794 0 1 tie_x0
xfeed_2793 0 1 tie_x0
xfeed_2792 0 1 tie_x0
xfeed_2791 0 1 tie_x0
xfeed_2790 0 1 tie_x0
xfeed_779 0 1 tie_x0
xfeed_778 0 1 tie_x0
xfeed_777 0 1 tie_x0
xfeed_776 0 1 tie_x0
xfeed_775 0 1 tie_x0
xfeed_774 0 1 tie_x0
xfeed_773 0 1 tie_x0
xfeed_772 0 1 tie_x0
xfeed_771 0 1 tie_x0
xfeed_770 0 1 tie_x0
xfeed_8259 0 1 tie_x0
xfeed_8258 0 1 tie_x0
xfeed_8257 0 1 tie_x0
xfeed_8256 0 1 tie_x0
xfeed_8255 0 1 tie_x0
xfeed_8254 0 1 tie_x0
xfeed_8253 0 1 tie_x0
xfeed_8252 0 1 tie_x0
xfeed_8251 0 1 tie_x0
xfeed_8250 0 1 tie_x0
xfeed_7729 0 1 tie_x0
xfeed_7728 0 1 tie_x0
xfeed_7727 0 1 tie_x0
xfeed_7726 0 1 tie_x0
xfeed_7725 0 1 tie_x0
xfeed_7724 0 1 tie_x0
xfeed_7723 0 1 tie_x0
xfeed_7722 0 1 tie_x0
xfeed_7721 0 1 tie_x0
xfeed_7720 0 1 tie_x0
xfeed_3419 0 1 tie_x0
xfeed_3418 0 1 tie_x0
xfeed_3417 0 1 tie_x0
xfeed_3416 0 1 tie_x0
xfeed_3415 0 1 tie_x0
xfeed_3414 0 1 tie_x0
xfeed_3413 0 1 tie_x0
xfeed_3412 0 1 tie_x0
xfeed_3411 0 1 tie_x0
xfeed_3410 0 1 tie_x0
xsubckt_139_ao22_x2 0 1 142 144 148 153 ao22_x2
xfeed_789 0 1 tie_x0
xfeed_788 0 1 tie_x0
xfeed_787 0 1 tie_x0
xfeed_786 0 1 tie_x0
xfeed_785 0 1 tie_x0
xfeed_784 0 1 tie_x0
xfeed_783 0 1 tie_x0
xfeed_782 0 1 tie_x0
xfeed_781 0 1 tie_x0
xfeed_780 0 1 tie_x0
xsubckt_92_na2_x1 0 1 181 4 2 na2_x1
xfeed_8269 0 1 tie_x0
xfeed_8268 0 1 tie_x0
xfeed_8267 0 1 tie_x0
xfeed_8266 0 1 tie_x0
xfeed_8265 0 1 tie_x0
xfeed_8264 0 1 tie_x0
xfeed_8263 0 1 tie_x0
xfeed_8262 0 1 tie_x0
xfeed_8261 0 1 tie_x0
xfeed_8260 0 1 tie_x0
xfeed_7739 0 1 tie_x0
xfeed_7738 0 1 tie_x0
xfeed_7737 0 1 tie_x0
xfeed_7736 0 1 tie_x0
xfeed_7735 0 1 tie_x0
xfeed_7734 0 1 tie_x0
xfeed_7733 0 1 tie_x0
xfeed_7732 0 1 tie_x0
xfeed_7731 0 1 tie_x0
xfeed_7730 0 1 tie_x0
xfeed_3429 0 1 tie_x0
xfeed_3428 0 1 tie_x0
xfeed_3427 0 1 tie_x0
xfeed_3426 0 1 tie_x0
xfeed_3425 0 1 tie_x0
xfeed_3424 0 1 tie_x0
xfeed_3423 0 1 tie_x0
xfeed_3422 0 1 tie_x0
xfeed_3421 0 1 tie_x0
xfeed_3420 0 1 tie_x0
xsubckt_96_na2_x1 0 1 179 81 10 na2_x1
xfeed_799 0 1 tie_x0
xfeed_798 0 1 tie_x0
xfeed_797 0 1 tie_x0
xfeed_796 0 1 tie_x0
xfeed_795 0 1 tie_x0
xfeed_794 0 1 tie_x0
xfeed_793 0 1 tie_x0
xfeed_792 0 1 tie_x0
xfeed_791 0 1 tie_x0
xfeed_790 0 1 tie_x0
xfeed_8279 0 1 tie_x0
xfeed_8278 0 1 tie_x0
xfeed_8277 0 1 tie_x0
xfeed_8276 0 1 tie_x0
xfeed_8275 0 1 tie_x0
xfeed_8274 0 1 tie_x0
xfeed_8273 0 1 tie_x0
xfeed_8272 0 1 tie_x0
xfeed_8271 0 1 tie_x0
xfeed_8270 0 1 tie_x0
xfeed_7749 0 1 tie_x0
xfeed_7748 0 1 rowend_x0
xfeed_7747 0 1 tie_x0
xfeed_7746 0 1 tie_x0
xfeed_7745 0 1 tie_x0
xfeed_7744 0 1 tie_x0
xfeed_7743 0 1 tie_x0
xfeed_7742 0 1 tie_x0
xfeed_7741 0 1 tie_x0
xfeed_7740 0 1 tie_x0
xfeed_3439 0 1 tie_x0
xfeed_3438 0 1 tie_x0
xfeed_3437 0 1 tie_x0
xfeed_3436 0 1 tie_x0
xfeed_3435 0 1 tie_x0
xfeed_3434 0 1 tie_x0
xfeed_3433 0 1 tie_x0
xfeed_3432 0 1 tie_x0
xfeed_3431 0 1 tie_x0
xfeed_3430 0 1 tie_x0
xfeed_2909 0 1 tie_x0
xfeed_2908 0 1 tie_x0
xfeed_2907 0 1 tie_x0
xfeed_2906 0 1 tie_x0
xfeed_2905 0 1 tie_x0
xfeed_2904 0 1 tie_x0
xfeed_2903 0 1 tie_x0
xfeed_2902 0 1 tie_x0
xfeed_2901 0 1 tie_x0
xfeed_2900 0 1 tie_x0
xsubckt_50_o2_x2 0 1 226 115 89 o2_x2
xsubckt_91_nao22_x1 0 1 182 131 188 184 nao22_x1
xfeed_8289 0 1 tie_x0
xfeed_8288 0 1 tie_x0
xfeed_8287 0 1 tie_x0
xfeed_8286 0 1 tie_x0
xfeed_8285 0 1 tie_x0
xfeed_8284 0 1 tie_x0
xfeed_8283 0 1 tie_x0
xfeed_8282 0 1 tie_x0
xfeed_8281 0 1 tie_x0
xfeed_8280 0 1 tie_x0
xfeed_7759 0 1 tie_x0
xfeed_7758 0 1 tie_x0
xfeed_7757 0 1 tie_x0
xfeed_7756 0 1 tie_x0
xfeed_7755 0 1 tie_x0
xfeed_7754 0 1 tie_x0
xfeed_7753 0 1 tie_x0
xfeed_7752 0 1 tie_x0
xfeed_7751 0 1 tie_x0
xfeed_7750 0 1 tie_x0
xfeed_3449 0 1 tie_x0
xfeed_3448 0 1 tie_x0
xfeed_3447 0 1 tie_x0
xfeed_3446 0 1 tie_x0
xfeed_3445 0 1 tie_x0
xfeed_3444 0 1 tie_x0
xfeed_3443 0 1 tie_x0
xfeed_3442 0 1 tie_x0
xfeed_3441 0 1 tie_x0
xfeed_3440 0 1 tie_x0
xfeed_2919 0 1 tie_x0
xfeed_2918 0 1 tie_x0
xfeed_2917 0 1 tie_x0
xfeed_2916 0 1 tie_x0
xfeed_2915 0 1 tie_x0
xfeed_2914 0 1 tie_x0
xfeed_2913 0 1 tie_x0
xfeed_2912 0 1 tie_x0
xfeed_2911 0 1 tie_x0
xfeed_2910 0 1 tie_x0
xfeed_8299 0 1 tie_x0
xfeed_8298 0 1 tie_x0
xfeed_8297 0 1 tie_x0
xfeed_8296 0 1 tie_x0
xfeed_8295 0 1 tie_x0
xfeed_8294 0 1 tie_x0
xfeed_8293 0 1 tie_x0
xfeed_8292 0 1 tie_x0
xfeed_8291 0 1 tie_x0
xfeed_8290 0 1 tie_x0
xfeed_7769 0 1 tie_x0
xfeed_7768 0 1 tie_x0
xfeed_7767 0 1 tie_x0
xfeed_7766 0 1 tie_x0
xfeed_7765 0 1 tie_x0
xfeed_7764 0 1 tie_x0
xfeed_7763 0 1 tie_x0
xfeed_7762 0 1 tie_x0
xfeed_7761 0 1 tie_x0
xfeed_7760 0 1 tie_x0
xfeed_3459 0 1 tie_x0
xfeed_3458 0 1 tie_x0
xfeed_3457 0 1 tie_x0
xfeed_3456 0 1 tie_x0
xfeed_3455 0 1 tie_x0
xfeed_3454 0 1 tie_x0
xfeed_3453 0 1 tie_x0
xfeed_3452 0 1 tie_x0
xfeed_3451 0 1 tie_x0
xfeed_3450 0 1 tie_x0
xfeed_2929 0 1 tie_x0
xfeed_2928 0 1 tie_x0
xfeed_2927 0 1 tie_x0
xfeed_2926 0 1 tie_x0
xfeed_2925 0 1 tie_x0
xfeed_2924 0 1 tie_x0
xfeed_2923 0 1 tie_x0
xfeed_2922 0 1 tie_x0
xfeed_2921 0 1 tie_x0
xfeed_2920 0 1 tie_x0
xfeed_900 0 1 tie_x0
xfeed_901 0 1 tie_x0
xfeed_902 0 1 tie_x0
xfeed_903 0 1 tie_x0
xfeed_904 0 1 tie_x0
xfeed_905 0 1 tie_x0
xfeed_906 0 1 tie_x0
xfeed_907 0 1 tie_x0
xfeed_908 0 1 tie_x0
xfeed_909 0 1 tie_x0
xfeed_7779 0 1 tie_x0
xfeed_7778 0 1 tie_x0
xfeed_7777 0 1 tie_x0
xfeed_7776 0 1 tie_x0
xfeed_7775 0 1 tie_x0
xfeed_7774 0 1 tie_x0
xfeed_7773 0 1 tie_x0
xfeed_7772 0 1 tie_x0
xfeed_7771 0 1 tie_x0
xfeed_7770 0 1 tie_x0
xfeed_3469 0 1 tie_x0
xfeed_3468 0 1 tie_x0
xfeed_3467 0 1 tie_x0
xfeed_3466 0 1 tie_x0
xfeed_3465 0 1 tie_x0
xfeed_3464 0 1 tie_x0
xfeed_3463 0 1 tie_x0
xfeed_3462 0 1 tie_x0
xfeed_3461 0 1 tie_x0
xfeed_3460 0 1 tie_x0
xfeed_2939 0 1 tie_x0
xfeed_2938 0 1 tie_x0
xfeed_2937 0 1 tie_x0
xfeed_2936 0 1 tie_x0
xfeed_2935 0 1 tie_x0
xfeed_2934 0 1 tie_x0
xfeed_2933 0 1 tie_x0
xfeed_2932 0 1 tie_x0
xfeed_2931 0 1 tie_x0
xfeed_2930 0 1 tie_x0
xfeed_910 0 1 tie_x0
xfeed_911 0 1 tie_x0
xfeed_912 0 1 tie_x0
xfeed_913 0 1 tie_x0
xfeed_914 0 1 tie_x0
xfeed_915 0 1 tie_x0
xfeed_916 0 1 tie_x0
xfeed_917 0 1 tie_x0
xfeed_918 0 1 tie_x0
xfeed_919 0 1 tie_x0
xfeed_7789 0 1 tie_x0
xfeed_7788 0 1 tie_x0
xfeed_7787 0 1 tie_x0
xfeed_7786 0 1 tie_x0
xfeed_7785 0 1 tie_x0
xfeed_7784 0 1 tie_x0
xfeed_7783 0 1 tie_x0
xfeed_7782 0 1 tie_x0
xfeed_7781 0 1 tie_x0
xfeed_7780 0 1 tie_x0
xfeed_3479 0 1 tie_x0
xfeed_3478 0 1 tie_x0
xfeed_3477 0 1 tie_x0
xfeed_3476 0 1 tie_x0
xfeed_3475 0 1 tie_x0
xfeed_3474 0 1 tie_x0
xfeed_3473 0 1 tie_x0
xfeed_3472 0 1 tie_x0
xfeed_3471 0 1 tie_x0
xfeed_3470 0 1 tie_x0
xfeed_2949 0 1 tie_x0
xfeed_2948 0 1 tie_x0
xfeed_2947 0 1 tie_x0
xfeed_2946 0 1 tie_x0
xfeed_2945 0 1 tie_x0
xfeed_2944 0 1 tie_x0
xfeed_2943 0 1 tie_x0
xfeed_2942 0 1 tie_x0
xfeed_2941 0 1 tie_x0
xfeed_2940 0 1 tie_x0
xsubckt_19_a2_x2 0 1 118 129 119 a2_x2
xfeed_920 0 1 tie_x0
xfeed_921 0 1 tie_x0
xfeed_922 0 1 tie_x0
xfeed_923 0 1 tie_x0
xfeed_924 0 1 tie_x0
xfeed_925 0 1 tie_x0
xfeed_926 0 1 tie_x0
xfeed_927 0 1 tie_x0
xfeed_928 0 1 tie_x0
xfeed_929 0 1 tie_x0
xfeed_8409 0 1 tie_x0
xfeed_8408 0 1 tie_x0
xfeed_8407 0 1 tie_x0
xfeed_8406 0 1 tie_x0
xfeed_8405 0 1 tie_x0
xfeed_8404 0 1 tie_x0
xfeed_8403 0 1 tie_x0
xfeed_8402 0 1 tie_x0
xfeed_8401 0 1 tie_x0
xfeed_8400 0 1 tie_x0
xfeed_7799 0 1 tie_x0
xfeed_7798 0 1 tie_x0
xfeed_7797 0 1 tie_x0
xfeed_7796 0 1 tie_x0
xfeed_7795 0 1 tie_x0
xfeed_7794 0 1 tie_x0
xfeed_7793 0 1 tie_x0
xfeed_7792 0 1 tie_x0
xfeed_7791 0 1 tie_x0
xfeed_7790 0 1 tie_x0
xfeed_3489 0 1 rowend_x0
xfeed_3488 0 1 tie_x0
xfeed_3487 0 1 tie_x0
xfeed_3486 0 1 tie_x0
xfeed_3485 0 1 tie_x0
xfeed_3484 0 1 tie_x0
xfeed_3483 0 1 tie_x0
xfeed_3482 0 1 tie_x0
xfeed_3481 0 1 tie_x0
xfeed_3480 0 1 tie_x0
xfeed_2959 0 1 tie_x0
xfeed_2958 0 1 tie_x0
xfeed_2957 0 1 tie_x0
xfeed_2956 0 1 tie_x0
xfeed_2955 0 1 tie_x0
xfeed_2954 0 1 tie_x0
xfeed_2953 0 1 tie_x0
xfeed_2952 0 1 tie_x0
xfeed_2951 0 1 tie_x0
xfeed_2950 0 1 tie_x0
xsubckt_59_a2_x2 0 1 212 17 11 a2_x2
xfeed_930 0 1 tie_x0
xfeed_931 0 1 tie_x0
xfeed_932 0 1 tie_x0
xfeed_933 0 1 tie_x0
xfeed_934 0 1 tie_x0
xfeed_935 0 1 tie_x0
xfeed_936 0 1 tie_x0
xfeed_937 0 1 tie_x0
xfeed_938 0 1 tie_x0
xfeed_939 0 1 tie_x0
xfeed_8419 0 1 tie_x0
xfeed_8418 0 1 tie_x0
xfeed_8417 0 1 tie_x0
xfeed_8416 0 1 tie_x0
xfeed_8415 0 1 tie_x0
xfeed_8414 0 1 tie_x0
xfeed_8413 0 1 tie_x0
xfeed_8412 0 1 tie_x0
xfeed_8411 0 1 tie_x0
xfeed_8410 0 1 tie_x0
xfeed_4109 0 1 tie_x0
xfeed_4108 0 1 tie_x0
xfeed_4107 0 1 tie_x0
xfeed_4106 0 1 tie_x0
xfeed_4105 0 1 tie_x0
xfeed_4104 0 1 tie_x0
xfeed_4103 0 1 tie_x0
xfeed_4102 0 1 tie_x0
xfeed_4101 0 1 tie_x0
xfeed_4100 0 1 tie_x0
xfeed_3499 0 1 tie_x0
xfeed_3498 0 1 tie_x0
xfeed_3497 0 1 tie_x0
xfeed_3496 0 1 tie_x0
xfeed_3495 0 1 tie_x0
xfeed_3494 0 1 tie_x0
xfeed_3493 0 1 tie_x0
xfeed_3492 0 1 tie_x0
xfeed_3491 0 1 tie_x0
xfeed_3490 0 1 tie_x0
xfeed_2969 0 1 tie_x0
xfeed_2968 0 1 tie_x0
xfeed_2967 0 1 tie_x0
xfeed_2966 0 1 rowend_x0
xfeed_2965 0 1 tie_x0
xfeed_2964 0 1 tie_x0
xfeed_2963 0 1 tie_x0
xfeed_2962 0 1 tie_x0
xfeed_2961 0 1 tie_x0
xfeed_2960 0 1 tie_x0
xfeed_940 0 1 rowend_x0
xfeed_941 0 1 tie_x0
xfeed_942 0 1 tie_x0
xfeed_943 0 1 tie_x0
xfeed_944 0 1 tie_x0
xfeed_945 0 1 tie_x0
xfeed_946 0 1 tie_x0
xfeed_947 0 1 tie_x0
xfeed_948 0 1 tie_x0
xfeed_949 0 1 tie_x0
xfeed_8429 0 1 tie_x0
xfeed_8428 0 1 tie_x0
xfeed_8427 0 1 tie_x0
xfeed_8426 0 1 tie_x0
xfeed_8425 0 1 tie_x0
xfeed_8424 0 1 tie_x0
xfeed_8423 0 1 tie_x0
xfeed_8422 0 1 tie_x0
xfeed_8421 0 1 tie_x0
xfeed_8420 0 1 tie_x0
xfeed_4119 0 1 tie_x0
xfeed_4118 0 1 tie_x0
xfeed_4117 0 1 tie_x0
xfeed_4116 0 1 tie_x0
xfeed_4115 0 1 tie_x0
xfeed_4114 0 1 tie_x0
xfeed_4113 0 1 tie_x0
xfeed_4112 0 1 tie_x0
xfeed_4111 0 1 rowend_x0
xfeed_4110 0 1 tie_x0
xfeed_2979 0 1 tie_x0
xfeed_2978 0 1 tie_x0
xfeed_2977 0 1 tie_x0
xfeed_2976 0 1 tie_x0
xfeed_2975 0 1 tie_x0
xfeed_2974 0 1 tie_x0
xfeed_2973 0 1 tie_x0
xfeed_2972 0 1 tie_x0
xfeed_2971 0 1 tie_x0
xfeed_2970 0 1 tie_x0
xsubckt_35_nao22_x1 0 1 103 107 110 112 nao22_x1
xfeed_950 0 1 tie_x0
xfeed_951 0 1 tie_x0
xfeed_952 0 1 tie_x0
xfeed_953 0 1 tie_x0
xfeed_954 0 1 tie_x0
xfeed_955 0 1 tie_x0
xfeed_956 0 1 tie_x0
xfeed_957 0 1 tie_x0
xfeed_958 0 1 tie_x0
xfeed_959 0 1 tie_x0
xfeed_8439 0 1 tie_x0
xfeed_8438 0 1 tie_x0
xfeed_8437 0 1 tie_x0
xfeed_8436 0 1 tie_x0
xfeed_8435 0 1 tie_x0
xfeed_8434 0 1 tie_x0
xfeed_8433 0 1 tie_x0
xfeed_8432 0 1 tie_x0
xfeed_8431 0 1 tie_x0
xfeed_8430 0 1 tie_x0
xfeed_7909 0 1 tie_x0
xfeed_7908 0 1 tie_x0
xfeed_7907 0 1 tie_x0
xfeed_7906 0 1 tie_x0
xfeed_7905 0 1 tie_x0
xfeed_7904 0 1 tie_x0
xfeed_7903 0 1 tie_x0
xfeed_7902 0 1 tie_x0
xfeed_7901 0 1 tie_x0
xfeed_7900 0 1 tie_x0
xfeed_4129 0 1 tie_x0
xfeed_4128 0 1 tie_x0
xfeed_4127 0 1 tie_x0
xfeed_4126 0 1 tie_x0
xfeed_4125 0 1 tie_x0
xfeed_4124 0 1 tie_x0
xfeed_4123 0 1 tie_x0
xfeed_4122 0 1 tie_x0
xfeed_4121 0 1 tie_x0
xfeed_4120 0 1 tie_x0
xfeed_2989 0 1 tie_x0
xfeed_2988 0 1 tie_x0
xfeed_2987 0 1 tie_x0
xfeed_2986 0 1 tie_x0
xfeed_2985 0 1 tie_x0
xfeed_2984 0 1 tie_x0
xfeed_2983 0 1 tie_x0
xfeed_2982 0 1 tie_x0
xfeed_2981 0 1 tie_x0
xfeed_2980 0 1 tie_x0
xsubckt_117_noa2ao222_x1 0 1 162 172 169 173 134 135 noa2ao222_x1
xsubckt_119_a2_x2 0 1 160 165 161 a2_x2
xfeed_960 0 1 tie_x0
xfeed_961 0 1 tie_x0
xfeed_962 0 1 tie_x0
xfeed_963 0 1 tie_x0
xfeed_964 0 1 tie_x0
xfeed_965 0 1 tie_x0
xfeed_966 0 1 tie_x0
xfeed_967 0 1 tie_x0
xfeed_968 0 1 tie_x0
xfeed_969 0 1 tie_x0
xfeed_8449 0 1 tie_x0
xfeed_8448 0 1 tie_x0
xfeed_8447 0 1 tie_x0
xfeed_8446 0 1 tie_x0
xfeed_8445 0 1 tie_x0
xfeed_8444 0 1 tie_x0
xfeed_8443 0 1 tie_x0
xfeed_8442 0 1 tie_x0
xfeed_8441 0 1 tie_x0
xfeed_8440 0 1 tie_x0
xfeed_7919 0 1 tie_x0
xfeed_7918 0 1 tie_x0
xfeed_7917 0 1 tie_x0
xfeed_7916 0 1 tie_x0
xfeed_7915 0 1 tie_x0
xfeed_7914 0 1 tie_x0
xfeed_7913 0 1 tie_x0
xfeed_7912 0 1 tie_x0
xfeed_7911 0 1 tie_x0
xfeed_7910 0 1 tie_x0
xfeed_4139 0 1 tie_x0
xfeed_4138 0 1 tie_x0
xfeed_4137 0 1 tie_x0
xfeed_4136 0 1 tie_x0
xfeed_4135 0 1 rowend_x0
xfeed_4134 0 1 tie_x0
xfeed_4133 0 1 tie_x0
xfeed_4132 0 1 tie_x0
xfeed_4131 0 1 tie_x0
xfeed_4130 0 1 tie_x0
xfeed_3609 0 1 tie_x0
xfeed_3608 0 1 tie_x0
xfeed_3607 0 1 tie_x0
xfeed_3606 0 1 tie_x0
xfeed_3605 0 1 tie_x0
xfeed_3604 0 1 tie_x0
xfeed_3603 0 1 tie_x0
xfeed_3602 0 1 tie_x0
xfeed_3601 0 1 tie_x0
xfeed_3600 0 1 tie_x0
xfeed_2998 0 1 tie_x0
xfeed_2997 0 1 tie_x0
xfeed_2996 0 1 tie_x0
xfeed_2995 0 1 tie_x0
xfeed_2994 0 1 tie_x0
xfeed_2993 0 1 tie_x0
xfeed_2992 0 1 tie_x0
xfeed_2991 0 1 tie_x0
xfeed_2990 0 1 tie_x0
xfeed_2999 0 1 tie_x0
xfeed_970 0 1 tie_x0
xfeed_971 0 1 tie_x0
xfeed_972 0 1 tie_x0
xfeed_973 0 1 tie_x0
xfeed_974 0 1 tie_x0
xfeed_975 0 1 tie_x0
xfeed_976 0 1 tie_x0
xfeed_977 0 1 tie_x0
xfeed_978 0 1 tie_x0
xfeed_979 0 1 tie_x0
xfeed_8459 0 1 tie_x0
xfeed_8458 0 1 tie_x0
xfeed_8457 0 1 tie_x0
xfeed_8456 0 1 tie_x0
xfeed_8455 0 1 tie_x0
xfeed_8454 0 1 tie_x0
xfeed_8453 0 1 tie_x0
xfeed_8452 0 1 tie_x0
xfeed_8451 0 1 tie_x0
xfeed_8450 0 1 tie_x0
xfeed_7929 0 1 tie_x0
xfeed_7928 0 1 tie_x0
xfeed_7927 0 1 tie_x0
xfeed_7926 0 1 tie_x0
xfeed_7925 0 1 tie_x0
xfeed_7924 0 1 tie_x0
xfeed_7923 0 1 tie_x0
xfeed_7922 0 1 tie_x0
xfeed_7921 0 1 tie_x0
xfeed_7920 0 1 tie_x0
xfeed_4149 0 1 tie_x0
xfeed_4148 0 1 tie_x0
xfeed_4147 0 1 tie_x0
xfeed_4146 0 1 tie_x0
xfeed_4145 0 1 tie_x0
xfeed_4144 0 1 tie_x0
xfeed_4143 0 1 tie_x0
xfeed_4142 0 1 tie_x0
xfeed_4141 0 1 tie_x0
xfeed_4140 0 1 tie_x0
xfeed_3619 0 1 tie_x0
xfeed_3618 0 1 tie_x0
xfeed_3617 0 1 tie_x0
xfeed_3616 0 1 tie_x0
xfeed_3615 0 1 tie_x0
xfeed_3614 0 1 tie_x0
xfeed_3613 0 1 tie_x0
xfeed_3612 0 1 tie_x0
xfeed_3611 0 1 tie_x0
xfeed_3610 0 1 tie_x0
xsubckt_162_sff1_x4 0 1 75 215 56 sff1_x4
xsubckt_158_sff1_x4 0 1 79 219 24 sff1_x4
xfeed_980 0 1 tie_x0
xfeed_981 0 1 tie_x0
xfeed_982 0 1 tie_x0
xfeed_983 0 1 tie_x0
xfeed_984 0 1 tie_x0
xfeed_985 0 1 tie_x0
xfeed_986 0 1 tie_x0
xfeed_987 0 1 tie_x0
xfeed_988 0 1 tie_x0
xfeed_989 0 1 tie_x0
xfeed_8469 0 1 tie_x0
xfeed_8468 0 1 tie_x0
xfeed_8467 0 1 tie_x0
xfeed_8466 0 1 tie_x0
xfeed_8465 0 1 tie_x0
xfeed_8464 0 1 tie_x0
xfeed_8463 0 1 tie_x0
xfeed_8462 0 1 tie_x0
xfeed_8461 0 1 tie_x0
xfeed_8460 0 1 tie_x0
xfeed_7939 0 1 tie_x0
xfeed_7938 0 1 tie_x0
xfeed_7937 0 1 tie_x0
xfeed_7936 0 1 tie_x0
xfeed_7935 0 1 tie_x0
xfeed_7934 0 1 tie_x0
xfeed_7933 0 1 tie_x0
xfeed_7932 0 1 tie_x0
xfeed_7931 0 1 tie_x0
xfeed_7930 0 1 tie_x0
xfeed_4159 0 1 tie_x0
xfeed_4158 0 1 tie_x0
xfeed_4157 0 1 tie_x0
xfeed_4156 0 1 tie_x0
xfeed_4155 0 1 tie_x0
xfeed_4154 0 1 tie_x0
xfeed_4153 0 1 tie_x0
xfeed_4152 0 1 tie_x0
xfeed_4151 0 1 tie_x0
xfeed_4150 0 1 tie_x0
xfeed_3629 0 1 tie_x0
xfeed_3628 0 1 tie_x0
xfeed_3627 0 1 tie_x0
xfeed_3626 0 1 tie_x0
xfeed_3625 0 1 tie_x0
xfeed_3624 0 1 tie_x0
xfeed_3623 0 1 tie_x0
xfeed_3622 0 1 tie_x0
xfeed_3621 0 1 tie_x0
xfeed_3620 0 1 tie_x0
xfeed_990 0 1 tie_x0
xfeed_991 0 1 tie_x0
xfeed_992 0 1 tie_x0
xfeed_993 0 1 tie_x0
xfeed_994 0 1 tie_x0
xfeed_995 0 1 tie_x0
xfeed_996 0 1 tie_x0
xfeed_997 0 1 tie_x0
xfeed_998 0 1 tie_x0
xfeed_999 0 1 tie_x0
xfeed_8479 0 1 tie_x0
xfeed_8478 0 1 tie_x0
xfeed_8477 0 1 tie_x0
xfeed_8476 0 1 tie_x0
xfeed_8475 0 1 tie_x0
xfeed_8474 0 1 rowend_x0
xfeed_8473 0 1 tie_x0
xfeed_8472 0 1 tie_x0
xfeed_8471 0 1 tie_x0
xfeed_8470 0 1 tie_x0
xfeed_7949 0 1 tie_x0
xfeed_7948 0 1 tie_x0
xfeed_7947 0 1 tie_x0
xfeed_7946 0 1 tie_x0
xfeed_7945 0 1 tie_x0
xfeed_7944 0 1 tie_x0
xfeed_7943 0 1 tie_x0
xfeed_7942 0 1 tie_x0
xfeed_7941 0 1 tie_x0
xfeed_7940 0 1 tie_x0
xfeed_4169 0 1 tie_x0
xfeed_4168 0 1 tie_x0
xfeed_4167 0 1 tie_x0
xfeed_4166 0 1 tie_x0
xfeed_4165 0 1 tie_x0
xfeed_4164 0 1 tie_x0
xfeed_4163 0 1 tie_x0
xfeed_4162 0 1 tie_x0
xfeed_4161 0 1 tie_x0
xfeed_4160 0 1 tie_x0
xfeed_3639 0 1 tie_x0
xfeed_3638 0 1 tie_x0
xfeed_3637 0 1 tie_x0
xfeed_3636 0 1 tie_x0
xfeed_3635 0 1 tie_x0
xfeed_3634 0 1 tie_x0
xfeed_3633 0 1 tie_x0
xfeed_3632 0 1 tie_x0
xfeed_3631 0 1 tie_x0
xfeed_3630 0 1 tie_x0
xfeed_8489 0 1 tie_x0
xfeed_8488 0 1 tie_x0
xfeed_8487 0 1 tie_x0
xfeed_8486 0 1 tie_x0
xfeed_8485 0 1 tie_x0
xfeed_8484 0 1 tie_x0
xfeed_8483 0 1 tie_x0
xfeed_8482 0 1 tie_x0
xfeed_8481 0 1 tie_x0
xfeed_8480 0 1 tie_x0
xfeed_7959 0 1 tie_x0
xfeed_7958 0 1 tie_x0
xfeed_7957 0 1 tie_x0
xfeed_7956 0 1 tie_x0
xfeed_7955 0 1 tie_x0
xfeed_7954 0 1 tie_x0
xfeed_7953 0 1 tie_x0
xfeed_7952 0 1 tie_x0
xfeed_7951 0 1 rowend_x0
xfeed_7950 0 1 tie_x0
xfeed_4179 0 1 tie_x0
xfeed_4178 0 1 tie_x0
xfeed_4177 0 1 tie_x0
xfeed_4176 0 1 tie_x0
xfeed_4175 0 1 tie_x0
xfeed_4174 0 1 tie_x0
xfeed_4173 0 1 tie_x0
xfeed_4172 0 1 tie_x0
xfeed_4171 0 1 tie_x0
xfeed_4170 0 1 tie_x0
xfeed_3649 0 1 tie_x0
xfeed_3648 0 1 tie_x0
xfeed_3647 0 1 tie_x0
xfeed_3646 0 1 tie_x0
xfeed_3645 0 1 tie_x0
xfeed_3644 0 1 tie_x0
xfeed_3643 0 1 tie_x0
xfeed_3642 0 1 tie_x0
xfeed_3641 0 1 tie_x0
xfeed_3640 0 1 tie_x0
xfeed_8499 0 1 tie_x0
xfeed_8498 0 1 tie_x0
xfeed_8497 0 1 tie_x0
xfeed_8496 0 1 tie_x0
xfeed_8495 0 1 tie_x0
xfeed_8494 0 1 rowend_x0
xfeed_8493 0 1 tie_x0
xfeed_8492 0 1 tie_x0
xfeed_8491 0 1 tie_x0
xfeed_8490 0 1 tie_x0
xfeed_7969 0 1 tie_x0
xfeed_7968 0 1 tie_x0
xfeed_7967 0 1 tie_x0
xfeed_7966 0 1 tie_x0
xfeed_7965 0 1 tie_x0
xfeed_7964 0 1 tie_x0
xfeed_7963 0 1 tie_x0
xfeed_7962 0 1 tie_x0
xfeed_7961 0 1 tie_x0
xfeed_7960 0 1 tie_x0
xfeed_4189 0 1 tie_x0
xfeed_4188 0 1 tie_x0
xfeed_4187 0 1 tie_x0
xfeed_4186 0 1 tie_x0
xfeed_4185 0 1 tie_x0
xfeed_4184 0 1 rowend_x0
xfeed_4183 0 1 tie_x0
xfeed_4182 0 1 tie_x0
xfeed_4181 0 1 tie_x0
xfeed_4180 0 1 tie_x0
xfeed_3659 0 1 tie_x0
xfeed_3658 0 1 tie_x0
xfeed_3657 0 1 tie_x0
xfeed_3656 0 1 tie_x0
xfeed_3655 0 1 tie_x0
xfeed_3654 0 1 tie_x0
xfeed_3653 0 1 tie_x0
xfeed_3652 0 1 tie_x0
xfeed_3651 0 1 tie_x0
xfeed_3650 0 1 tie_x0
xfeed_7977 0 1 tie_x0
xfeed_7976 0 1 tie_x0
xfeed_7975 0 1 tie_x0
xfeed_7974 0 1 tie_x0
xfeed_7973 0 1 tie_x0
xfeed_7972 0 1 tie_x0
xfeed_7971 0 1 tie_x0
xfeed_7970 0 1 tie_x0
xfeed_4199 0 1 tie_x0
xfeed_4198 0 1 tie_x0
xfeed_4197 0 1 tie_x0
xfeed_4196 0 1 tie_x0
xfeed_4195 0 1 tie_x0
xfeed_4194 0 1 tie_x0
xfeed_4193 0 1 tie_x0
xfeed_4192 0 1 tie_x0
xfeed_4191 0 1 tie_x0
xfeed_4190 0 1 tie_x0
xfeed_3669 0 1 tie_x0
xfeed_3668 0 1 tie_x0
xfeed_3667 0 1 tie_x0
xfeed_3666 0 1 tie_x0
xfeed_3665 0 1 tie_x0
xfeed_3664 0 1 tie_x0
xfeed_3663 0 1 tie_x0
xfeed_3662 0 1 tie_x0
xfeed_3661 0 1 tie_x0
xfeed_3660 0 1 tie_x0
xsubckt_10_a2_x2 0 1 126 128 127 a2_x2
xfeed_7979 0 1 tie_x0
xfeed_7978 0 1 tie_x0
xsubckt_70_a2_x2 0 1 201 91 203 a2_x2
xsubckt_30_a2_x2 0 1 108 13 16 a2_x2
xfeed_7984 0 1 tie_x0
xfeed_7983 0 1 tie_x0
xfeed_7982 0 1 tie_x0
xfeed_7981 0 1 tie_x0
xfeed_7980 0 1 tie_x0
xfeed_3679 0 1 tie_x0
xfeed_3678 0 1 tie_x0
xfeed_3677 0 1 tie_x0
xfeed_3676 0 1 tie_x0
xfeed_3675 0 1 tie_x0
xfeed_3674 0 1 tie_x0
xfeed_3673 0 1 tie_x0
xfeed_3672 0 1 tie_x0
xfeed_3671 0 1 rowend_x0
xfeed_3670 0 1 tie_x0
xsubckt_90_a2_x2 0 1 183 188 184 a2_x2
xsubckt_94_on12_x1 0 1 180 3 2 on12_x1
xfeed_7989 0 1 tie_x0
xfeed_7988 0 1 tie_x0
xfeed_7987 0 1 tie_x0
xfeed_7986 0 1 tie_x0
xfeed_7985 0 1 tie_x0
xfeed_8609 0 1 tie_x0
xfeed_8608 0 1 tie_x0
xfeed_8607 0 1 tie_x0
xfeed_8606 0 1 tie_x0
xfeed_8605 0 1 tie_x0
xfeed_8604 0 1 tie_x0
xfeed_8603 0 1 tie_x0
xfeed_8602 0 1 tie_x0
xfeed_8601 0 1 tie_x0
xfeed_8600 0 1 tie_x0
xfeed_7991 0 1 tie_x0
xfeed_7990 0 1 tie_x0
xfeed_3689 0 1 tie_x0
xfeed_3688 0 1 tie_x0
xfeed_3687 0 1 tie_x0
xfeed_3686 0 1 tie_x0
xfeed_3685 0 1 tie_x0
xfeed_3684 0 1 tie_x0
xfeed_3683 0 1 tie_x0
xfeed_3682 0 1 tie_x0
xfeed_3681 0 1 tie_x0
xfeed_3680 0 1 tie_x0
xfeed_7999 0 1 tie_x0
xfeed_7998 0 1 tie_x0
xfeed_7997 0 1 tie_x0
xfeed_7996 0 1 tie_x0
xfeed_7995 0 1 tie_x0
xfeed_7994 0 1 tie_x0
xfeed_7993 0 1 tie_x0
xfeed_7992 0 1 tie_x0
xfeed_8619 0 1 tie_x0
xfeed_8618 0 1 tie_x0
xfeed_8617 0 1 tie_x0
xfeed_8616 0 1 tie_x0
xfeed_8615 0 1 tie_x0
xfeed_8614 0 1 tie_x0
xfeed_8613 0 1 tie_x0
xfeed_8612 0 1 tie_x0
xfeed_8611 0 1 tie_x0
xfeed_8610 0 1 tie_x0
xfeed_4309 0 1 tie_x0
xfeed_4308 0 1 tie_x0
xfeed_4307 0 1 tie_x0
xfeed_4306 0 1 tie_x0
xfeed_4305 0 1 tie_x0
xfeed_4304 0 1 tie_x0
xfeed_4303 0 1 tie_x0
xfeed_4302 0 1 tie_x0
xfeed_4301 0 1 tie_x0
xfeed_4300 0 1 tie_x0
xfeed_3698 0 1 tie_x0
xfeed_3697 0 1 rowend_x0
xfeed_3696 0 1 tie_x0
xfeed_3695 0 1 tie_x0
xfeed_3694 0 1 tie_x0
xfeed_3693 0 1 tie_x0
xfeed_3692 0 1 tie_x0
xfeed_3691 0 1 tie_x0
xfeed_3690 0 1 tie_x0
xfeed_3699 0 1 tie_x0
xsubckt_39_nao22_x1 0 1 99 114 106 104 nao22_x1
xfeed_8629 0 1 tie_x0
xfeed_8628 0 1 tie_x0
xfeed_8627 0 1 tie_x0
xfeed_8626 0 1 tie_x0
xfeed_8625 0 1 tie_x0
xfeed_8624 0 1 tie_x0
xfeed_8623 0 1 tie_x0
xfeed_8622 0 1 tie_x0
xfeed_8621 0 1 tie_x0
xfeed_8620 0 1 tie_x0
xfeed_4319 0 1 tie_x0
xfeed_4318 0 1 tie_x0
xfeed_4317 0 1 tie_x0
xfeed_4316 0 1 tie_x0
xfeed_4315 0 1 rowend_x0
xfeed_4314 0 1 tie_x0
xfeed_4313 0 1 tie_x0
xfeed_4312 0 1 tie_x0
xfeed_4311 0 1 tie_x0
xfeed_4310 0 1 tie_x0
xsubckt_110_a2_x2 0 1 219 131 168 a2_x2
xfeed_8639 0 1 tie_x0
xfeed_8638 0 1 tie_x0
xfeed_8637 0 1 tie_x0
xfeed_8636 0 1 tie_x0
xfeed_8635 0 1 tie_x0
xfeed_8634 0 1 tie_x0
xfeed_8633 0 1 tie_x0
xfeed_8632 0 1 tie_x0
xfeed_8631 0 1 tie_x0
xfeed_8630 0 1 tie_x0
xfeed_4329 0 1 tie_x0
xfeed_4328 0 1 tie_x0
xfeed_4327 0 1 tie_x0
xfeed_4326 0 1 tie_x0
xfeed_4325 0 1 tie_x0
xfeed_4324 0 1 tie_x0
xfeed_4323 0 1 tie_x0
xfeed_4322 0 1 tie_x0
xfeed_4321 0 1 tie_x0
xfeed_4320 0 1 tie_x0
xsubckt_145_ao22_x2 0 1 137 138 142 146 ao22_x2
xsubckt_86_a4_x2 0 1 187 12 16 11 15 a4_x2
xfeed_8649 0 1 tie_x0
xfeed_8648 0 1 tie_x0
xfeed_8647 0 1 tie_x0
xfeed_8646 0 1 tie_x0
xfeed_8645 0 1 tie_x0
xfeed_8644 0 1 tie_x0
xfeed_8643 0 1 tie_x0
xfeed_8642 0 1 tie_x0
xfeed_8641 0 1 tie_x0
xfeed_8640 0 1 tie_x0
xfeed_4339 0 1 rowend_x0
xfeed_4338 0 1 tie_x0
xfeed_4337 0 1 tie_x0
xfeed_4336 0 1 tie_x0
xfeed_4335 0 1 tie_x0
xfeed_4334 0 1 tie_x0
xfeed_4333 0 1 tie_x0
xfeed_4332 0 1 tie_x0
xfeed_4331 0 1 tie_x0
xfeed_4330 0 1 tie_x0
xfeed_3809 0 1 tie_x0
xfeed_3808 0 1 tie_x0
xfeed_3807 0 1 tie_x0
xfeed_3806 0 1 tie_x0
xfeed_3805 0 1 tie_x0
xfeed_3804 0 1 tie_x0
xfeed_3803 0 1 tie_x0
xfeed_3802 0 1 tie_x0
xfeed_3801 0 1 tie_x0
xfeed_3800 0 1 tie_x0
xsubckt_65_nxr2_x1 0 1 206 84 210 nxr2_x1
xfeed_8659 0 1 tie_x0
xfeed_8658 0 1 tie_x0
xfeed_8657 0 1 tie_x0
xfeed_8656 0 1 tie_x0
xfeed_8655 0 1 tie_x0
xfeed_8654 0 1 tie_x0
xfeed_8653 0 1 tie_x0
xfeed_8652 0 1 tie_x0
xfeed_8651 0 1 tie_x0
xfeed_8650 0 1 tie_x0
xfeed_4349 0 1 tie_x0
xfeed_4348 0 1 tie_x0
xfeed_4347 0 1 tie_x0
xfeed_4346 0 1 tie_x0
xfeed_4345 0 1 tie_x0
xfeed_4344 0 1 tie_x0
xfeed_4343 0 1 tie_x0
xfeed_4342 0 1 tie_x0
xfeed_4341 0 1 tie_x0
xfeed_4340 0 1 tie_x0
xfeed_3819 0 1 tie_x0
xfeed_3818 0 1 tie_x0
xfeed_3817 0 1 tie_x0
xfeed_3816 0 1 tie_x0
xfeed_3815 0 1 tie_x0
xfeed_3814 0 1 tie_x0
xfeed_3813 0 1 tie_x0
xfeed_3812 0 1 tie_x0
xfeed_3811 0 1 tie_x0
xfeed_3810 0 1 tie_x0
xsubckt_126_an12_x1 0 1 154 158 156 an12_x1
xfeed_8669 0 1 tie_x0
xfeed_8668 0 1 tie_x0
xfeed_8667 0 1 tie_x0
xfeed_8666 0 1 tie_x0
xfeed_8665 0 1 tie_x0
xfeed_8664 0 1 tie_x0
xfeed_8663 0 1 tie_x0
xfeed_8662 0 1 tie_x0
xfeed_8661 0 1 tie_x0
xfeed_8660 0 1 tie_x0
xfeed_4359 0 1 tie_x0
xfeed_4358 0 1 tie_x0
xfeed_4357 0 1 tie_x0
xfeed_4356 0 1 tie_x0
xfeed_4355 0 1 tie_x0
xfeed_4354 0 1 tie_x0
xfeed_4353 0 1 tie_x0
xfeed_4352 0 1 tie_x0
xfeed_4351 0 1 tie_x0
xfeed_4350 0 1 tie_x0
xfeed_3829 0 1 tie_x0
xfeed_3828 0 1 tie_x0
xfeed_3827 0 1 tie_x0
xfeed_3826 0 1 tie_x0
xfeed_3825 0 1 tie_x0
xfeed_3824 0 1 tie_x0
xfeed_3823 0 1 tie_x0
xfeed_3822 0 1 tie_x0
xfeed_3821 0 1 tie_x0
xfeed_3820 0 1 tie_x0
xfeed_8677 0 1 tie_x0
xfeed_8676 0 1 tie_x0
xfeed_8675 0 1 tie_x0
xfeed_8674 0 1 tie_x0
xfeed_8673 0 1 tie_x0
xfeed_8672 0 1 tie_x0
xfeed_8671 0 1 tie_x0
xfeed_8670 0 1 tie_x0
xfeed_4369 0 1 tie_x0
xfeed_4368 0 1 tie_x0
xfeed_4367 0 1 tie_x0
xfeed_4366 0 1 tie_x0
xfeed_4365 0 1 rowend_x0
xfeed_4364 0 1 tie_x0
xfeed_4363 0 1 tie_x0
xfeed_4362 0 1 tie_x0
xfeed_4361 0 1 tie_x0
xfeed_4360 0 1 tie_x0
xfeed_3838 0 1 tie_x0
xfeed_3837 0 1 tie_x0
xfeed_3836 0 1 tie_x0
xfeed_3835 0 1 tie_x0
xfeed_3834 0 1 tie_x0
xfeed_3833 0 1 tie_x0
xfeed_3832 0 1 tie_x0
xfeed_3831 0 1 tie_x0
xfeed_3830 0 1 tie_x0
xfeed_8679 0 1 tie_x0
xfeed_8678 0 1 tie_x0
xfeed_3839 0 1 tie_x0
xfeed_8684 0 1 tie_x0
xfeed_8683 0 1 tie_x0
xfeed_8682 0 1 rowend_x0
xfeed_8681 0 1 tie_x0
xfeed_8680 0 1 tie_x0
xfeed_4379 0 1 tie_x0
xfeed_4378 0 1 tie_x0
xfeed_4377 0 1 tie_x0
xfeed_4376 0 1 tie_x0
xfeed_4375 0 1 tie_x0
xfeed_4374 0 1 tie_x0
xfeed_4373 0 1 tie_x0
xfeed_4372 0 1 tie_x0
xfeed_4371 0 1 tie_x0
xfeed_4370 0 1 tie_x0
xfeed_3845 0 1 tie_x0
xfeed_3844 0 1 tie_x0
xfeed_3843 0 1 tie_x0
xfeed_3842 0 1 tie_x0
xfeed_3841 0 1 tie_x0
xfeed_3840 0 1 tie_x0
xsubckt_127_a2_x2 0 1 153 76 5 a2_x2
xfeed_8689 0 1 tie_x0
xfeed_8688 0 1 tie_x0
xfeed_8687 0 1 tie_x0
xfeed_8686 0 1 tie_x0
xfeed_8685 0 1 tie_x0
xfeed_3849 0 1 tie_x0
xfeed_3848 0 1 tie_x0
xfeed_3847 0 1 tie_x0
xfeed_3846 0 1 tie_x0
xfeed_8691 0 1 tie_x0
xfeed_8690 0 1 tie_x0
xfeed_4389 0 1 tie_x0
xfeed_4388 0 1 tie_x0
xfeed_4387 0 1 tie_x0
xfeed_4386 0 1 tie_x0
xfeed_4385 0 1 tie_x0
xfeed_4384 0 1 tie_x0
xfeed_4383 0 1 tie_x0
xfeed_4382 0 1 tie_x0
xfeed_4381 0 1 tie_x0
xfeed_4380 0 1 tie_x0
xfeed_3852 0 1 tie_x0
xfeed_3851 0 1 tie_x0
xfeed_3850 0 1 tie_x0
xsubckt_32_a3_x2 0 1 106 111 109 108 a3_x2
xfeed_8699 0 1 tie_x0
xfeed_8698 0 1 tie_x0
xfeed_8697 0 1 tie_x0
xfeed_8696 0 1 tie_x0
xfeed_8695 0 1 tie_x0
xfeed_8694 0 1 tie_x0
xfeed_8693 0 1 tie_x0
xfeed_8692 0 1 tie_x0
xfeed_3859 0 1 tie_x0
xfeed_3858 0 1 tie_x0
xfeed_3857 0 1 tie_x0
xfeed_3856 0 1 tie_x0
xfeed_3855 0 1 tie_x0
xfeed_3854 0 1 tie_x0
xfeed_3853 0 1 tie_x0
xfeed_5009 0 1 tie_x0
xfeed_5008 0 1 tie_x0
xfeed_5007 0 1 tie_x0
xfeed_5006 0 1 tie_x0
xfeed_5005 0 1 tie_x0
xfeed_5004 0 1 tie_x0
xfeed_5003 0 1 tie_x0
xfeed_5002 0 1 tie_x0
xfeed_5001 0 1 tie_x0
xfeed_5000 0 1 tie_x0
xfeed_4398 0 1 tie_x0
xfeed_4397 0 1 tie_x0
xfeed_4396 0 1 tie_x0
xfeed_4395 0 1 tie_x0
xfeed_4394 0 1 tie_x0
xfeed_4393 0 1 tie_x0
xfeed_4392 0 1 tie_x0
xfeed_4391 0 1 tie_x0
xfeed_4390 0 1 tie_x0
xfeed_4399 0 1 tie_x0
xfeed_3869 0 1 tie_x0
xfeed_3868 0 1 tie_x0
xfeed_3867 0 1 tie_x0
xfeed_3866 0 1 tie_x0
xfeed_3865 0 1 tie_x0
xfeed_3864 0 1 tie_x0
xfeed_3863 0 1 tie_x0
xfeed_3862 0 1 tie_x0
xfeed_3861 0 1 tie_x0
xfeed_3860 0 1 tie_x0
xspare_buffer_8 0 1 57 71 buf_x8
xspare_buffer_4 0 1 70 71 buf_x8
xspare_buffer_0 0 1 71 72 buf_x8
xfeed_5019 0 1 tie_x0
xfeed_5018 0 1 tie_x0
xfeed_5017 0 1 tie_x0
xfeed_5016 0 1 tie_x0
xfeed_5015 0 1 tie_x0
xfeed_5014 0 1 tie_x0
xfeed_5013 0 1 tie_x0
xfeed_5012 0 1 tie_x0
xfeed_5011 0 1 rowend_x0
xfeed_5010 0 1 tie_x0
xfeed_3879 0 1 tie_x0
xfeed_3878 0 1 tie_x0
xfeed_3877 0 1 rowend_x0
xfeed_3876 0 1 tie_x0
xfeed_3875 0 1 tie_x0
xfeed_3874 0 1 tie_x0
xfeed_3873 0 1 tie_x0
xfeed_3872 0 1 tie_x0
xfeed_3871 0 1 tie_x0
xfeed_3870 0 1 tie_x0
xsubckt_118_oa2ao222_x2 0 1 161 172 169 173 134 135 oa2ao222_x2
xfeed_5029 0 1 tie_x0
xfeed_5028 0 1 tie_x0
xfeed_5027 0 1 tie_x0
xfeed_5026 0 1 tie_x0
xfeed_5025 0 1 tie_x0
xfeed_5024 0 1 tie_x0
xfeed_5023 0 1 tie_x0
xfeed_5022 0 1 tie_x0
xfeed_5021 0 1 tie_x0
xfeed_5020 0 1 tie_x0
xsubckt_100_no2_x1 0 1 176 80 9 no2_x1
xfeed_3889 0 1 tie_x0
xfeed_3888 0 1 tie_x0
xfeed_3887 0 1 tie_x0
xfeed_3886 0 1 tie_x0
xfeed_3885 0 1 tie_x0
xfeed_3884 0 1 tie_x0
xfeed_3883 0 1 tie_x0
xfeed_3882 0 1 tie_x0
xfeed_3881 0 1 tie_x0
xfeed_3880 0 1 tie_x0
xsubckt_106_no2_x1 0 1 171 79 8 no2_x1
xfeed_5039 0 1 tie_x0
xfeed_5038 0 1 tie_x0
xfeed_5037 0 1 tie_x0
xfeed_5036 0 1 rowend_x0
xfeed_5035 0 1 tie_x0
xfeed_5034 0 1 tie_x0
xfeed_5033 0 1 tie_x0
xfeed_5032 0 1 tie_x0
xfeed_5031 0 1 tie_x0
xfeed_5030 0 1 tie_x0
xfeed_4509 0 1 tie_x0
xfeed_4508 0 1 tie_x0
xfeed_4507 0 1 tie_x0
xfeed_4506 0 1 tie_x0
xfeed_4505 0 1 tie_x0
xfeed_4504 0 1 tie_x0
xfeed_4503 0 1 tie_x0
xfeed_4502 0 1 tie_x0
xfeed_4501 0 1 tie_x0
xfeed_4500 0 1 tie_x0
xfeed_3899 0 1 tie_x0
xfeed_3898 0 1 tie_x0
xfeed_3897 0 1 tie_x0
xfeed_3896 0 1 tie_x0
xfeed_3895 0 1 tie_x0
xfeed_3894 0 1 tie_x0
xfeed_3893 0 1 tie_x0
xfeed_3892 0 1 tie_x0
xfeed_3891 0 1 tie_x0
xfeed_3890 0 1 tie_x0
xsubckt_111_ao22_x2 0 1 167 172 171 173 ao22_x2
xfeed_5049 0 1 tie_x0
xfeed_5048 0 1 tie_x0
xfeed_5047 0 1 tie_x0
xfeed_5046 0 1 tie_x0
xfeed_5045 0 1 tie_x0
xfeed_5044 0 1 tie_x0
xfeed_5043 0 1 tie_x0
xfeed_5042 0 1 tie_x0
xfeed_5041 0 1 tie_x0
xfeed_5040 0 1 tie_x0
xfeed_4519 0 1 rowend_x0
xfeed_4518 0 1 tie_x0
xfeed_4517 0 1 tie_x0
xfeed_4516 0 1 tie_x0
xfeed_4515 0 1 tie_x0
xfeed_4514 0 1 tie_x0
xfeed_4513 0 1 tie_x0
xfeed_4512 0 1 tie_x0
xfeed_4511 0 1 tie_x0
xfeed_4510 0 1 tie_x0
xspare_feed_13 0 1 tie_x0
xspare_feed_12 0 1 tie_x0
xspare_feed_11 0 1 tie_x0
xspare_feed_10 0 1 tie_x0
xspare_feed_19 0 1 tie_x0
xspare_feed_18 0 1 tie_x0
xspare_feed_17 0 1 tie_x0
xspare_feed_16 0 1 tie_x0
xspare_feed_15 0 1 tie_x0
xspare_feed_14 0 1 tie_x0
xfeed_5059 0 1 tie_x0
xfeed_5058 0 1 tie_x0
xfeed_5057 0 1 tie_x0
xfeed_5056 0 1 tie_x0
xfeed_5055 0 1 tie_x0
xfeed_5054 0 1 tie_x0
xfeed_5053 0 1 tie_x0
xfeed_5052 0 1 tie_x0
xfeed_5051 0 1 tie_x0
xfeed_5050 0 1 tie_x0
xfeed_4529 0 1 tie_x0
xfeed_4528 0 1 tie_x0
xfeed_4527 0 1 tie_x0
xfeed_4526 0 1 tie_x0
xfeed_4525 0 1 tie_x0
xfeed_4524 0 1 tie_x0
xfeed_4523 0 1 rowend_x0
xfeed_4522 0 1 tie_x0
xfeed_4521 0 1 tie_x0
xfeed_4520 0 1 tie_x0
xspare_feed_20 0 1 tie_x0
xsubckt_49_a3_x2 0 1 89 131 92 90 a3_x2
xspare_feed_29 0 1 tie_x0
xspare_feed_28 0 1 tie_x0
xspare_feed_27 0 1 tie_x0
xspare_feed_26 0 1 tie_x0
xspare_feed_25 0 1 tie_x0
xspare_feed_24 0 1 tie_x0
xspare_feed_23 0 1 tie_x0
xspare_feed_22 0 1 tie_x0
xspare_feed_21 0 1 tie_x0
xfeed_5069 0 1 tie_x0
xfeed_5068 0 1 tie_x0
xfeed_5067 0 1 tie_x0
xfeed_5066 0 1 tie_x0
xfeed_5065 0 1 tie_x0
xfeed_5064 0 1 tie_x0
xfeed_5063 0 1 tie_x0
xfeed_5062 0 1 tie_x0
xfeed_5061 0 1 tie_x0
xfeed_5060 0 1 tie_x0
xfeed_4538 0 1 tie_x0
xfeed_4537 0 1 tie_x0
xfeed_4536 0 1 tie_x0
xfeed_4535 0 1 tie_x0
xfeed_4534 0 1 tie_x0
xfeed_4533 0 1 tie_x0
xfeed_4532 0 1 tie_x0
xfeed_4531 0 1 tie_x0
xfeed_4530 0 1 tie_x0
xspare_feed_9 0 1 tie_x0
xspare_feed_8 0 1 tie_x0
xspare_feed_7 0 1 tie_x0
xspare_feed_6 0 1 tie_x0
xspare_feed_5 0 1 tie_x0
xspare_feed_4 0 1 tie_x0
xspare_feed_3 0 1 tie_x0
xspare_feed_2 0 1 tie_x0
xspare_feed_1 0 1 tie_x0
xspare_feed_0 0 1 tie_x0
xfeed_4539 0 1 tie_x0
xspare_feed_39 0 1 tie_x0
xspare_feed_38 0 1 tie_x0
xspare_feed_37 0 1 tie_x0
xspare_feed_36 0 1 tie_x0
xspare_feed_35 0 1 tie_x0
xspare_feed_34 0 1 tie_x0
xspare_feed_33 0 1 tie_x0
xspare_feed_32 0 1 tie_x0
xspare_feed_31 0 1 tie_x0
xspare_feed_30 0 1 tie_x0
xfeed_5079 0 1 tie_x0
xfeed_5078 0 1 tie_x0
xfeed_5077 0 1 tie_x0
xfeed_5076 0 1 tie_x0
xfeed_5075 0 1 tie_x0
xfeed_5074 0 1 tie_x0
xfeed_5073 0 1 tie_x0
xfeed_5072 0 1 tie_x0
xfeed_5071 0 1 tie_x0
xfeed_5070 0 1 tie_x0
xfeed_4545 0 1 tie_x0
xfeed_4544 0 1 tie_x0
xfeed_4543 0 1 tie_x0
xfeed_4542 0 1 tie_x0
xfeed_4541 0 1 tie_x0
xfeed_4540 0 1 tie_x0
xfeed_4549 0 1 tie_x0
xfeed_4548 0 1 tie_x0
xfeed_4547 0 1 tie_x0
xfeed_4546 0 1 tie_x0
xspare_feed_49 0 1 tie_x0
xspare_feed_48 0 1 tie_x0
xspare_feed_47 0 1 tie_x0
xspare_feed_46 0 1 tie_x0
xspare_feed_45 0 1 tie_x0
xspare_feed_44 0 1 tie_x0
xspare_feed_43 0 1 tie_x0
xspare_feed_42 0 1 tie_x0
xspare_feed_41 0 1 tie_x0
xspare_feed_40 0 1 tie_x0
xfeed_5089 0 1 tie_x0
xfeed_5088 0 1 tie_x0
xfeed_5087 0 1 tie_x0
xfeed_5086 0 1 tie_x0
xfeed_5085 0 1 tie_x0
xfeed_5084 0 1 tie_x0
xfeed_5083 0 1 tie_x0
xfeed_5082 0 1 tie_x0
xfeed_5081 0 1 tie_x0
xfeed_5080 0 1 tie_x0
xfeed_4552 0 1 tie_x0
xfeed_4551 0 1 tie_x0
xfeed_4550 0 1 tie_x0
xfeed_4559 0 1 tie_x0
xfeed_4558 0 1 tie_x0
xfeed_4557 0 1 tie_x0
xfeed_4556 0 1 tie_x0
xfeed_4555 0 1 tie_x0
xfeed_4554 0 1 tie_x0
xfeed_4553 0 1 tie_x0
xspare_feed_59 0 1 tie_x0
xspare_feed_58 0 1 tie_x0
xspare_feed_57 0 1 tie_x0
xspare_feed_56 0 1 tie_x0
xspare_feed_55 0 1 tie_x0
xspare_feed_54 0 1 tie_x0
xspare_feed_53 0 1 tie_x0
xspare_feed_52 0 1 tie_x0
xspare_feed_51 0 1 tie_x0
xspare_feed_50 0 1 tie_x0
xfeed_5098 0 1 tie_x0
xfeed_5097 0 1 tie_x0
xfeed_5096 0 1 tie_x0
xfeed_5095 0 1 tie_x0
xfeed_5094 0 1 tie_x0
xfeed_5093 0 1 tie_x0
xfeed_5092 0 1 tie_x0
xfeed_5091 0 1 tie_x0
xfeed_5090 0 1 tie_x0
xfeed_5099 0 1 tie_x0
xfeed_4569 0 1 tie_x0
xfeed_4568 0 1 tie_x0
xfeed_4567 0 1 tie_x0
xfeed_4566 0 1 tie_x0
xfeed_4565 0 1 tie_x0
xfeed_4564 0 1 tie_x0
xfeed_4563 0 1 tie_x0
xfeed_4562 0 1 tie_x0
xfeed_4561 0 1 tie_x0
xfeed_4560 0 1 tie_x0
xspare_feed_69 0 1 tie_x0
xspare_feed_68 0 1 tie_x0
xspare_feed_67 0 1 tie_x0
xspare_feed_66 0 1 tie_x0
xspare_feed_65 0 1 tie_x0
xspare_feed_64 0 1 tie_x0
xspare_feed_63 0 1 tie_x0
xspare_feed_62 0 1 tie_x0
xspare_feed_61 0 1 tie_x0
xspare_feed_60 0 1 tie_x0
xsubckt_13_na2_x1 0 1 124 13 17 na2_x1
xfeed_4579 0 1 tie_x0
xfeed_4578 0 1 tie_x0
xfeed_4577 0 1 tie_x0
xfeed_4576 0 1 tie_x0
xfeed_4575 0 1 tie_x0
xfeed_4574 0 1 tie_x0
xfeed_4573 0 1 tie_x0
xfeed_4572 0 1 tie_x0
xfeed_4571 0 1 tie_x0
xfeed_4570 0 1 tie_x0
xspare_feed_78 0 1 tie_x0
xspare_feed_77 0 1 tie_x0
xspare_feed_76 0 1 tie_x0
xspare_feed_75 0 1 tie_x0
xspare_feed_74 0 1 tie_x0
xspare_feed_73 0 1 tie_x0
xspare_feed_72 0 1 tie_x0
xspare_feed_71 0 1 tie_x0
xspare_feed_70 0 1 tie_x0
xspare_feed_79 0 1 tie_x0
xfeed_4589 0 1 tie_x0
xfeed_4588 0 1 tie_x0
xfeed_4587 0 1 tie_x0
xfeed_4586 0 1 tie_x0
xfeed_4585 0 1 tie_x0
xfeed_4584 0 1 tie_x0
xfeed_4583 0 1 tie_x0
xfeed_4582 0 1 tie_x0
xfeed_4581 0 1 tie_x0
xfeed_4580 0 1 tie_x0
xspare_feed_80 0 1 tie_x0
xspare_feed_81 0 1 tie_x0
xspare_feed_82 0 1 tie_x0
xspare_feed_83 0 1 tie_x0
xspare_feed_84 0 1 tie_x0
xspare_feed_85 0 1 rowend_x0
xspare_feed_86 0 1 tie_x0
xspare_feed_87 0 1 rowend_x0
xspare_feed_88 0 1 rowend_x0
xspare_feed_89 0 1 tie_x0
xfeed_5209 0 1 tie_x0
xfeed_5208 0 1 tie_x0
xfeed_5207 0 1 tie_x0
xfeed_5206 0 1 tie_x0
xfeed_5205 0 1 tie_x0
xfeed_5204 0 1 tie_x0
xfeed_5203 0 1 tie_x0
xfeed_5202 0 1 tie_x0
xfeed_5201 0 1 tie_x0
xfeed_5200 0 1 tie_x0
xfeed_4599 0 1 tie_x0
xfeed_4598 0 1 tie_x0
xfeed_4597 0 1 tie_x0
xfeed_4596 0 1 tie_x0
xfeed_4595 0 1 tie_x0
xfeed_4594 0 1 tie_x0
xfeed_4593 0 1 tie_x0
xfeed_4592 0 1 tie_x0
xfeed_4591 0 1 tie_x0
xfeed_4590 0 1 tie_x0
xspare_feed_90 0 1 rowend_x0
xspare_feed_91 0 1 tie_x0
xspare_feed_92 0 1 rowend_x0
xspare_feed_93 0 1 rowend_x0
xspare_feed_94 0 1 tie_x0
xspare_feed_95 0 1 rowend_x0
xspare_feed_96 0 1 tie_x0
xspare_feed_97 0 1 rowend_x0
xspare_feed_98 0 1 rowend_x0
xspare_feed_99 0 1 tie_x0
xfeed_5219 0 1 tie_x0
xfeed_5218 0 1 tie_x0
xfeed_5217 0 1 tie_x0
xfeed_5216 0 1 tie_x0
xfeed_5215 0 1 tie_x0
xfeed_5214 0 1 tie_x0
xfeed_5213 0 1 tie_x0
xfeed_5212 0 1 tie_x0
xfeed_5211 0 1 tie_x0
xfeed_5210 0 1 tie_x0
xfeed_5229 0 1 tie_x0
xfeed_5228 0 1 tie_x0
xfeed_5227 0 1 tie_x0
xfeed_5226 0 1 tie_x0
xfeed_5225 0 1 tie_x0
xfeed_5224 0 1 tie_x0
xfeed_5223 0 1 tie_x0
xfeed_5222 0 1 tie_x0
xfeed_5221 0 1 tie_x0
xfeed_5220 0 1 tie_x0
xfeed_5238 0 1 tie_x0
xfeed_5237 0 1 tie_x0
xfeed_5236 0 1 tie_x0
xfeed_5235 0 1 tie_x0
xfeed_5234 0 1 tie_x0
xfeed_5233 0 1 tie_x0
xfeed_5232 0 1 tie_x0
xfeed_5231 0 1 tie_x0
xfeed_5230 0 1 tie_x0
xsubckt_87_na4_x1 0 1 186 12 16 11 15 na4_x1
xsubckt_135_a2_x2 0 1 146 75 4 a2_x2
xfeed_5239 0 1 tie_x0
xfeed_4709 0 1 tie_x0
xfeed_4708 0 1 tie_x0
xfeed_4707 0 1 tie_x0
xfeed_4706 0 1 tie_x0
xfeed_4705 0 1 tie_x0
xfeed_4704 0 1 tie_x0
xfeed_4703 0 1 tie_x0
xfeed_4702 0 1 tie_x0
xfeed_4701 0 1 tie_x0
xfeed_4700 0 1 tie_x0
xsubckt_147_ao22_x2 0 1 214 131 137 136 ao22_x2
xfeed_5245 0 1 tie_x0
xfeed_5244 0 1 tie_x0
xfeed_5243 0 1 tie_x0
xfeed_5242 0 1 tie_x0
xfeed_5241 0 1 tie_x0
xfeed_5240 0 1 tie_x0
xfeed_5249 0 1 tie_x0
xfeed_5248 0 1 tie_x0
xfeed_5247 0 1 tie_x0
xfeed_5246 0 1 tie_x0
xfeed_4719 0 1 tie_x0
xfeed_4718 0 1 tie_x0
xfeed_4717 0 1 tie_x0
xfeed_4716 0 1 tie_x0
xfeed_4715 0 1 tie_x0
xfeed_4714 0 1 tie_x0
xfeed_4713 0 1 tie_x0
xfeed_4712 0 1 tie_x0
xfeed_4711 0 1 tie_x0
xfeed_4710 0 1 tie_x0
xfeed_5252 0 1 tie_x0
xfeed_5251 0 1 tie_x0
xfeed_5250 0 1 tie_x0
xfeed_5259 0 1 tie_x0
xfeed_5258 0 1 tie_x0
xfeed_5257 0 1 tie_x0
xfeed_5256 0 1 tie_x0
xfeed_5255 0 1 tie_x0
xfeed_5254 0 1 tie_x0
xfeed_5253 0 1 tie_x0
xfeed_4729 0 1 tie_x0
xfeed_4728 0 1 tie_x0
xfeed_4727 0 1 tie_x0
xfeed_4726 0 1 tie_x0
xfeed_4725 0 1 rowend_x0
xfeed_4724 0 1 tie_x0
xfeed_4723 0 1 tie_x0
xfeed_4722 0 1 tie_x0
xfeed_4721 0 1 tie_x0
xfeed_4720 0 1 tie_x0
xfeed_5269 0 1 tie_x0
xfeed_5268 0 1 tie_x0
xfeed_5267 0 1 tie_x0
xfeed_5266 0 1 tie_x0
xfeed_5265 0 1 tie_x0
xfeed_5264 0 1 tie_x0
xfeed_5263 0 1 tie_x0
xfeed_5262 0 1 tie_x0
xfeed_5261 0 1 tie_x0
xfeed_5260 0 1 tie_x0
xfeed_4739 0 1 tie_x0
xfeed_4738 0 1 tie_x0
xfeed_4737 0 1 tie_x0
xfeed_4736 0 1 tie_x0
xfeed_4735 0 1 tie_x0
xfeed_4734 0 1 tie_x0
xfeed_4733 0 1 tie_x0
xfeed_4732 0 1 tie_x0
xfeed_4731 0 1 tie_x0
xfeed_4730 0 1 tie_x0
xfeed_5279 0 1 tie_x0
xfeed_5278 0 1 tie_x0
xfeed_5277 0 1 tie_x0
xfeed_5276 0 1 tie_x0
xfeed_5275 0 1 tie_x0
xfeed_5274 0 1 tie_x0
xfeed_5273 0 1 tie_x0
xfeed_5272 0 1 tie_x0
xfeed_5271 0 1 tie_x0
xfeed_5270 0 1 tie_x0
xfeed_4749 0 1 tie_x0
xfeed_4748 0 1 tie_x0
xfeed_4747 0 1 tie_x0
xfeed_4746 0 1 tie_x0
xfeed_4745 0 1 tie_x0
xfeed_4744 0 1 tie_x0
xfeed_4743 0 1 tie_x0
xfeed_4742 0 1 tie_x0
xfeed_4741 0 1 tie_x0
xfeed_4740 0 1 tie_x0
xfeed_5289 0 1 tie_x0
xfeed_5288 0 1 tie_x0
xfeed_5287 0 1 tie_x0
xfeed_5286 0 1 tie_x0
xfeed_5285 0 1 tie_x0
xfeed_5284 0 1 tie_x0
xfeed_5283 0 1 tie_x0
xfeed_5282 0 1 tie_x0
xfeed_5281 0 1 tie_x0
xfeed_5280 0 1 tie_x0
xfeed_4759 0 1 tie_x0
xfeed_4758 0 1 tie_x0
xfeed_4757 0 1 tie_x0
xfeed_4756 0 1 tie_x0
xfeed_4755 0 1 tie_x0
xfeed_4754 0 1 tie_x0
xfeed_4753 0 1 tie_x0
xfeed_4752 0 1 tie_x0
xfeed_4751 0 1 tie_x0
xfeed_4750 0 1 tie_x0
xsubckt_20_na2_x1 0 1 117 129 119 na2_x1
xfeed_5299 0 1 tie_x0
xfeed_5298 0 1 tie_x0
xfeed_5297 0 1 tie_x0
xfeed_5296 0 1 tie_x0
xfeed_5295 0 1 tie_x0
xfeed_5294 0 1 tie_x0
xfeed_5293 0 1 tie_x0
xfeed_5292 0 1 tie_x0
xfeed_5291 0 1 tie_x0
xfeed_5290 0 1 tie_x0
xfeed_4769 0 1 tie_x0
xfeed_4768 0 1 tie_x0
xfeed_4767 0 1 tie_x0
xfeed_4766 0 1 tie_x0
xfeed_4765 0 1 tie_x0
xfeed_4764 0 1 tie_x0
xfeed_4763 0 1 tie_x0
xfeed_4762 0 1 tie_x0
xfeed_4761 0 1 tie_x0
xfeed_4760 0 1 tie_x0
xfeed_4779 0 1 tie_x0
xfeed_4778 0 1 tie_x0
xfeed_4777 0 1 tie_x0
xfeed_4776 0 1 tie_x0
xfeed_4775 0 1 tie_x0
xfeed_4774 0 1 tie_x0
xfeed_4773 0 1 tie_x0
xfeed_4772 0 1 tie_x0
xfeed_4771 0 1 tie_x0
xfeed_4770 0 1 tie_x0
xfeed_4789 0 1 tie_x0
xfeed_4788 0 1 tie_x0
xfeed_4787 0 1 tie_x0
xfeed_4786 0 1 tie_x0
xfeed_4785 0 1 tie_x0
xfeed_4784 0 1 tie_x0
xfeed_4783 0 1 tie_x0
xfeed_4782 0 1 tie_x0
xfeed_4781 0 1 tie_x0
xfeed_4780 0 1 tie_x0
xsubckt_45_nao22_x1 0 1 93 97 100 102 nao22_x1
xfeed_5409 0 1 tie_x0
xfeed_5408 0 1 tie_x0
xfeed_5407 0 1 tie_x0
xfeed_5406 0 1 tie_x0
xfeed_5405 0 1 tie_x0
xfeed_5404 0 1 tie_x0
xfeed_5403 0 1 tie_x0
xfeed_5402 0 1 tie_x0
xfeed_5401 0 1 tie_x0
xfeed_5400 0 1 tie_x0
xfeed_4799 0 1 tie_x0
xfeed_4798 0 1 tie_x0
xfeed_4797 0 1 tie_x0
xfeed_4796 0 1 tie_x0
xfeed_4795 0 1 tie_x0
xfeed_4794 0 1 tie_x0
xfeed_4793 0 1 tie_x0
xfeed_4792 0 1 tie_x0
xfeed_4791 0 1 tie_x0
xfeed_4790 0 1 tie_x0
xsubckt_5_a2_x2 0 1 130 18 14 a2_x2
xfeed_1100 0 1 tie_x0
xfeed_1101 0 1 tie_x0
xfeed_1102 0 1 tie_x0
xfeed_1103 0 1 tie_x0
xfeed_1104 0 1 tie_x0
xfeed_1105 0 1 tie_x0
xfeed_1106 0 1 tie_x0
xfeed_5419 0 1 tie_x0
xfeed_5418 0 1 tie_x0
xfeed_5417 0 1 tie_x0
xfeed_5416 0 1 tie_x0
xfeed_5415 0 1 tie_x0
xfeed_5414 0 1 tie_x0
xfeed_5413 0 1 tie_x0
xfeed_5412 0 1 tie_x0
xfeed_5411 0 1 tie_x0
xfeed_5410 0 1 tie_x0
xsubckt_24_ao22_x2 0 1 114 122 121 125 ao22_x2
xfeed_1107 0 1 tie_x0
xfeed_1108 0 1 tie_x0
xfeed_1109 0 1 tie_x0
xfeed_1110 0 1 tie_x0
xfeed_1111 0 1 tie_x0
xfeed_1112 0 1 tie_x0
xfeed_1113 0 1 tie_x0
xfeed_5429 0 1 tie_x0
xfeed_5428 0 1 tie_x0
xfeed_5427 0 1 tie_x0
xfeed_5426 0 1 tie_x0
xfeed_5425 0 1 tie_x0
xfeed_5424 0 1 tie_x0
xfeed_5423 0 1 tie_x0
xfeed_5422 0 1 tie_x0
xfeed_5421 0 1 tie_x0
xfeed_5420 0 1 tie_x0
xfeed_1114 0 1 tie_x0
xfeed_1115 0 1 tie_x0
xfeed_1116 0 1 tie_x0
xfeed_1117 0 1 tie_x0
xfeed_1118 0 1 rowend_x0
xfeed_1119 0 1 tie_x0
xfeed_1120 0 1 tie_x0
xfeed_5439 0 1 tie_x0
xfeed_5438 0 1 tie_x0
xfeed_5437 0 1 tie_x0
xfeed_5436 0 1 tie_x0
xfeed_5435 0 1 tie_x0
xfeed_5434 0 1 tie_x0
xfeed_5433 0 1 tie_x0
xfeed_5432 0 1 tie_x0
xfeed_5431 0 1 tie_x0
xfeed_5430 0 1 tie_x0
xfeed_4909 0 1 tie_x0
xfeed_4908 0 1 tie_x0
xfeed_4907 0 1 tie_x0
xfeed_4906 0 1 tie_x0
xfeed_4905 0 1 tie_x0
xfeed_4904 0 1 tie_x0
xfeed_4903 0 1 tie_x0
xfeed_4902 0 1 tie_x0
xfeed_4901 0 1 tie_x0
xfeed_4900 0 1 tie_x0
xsubckt_23_a2_x2 0 1 115 7 2 a2_x2
xfeed_1121 0 1 tie_x0
xfeed_1122 0 1 tie_x0
xfeed_1123 0 1 tie_x0
xfeed_1124 0 1 tie_x0
xfeed_1125 0 1 tie_x0
xfeed_1126 0 1 tie_x0
xfeed_1127 0 1 tie_x0
xfeed_1128 0 1 tie_x0
xfeed_1129 0 1 tie_x0
xfeed_5449 0 1 tie_x0
xfeed_5448 0 1 tie_x0
xfeed_5447 0 1 tie_x0
xfeed_5446 0 1 tie_x0
xfeed_5445 0 1 tie_x0
xfeed_5444 0 1 tie_x0
xfeed_5443 0 1 tie_x0
xfeed_5442 0 1 tie_x0
xfeed_5441 0 1 tie_x0
xfeed_5440 0 1 tie_x0
xfeed_4919 0 1 tie_x0
xfeed_4918 0 1 tie_x0
xfeed_4917 0 1 tie_x0
xfeed_4916 0 1 tie_x0
xfeed_4915 0 1 tie_x0
xfeed_4914 0 1 tie_x0
xfeed_4913 0 1 tie_x0
xfeed_4912 0 1 tie_x0
xfeed_4911 0 1 tie_x0
xfeed_4910 0 1 tie_x0
xsubckt_27_oa2a22_x2 0 1 111 17 12 11 18 oa2a22_x2
xfeed_1130 0 1 tie_x0
xfeed_1131 0 1 tie_x0
xfeed_1132 0 1 tie_x0
xfeed_1133 0 1 tie_x0
xfeed_1134 0 1 tie_x0
xfeed_1135 0 1 tie_x0
xfeed_1136 0 1 tie_x0
xfeed_1137 0 1 tie_x0
xfeed_1138 0 1 tie_x0
xfeed_1139 0 1 tie_x0
xsubckt_113_na2_x1 0 1 165 78 7 na2_x1
xfeed_5459 0 1 tie_x0
xfeed_5458 0 1 tie_x0
xfeed_5457 0 1 tie_x0
xfeed_5456 0 1 tie_x0
xfeed_5455 0 1 tie_x0
xfeed_5454 0 1 tie_x0
xfeed_5453 0 1 tie_x0
xfeed_5452 0 1 tie_x0
xfeed_5451 0 1 tie_x0
xfeed_5450 0 1 tie_x0
xfeed_4929 0 1 tie_x0
xfeed_4928 0 1 tie_x0
xfeed_4927 0 1 tie_x0
xfeed_4926 0 1 tie_x0
xfeed_4925 0 1 tie_x0
xfeed_4924 0 1 tie_x0
xfeed_4923 0 1 tie_x0
xfeed_4922 0 1 tie_x0
xfeed_4921 0 1 tie_x0
xfeed_4920 0 1 tie_x0
xfeed_1140 0 1 tie_x0
xfeed_1141 0 1 tie_x0
xfeed_1142 0 1 tie_x0
xfeed_1143 0 1 tie_x0
xfeed_1144 0 1 tie_x0
xfeed_1145 0 1 tie_x0
xfeed_1146 0 1 tie_x0
xfeed_1147 0 1 tie_x0
xfeed_1148 0 1 tie_x0
xfeed_1149 0 1 tie_x0
xfeed_5469 0 1 tie_x0
xfeed_5468 0 1 tie_x0
xfeed_5467 0 1 tie_x0
xfeed_5466 0 1 tie_x0
xfeed_5465 0 1 tie_x0
xfeed_5464 0 1 tie_x0
xfeed_5463 0 1 tie_x0
xfeed_5462 0 1 tie_x0
xfeed_5461 0 1 tie_x0
xfeed_5460 0 1 tie_x0
xfeed_4939 0 1 tie_x0
xfeed_4938 0 1 tie_x0
xfeed_4937 0 1 tie_x0
xfeed_4936 0 1 tie_x0
xfeed_4935 0 1 tie_x0
xfeed_4934 0 1 tie_x0
xfeed_4933 0 1 tie_x0
xfeed_4932 0 1 rowend_x0
xfeed_4931 0 1 tie_x0
xfeed_4930 0 1 tie_x0
xfeed_1150 0 1 tie_x0
xfeed_1151 0 1 tie_x0
xfeed_1152 0 1 tie_x0
xfeed_1153 0 1 tie_x0
xfeed_1154 0 1 tie_x0
xfeed_1155 0 1 tie_x0
xfeed_1156 0 1 tie_x0
xfeed_1157 0 1 tie_x0
xfeed_1158 0 1 tie_x0
xfeed_1159 0 1 tie_x0
xfeed_5479 0 1 tie_x0
xfeed_5478 0 1 tie_x0
xfeed_5477 0 1 tie_x0
xfeed_5476 0 1 tie_x0
xfeed_5475 0 1 tie_x0
xfeed_5474 0 1 tie_x0
xfeed_5473 0 1 tie_x0
xfeed_5472 0 1 tie_x0
xfeed_5471 0 1 tie_x0
xfeed_5470 0 1 tie_x0
xfeed_4949 0 1 tie_x0
xfeed_4948 0 1 tie_x0
xfeed_4947 0 1 tie_x0
xfeed_4946 0 1 tie_x0
xfeed_4945 0 1 tie_x0
xfeed_4944 0 1 tie_x0
xfeed_4943 0 1 tie_x0
xfeed_4942 0 1 tie_x0
xfeed_4941 0 1 tie_x0
xfeed_4940 0 1 tie_x0
xsubckt_103_a2_x2 0 1 220 131 174 a2_x2
xfeed_1160 0 1 tie_x0
xfeed_1161 0 1 tie_x0
xfeed_1162 0 1 rowend_x0
xfeed_1163 0 1 tie_x0
xfeed_1164 0 1 tie_x0
xfeed_1165 0 1 tie_x0
xfeed_1166 0 1 tie_x0
xfeed_1167 0 1 tie_x0
xfeed_1168 0 1 tie_x0
xfeed_1169 0 1 tie_x0
xsubckt_31_na2_x1 0 1 107 13 16 na2_x1
xfeed_5489 0 1 tie_x0
xfeed_5488 0 1 tie_x0
xfeed_5487 0 1 tie_x0
xfeed_5486 0 1 tie_x0
xfeed_5485 0 1 tie_x0
xfeed_5484 0 1 tie_x0
xfeed_5483 0 1 tie_x0
xfeed_5482 0 1 tie_x0
xfeed_5481 0 1 tie_x0
xfeed_5480 0 1 tie_x0
xfeed_4959 0 1 tie_x0
xfeed_4958 0 1 tie_x0
xfeed_4957 0 1 tie_x0
xfeed_4956 0 1 tie_x0
xfeed_4955 0 1 tie_x0
xfeed_4954 0 1 tie_x0
xfeed_4953 0 1 tie_x0
xfeed_4952 0 1 tie_x0
xfeed_4951 0 1 tie_x0
xfeed_4950 0 1 tie_x0
xfeed_1170 0 1 tie_x0
xfeed_1171 0 1 tie_x0
xfeed_1172 0 1 tie_x0
xfeed_1173 0 1 tie_x0
xfeed_1174 0 1 tie_x0
xfeed_1175 0 1 tie_x0
xfeed_1176 0 1 tie_x0
xfeed_1177 0 1 tie_x0
xfeed_1178 0 1 tie_x0
xfeed_1179 0 1 tie_x0
xsubckt_151_sff1_x4 0 1 7 226 21 sff1_x4
xfeed_6109 0 1 tie_x0
xfeed_6108 0 1 tie_x0
xfeed_6107 0 1 tie_x0
xfeed_6106 0 1 tie_x0
xfeed_6105 0 1 tie_x0
xfeed_6104 0 1 tie_x0
xfeed_6103 0 1 tie_x0
xfeed_6102 0 1 tie_x0
xfeed_6101 0 1 tie_x0
xfeed_6100 0 1 tie_x0
xfeed_5499 0 1 tie_x0
xfeed_5498 0 1 tie_x0
xfeed_5497 0 1 tie_x0
xfeed_5496 0 1 tie_x0
xfeed_5495 0 1 tie_x0
xfeed_5494 0 1 tie_x0
xfeed_5493 0 1 tie_x0
xfeed_5492 0 1 tie_x0
xfeed_5491 0 1 tie_x0
xfeed_5490 0 1 tie_x0
xfeed_4969 0 1 tie_x0
xfeed_4968 0 1 tie_x0
xfeed_4967 0 1 tie_x0
xfeed_4966 0 1 tie_x0
xfeed_4965 0 1 tie_x0
xfeed_4964 0 1 tie_x0
xfeed_4963 0 1 tie_x0
xfeed_4962 0 1 tie_x0
xfeed_4961 0 1 tie_x0
xfeed_4960 0 1 tie_x0
xfeed_1180 0 1 tie_x0
xfeed_1181 0 1 tie_x0
xfeed_1182 0 1 tie_x0
xfeed_1183 0 1 tie_x0
xfeed_1184 0 1 tie_x0
xfeed_1185 0 1 tie_x0
xfeed_1186 0 1 tie_x0
xfeed_1187 0 1 tie_x0
xfeed_1188 0 1 tie_x0
xfeed_1189 0 1 tie_x0
xfeed_6119 0 1 tie_x0
xfeed_6118 0 1 tie_x0
xfeed_6117 0 1 tie_x0
xfeed_6116 0 1 tie_x0
xfeed_6115 0 1 tie_x0
xfeed_6114 0 1 tie_x0
xfeed_6113 0 1 tie_x0
xfeed_6112 0 1 tie_x0
xfeed_6111 0 1 tie_x0
xfeed_6110 0 1 tie_x0
xfeed_4979 0 1 tie_x0
xfeed_4978 0 1 tie_x0
xfeed_4977 0 1 rowend_x0
xfeed_4976 0 1 tie_x0
xfeed_4975 0 1 tie_x0
xfeed_4974 0 1 tie_x0
xfeed_4973 0 1 tie_x0
xfeed_4972 0 1 tie_x0
xfeed_4971 0 1 tie_x0
xfeed_4970 0 1 tie_x0
xfeed_1190 0 1 tie_x0
xfeed_1191 0 1 tie_x0
xfeed_1192 0 1 tie_x0
xfeed_1193 0 1 tie_x0
xfeed_1194 0 1 tie_x0
xfeed_1195 0 1 tie_x0
xfeed_1196 0 1 tie_x0
xfeed_1197 0 1 tie_x0
xfeed_1198 0 1 tie_x0
xfeed_1199 0 1 tie_x0
xfeed_6129 0 1 tie_x0
xfeed_6128 0 1 tie_x0
xfeed_6127 0 1 tie_x0
xfeed_6126 0 1 tie_x0
xfeed_6125 0 1 tie_x0
xfeed_6124 0 1 tie_x0
xfeed_6123 0 1 tie_x0
xfeed_6122 0 1 tie_x0
xfeed_6121 0 1 tie_x0
xfeed_6120 0 1 tie_x0
xfeed_4989 0 1 tie_x0
xfeed_4988 0 1 tie_x0
xfeed_4987 0 1 tie_x0
xfeed_4986 0 1 tie_x0
xfeed_4985 0 1 tie_x0
xfeed_4984 0 1 tie_x0
xfeed_4983 0 1 tie_x0
xfeed_4982 0 1 tie_x0
xfeed_4981 0 1 tie_x0
xfeed_4980 0 1 tie_x0
xfeed_6139 0 1 tie_x0
xfeed_6138 0 1 tie_x0
xfeed_6137 0 1 tie_x0
xfeed_6136 0 1 tie_x0
xfeed_6135 0 1 tie_x0
xfeed_6134 0 1 tie_x0
xfeed_6133 0 1 tie_x0
xfeed_6132 0 1 tie_x0
xfeed_6131 0 1 tie_x0
xfeed_6130 0 1 tie_x0
xfeed_5609 0 1 tie_x0
xfeed_5608 0 1 tie_x0
xfeed_5607 0 1 tie_x0
xfeed_5606 0 1 tie_x0
xfeed_5605 0 1 tie_x0
xfeed_5604 0 1 tie_x0
xfeed_5603 0 1 tie_x0
xfeed_5602 0 1 tie_x0
xfeed_5601 0 1 tie_x0
xfeed_5600 0 1 tie_x0
xfeed_4999 0 1 tie_x0
xfeed_4998 0 1 tie_x0
xfeed_4997 0 1 tie_x0
xfeed_4996 0 1 tie_x0
xfeed_4995 0 1 tie_x0
xfeed_4994 0 1 tie_x0
xfeed_4993 0 1 tie_x0
xfeed_4992 0 1 tie_x0
xfeed_4991 0 1 tie_x0
xfeed_4990 0 1 tie_x0
xfeed_6149 0 1 tie_x0
xfeed_6148 0 1 tie_x0
xfeed_6147 0 1 tie_x0
xfeed_6146 0 1 tie_x0
xfeed_6145 0 1 tie_x0
xfeed_6144 0 1 tie_x0
xfeed_6143 0 1 tie_x0
xfeed_6142 0 1 rowend_x0
xfeed_6141 0 1 tie_x0
xfeed_6140 0 1 tie_x0
xfeed_5619 0 1 tie_x0
xfeed_5618 0 1 tie_x0
xfeed_5617 0 1 tie_x0
xfeed_5616 0 1 tie_x0
xfeed_5615 0 1 tie_x0
xfeed_5614 0 1 tie_x0
xfeed_5613 0 1 tie_x0
xfeed_5612 0 1 tie_x0
xfeed_5611 0 1 tie_x0
xfeed_5610 0 1 tie_x0
xfeed_1300 0 1 tie_x0
xfeed_1301 0 1 tie_x0
xfeed_1302 0 1 tie_x0
xfeed_1303 0 1 tie_x0
xfeed_1304 0 1 tie_x0
xfeed_1305 0 1 tie_x0
xfeed_1306 0 1 tie_x0
xfeed_1307 0 1 tie_x0
xfeed_1308 0 1 tie_x0
xfeed_1309 0 1 tie_x0
xfeed_6159 0 1 tie_x0
xfeed_6158 0 1 tie_x0
xfeed_6157 0 1 tie_x0
xfeed_6156 0 1 tie_x0
xfeed_6155 0 1 tie_x0
xfeed_6154 0 1 tie_x0
xfeed_6153 0 1 tie_x0
xfeed_6152 0 1 tie_x0
xfeed_6151 0 1 tie_x0
xfeed_6150 0 1 tie_x0
xfeed_5629 0 1 tie_x0
xfeed_5628 0 1 tie_x0
xfeed_5627 0 1 tie_x0
xfeed_5626 0 1 tie_x0
xfeed_5625 0 1 tie_x0
xfeed_5624 0 1 tie_x0
xfeed_5623 0 1 tie_x0
xfeed_5622 0 1 tie_x0
xfeed_5621 0 1 tie_x0
xfeed_5620 0 1 tie_x0
xfeed_1310 0 1 tie_x0
xfeed_1311 0 1 tie_x0
xfeed_1312 0 1 tie_x0
xfeed_1313 0 1 tie_x0
xfeed_1314 0 1 tie_x0
xfeed_1315 0 1 tie_x0
xfeed_1316 0 1 tie_x0
xfeed_1317 0 1 tie_x0
xfeed_1318 0 1 rowend_x0
xfeed_1319 0 1 tie_x0
xfeed_6169 0 1 tie_x0
xfeed_6168 0 1 tie_x0
xfeed_6167 0 1 tie_x0
xfeed_6166 0 1 tie_x0
xfeed_6165 0 1 tie_x0
xfeed_6164 0 1 tie_x0
xfeed_6163 0 1 tie_x0
xfeed_6162 0 1 tie_x0
xfeed_6161 0 1 tie_x0
xfeed_6160 0 1 tie_x0
xfeed_5639 0 1 tie_x0
xfeed_5638 0 1 tie_x0
xfeed_5637 0 1 tie_x0
xfeed_5636 0 1 tie_x0
xfeed_5635 0 1 tie_x0
xfeed_5634 0 1 tie_x0
xfeed_5633 0 1 tie_x0
xfeed_5632 0 1 tie_x0
xfeed_5631 0 1 tie_x0
xfeed_5630 0 1 tie_x0
xsubckt_69_nxr2_x1 0 1 202 86 205 nxr2_x1
xfeed_1320 0 1 tie_x0
xfeed_1321 0 1 tie_x0
xfeed_1322 0 1 tie_x0
xfeed_1323 0 1 tie_x0
xfeed_1324 0 1 tie_x0
xfeed_1325 0 1 tie_x0
xfeed_1326 0 1 tie_x0
xfeed_1327 0 1 tie_x0
xfeed_1328 0 1 tie_x0
xfeed_1329 0 1 tie_x0
xfeed_6179 0 1 tie_x0
xfeed_6178 0 1 tie_x0
xfeed_6177 0 1 tie_x0
xfeed_6176 0 1 tie_x0
xfeed_6175 0 1 tie_x0
xfeed_6174 0 1 tie_x0
xfeed_6173 0 1 tie_x0
xfeed_6172 0 1 tie_x0
xfeed_6171 0 1 tie_x0
xfeed_6170 0 1 tie_x0
xfeed_5649 0 1 tie_x0
xfeed_5648 0 1 tie_x0
xfeed_5647 0 1 tie_x0
xfeed_5646 0 1 tie_x0
xfeed_5645 0 1 tie_x0
xfeed_5644 0 1 tie_x0
xfeed_5643 0 1 tie_x0
xfeed_5642 0 1 tie_x0
xfeed_5641 0 1 tie_x0
xfeed_5640 0 1 tie_x0
xsubckt_128_na2_x1 0 1 152 76 5 na2_x1
xfeed_1330 0 1 tie_x0
xfeed_1331 0 1 tie_x0
xfeed_1332 0 1 tie_x0
xfeed_1333 0 1 tie_x0
xfeed_1334 0 1 tie_x0
xfeed_1335 0 1 tie_x0
xfeed_1336 0 1 tie_x0
xfeed_1337 0 1 tie_x0
xfeed_1338 0 1 tie_x0
xfeed_1339 0 1 tie_x0
xfeed_6189 0 1 tie_x0
xfeed_6188 0 1 tie_x0
xfeed_6187 0 1 tie_x0
xfeed_6186 0 1 tie_x0
xfeed_6185 0 1 tie_x0
xfeed_6184 0 1 tie_x0
xfeed_6183 0 1 tie_x0
xfeed_6182 0 1 tie_x0
xfeed_6181 0 1 tie_x0
xfeed_6180 0 1 tie_x0
xfeed_5659 0 1 tie_x0
xfeed_5658 0 1 tie_x0
xfeed_5657 0 1 tie_x0
xfeed_5656 0 1 tie_x0
xfeed_5655 0 1 tie_x0
xfeed_5654 0 1 tie_x0
xfeed_5653 0 1 tie_x0
xfeed_5652 0 1 tie_x0
xfeed_5651 0 1 tie_x0
xfeed_5650 0 1 tie_x0
xfeed_1340 0 1 tie_x0
xfeed_1341 0 1 tie_x0
xfeed_1342 0 1 tie_x0
xfeed_1343 0 1 tie_x0
xfeed_1344 0 1 tie_x0
xfeed_1345 0 1 tie_x0
xfeed_1346 0 1 tie_x0
xfeed_1347 0 1 tie_x0
xfeed_1348 0 1 tie_x0
xfeed_1349 0 1 tie_x0
xfeed_6199 0 1 tie_x0
xfeed_6198 0 1 tie_x0
xfeed_6197 0 1 tie_x0
xfeed_6196 0 1 tie_x0
xfeed_6195 0 1 tie_x0
xfeed_6194 0 1 tie_x0
xfeed_6193 0 1 tie_x0
xfeed_6192 0 1 tie_x0
xfeed_6191 0 1 tie_x0
xfeed_6190 0 1 tie_x0
xfeed_5669 0 1 tie_x0
xfeed_5668 0 1 tie_x0
xfeed_5667 0 1 tie_x0
xfeed_5666 0 1 tie_x0
xfeed_5665 0 1 tie_x0
xfeed_5664 0 1 tie_x0
xfeed_5663 0 1 tie_x0
xfeed_5662 0 1 tie_x0
xfeed_5661 0 1 tie_x0
xfeed_5660 0 1 tie_x0
xfeed_1350 0 1 tie_x0
xfeed_1351 0 1 tie_x0
xfeed_1352 0 1 tie_x0
xfeed_1353 0 1 tie_x0
xfeed_1354 0 1 tie_x0
xfeed_1355 0 1 tie_x0
xfeed_1356 0 1 tie_x0
xfeed_1357 0 1 tie_x0
xfeed_1358 0 1 tie_x0
xfeed_1359 0 1 tie_x0
xfeed_5679 0 1 tie_x0
xfeed_5678 0 1 tie_x0
xfeed_5677 0 1 tie_x0
xfeed_5676 0 1 tie_x0
xfeed_5675 0 1 tie_x0
xfeed_5674 0 1 tie_x0
xfeed_5673 0 1 tie_x0
xfeed_5672 0 1 tie_x0
xfeed_5671 0 1 tie_x0
xfeed_5670 0 1 tie_x0
xfeed_1360 0 1 tie_x0
xfeed_1361 0 1 tie_x0
xfeed_1362 0 1 tie_x0
xfeed_1363 0 1 tie_x0
xfeed_1364 0 1 tie_x0
xfeed_1365 0 1 tie_x0
xfeed_1366 0 1 tie_x0
xfeed_1367 0 1 tie_x0
xfeed_1368 0 1 tie_x0
xfeed_1369 0 1 tie_x0
xfeed_5689 0 1 tie_x0
xfeed_5688 0 1 tie_x0
xfeed_5687 0 1 tie_x0
xfeed_5686 0 1 tie_x0
xfeed_5685 0 1 tie_x0
xfeed_5684 0 1 tie_x0
xfeed_5683 0 1 tie_x0
xfeed_5682 0 1 tie_x0
xfeed_5681 0 1 tie_x0
xfeed_5680 0 1 tie_x0
xfeed_1370 0 1 tie_x0
xfeed_1371 0 1 tie_x0
xfeed_1372 0 1 tie_x0
xfeed_1373 0 1 tie_x0
xfeed_1374 0 1 tie_x0
xfeed_1375 0 1 tie_x0
xfeed_1376 0 1 tie_x0
xfeed_1377 0 1 tie_x0
xfeed_1378 0 1 tie_x0
xfeed_1379 0 1 tie_x0
xfeed_6309 0 1 tie_x0
xfeed_6308 0 1 tie_x0
xfeed_6307 0 1 tie_x0
xfeed_6306 0 1 tie_x0
xfeed_6305 0 1 tie_x0
xfeed_6304 0 1 tie_x0
xfeed_6303 0 1 tie_x0
xfeed_6302 0 1 tie_x0
xfeed_6301 0 1 tie_x0
xfeed_6300 0 1 rowend_x0
xfeed_5699 0 1 tie_x0
xfeed_5698 0 1 tie_x0
xfeed_5697 0 1 tie_x0
xfeed_5696 0 1 tie_x0
xfeed_5695 0 1 tie_x0
xfeed_5694 0 1 tie_x0
xfeed_5693 0 1 tie_x0
xfeed_5692 0 1 tie_x0
xfeed_5691 0 1 tie_x0
xfeed_5690 0 1 tie_x0
xfeed_1380 0 1 tie_x0
xfeed_1381 0 1 tie_x0
xfeed_1382 0 1 tie_x0
xfeed_1383 0 1 tie_x0
xfeed_1384 0 1 tie_x0
xfeed_1385 0 1 tie_x0
xfeed_1386 0 1 tie_x0
xfeed_1387 0 1 tie_x0
xfeed_1388 0 1 tie_x0
xfeed_1389 0 1 tie_x0
xfeed_6319 0 1 tie_x0
xfeed_6318 0 1 tie_x0
xfeed_6317 0 1 tie_x0
xfeed_6316 0 1 tie_x0
xfeed_6315 0 1 tie_x0
xfeed_6314 0 1 tie_x0
xfeed_6313 0 1 tie_x0
xfeed_6312 0 1 tie_x0
xfeed_6311 0 1 tie_x0
xfeed_6310 0 1 tie_x0
xfeed_1390 0 1 rowend_x0
xfeed_1391 0 1 tie_x0
xfeed_1392 0 1 tie_x0
xfeed_1393 0 1 tie_x0
xfeed_1394 0 1 tie_x0
xfeed_1395 0 1 tie_x0
xfeed_1396 0 1 tie_x0
xfeed_1397 0 1 tie_x0
xfeed_1398 0 1 tie_x0
xfeed_1399 0 1 tie_x0
xfeed_2000 0 1 tie_x0
xfeed_2001 0 1 tie_x0
xfeed_2002 0 1 tie_x0
xfeed_2003 0 1 rowend_x0
xfeed_2004 0 1 tie_x0
xfeed_2005 0 1 tie_x0
xfeed_2006 0 1 tie_x0
xfeed_2007 0 1 tie_x0
xfeed_2008 0 1 tie_x0
xfeed_2009 0 1 tie_x0
xfeed_6329 0 1 tie_x0
xfeed_6328 0 1 tie_x0
xfeed_6327 0 1 tie_x0
xfeed_6326 0 1 tie_x0
xfeed_6325 0 1 rowend_x0
xfeed_6324 0 1 tie_x0
xfeed_6323 0 1 tie_x0
xfeed_6322 0 1 tie_x0
xfeed_6321 0 1 tie_x0
xfeed_6320 0 1 tie_x0
xfeed_2010 0 1 tie_x0
xfeed_2011 0 1 tie_x0
xfeed_2012 0 1 tie_x0
xfeed_2013 0 1 tie_x0
xfeed_2014 0 1 tie_x0
xfeed_2015 0 1 tie_x0
xfeed_2016 0 1 tie_x0
xfeed_2017 0 1 tie_x0
xfeed_2018 0 1 tie_x0
xfeed_2019 0 1 tie_x0
xfeed_6339 0 1 tie_x0
xfeed_6338 0 1 tie_x0
xfeed_6337 0 1 tie_x0
xfeed_6336 0 1 tie_x0
xfeed_6335 0 1 tie_x0
xfeed_6334 0 1 tie_x0
xfeed_6333 0 1 tie_x0
xfeed_6332 0 1 tie_x0
xfeed_6331 0 1 tie_x0
xfeed_6330 0 1 tie_x0
xfeed_5809 0 1 tie_x0
xfeed_5808 0 1 tie_x0
xfeed_5807 0 1 tie_x0
xfeed_5806 0 1 tie_x0
xfeed_5805 0 1 tie_x0
xfeed_5804 0 1 tie_x0
xfeed_5803 0 1 tie_x0
xfeed_5802 0 1 tie_x0
xfeed_5801 0 1 tie_x0
xfeed_5800 0 1 tie_x0
xfeed_2020 0 1 tie_x0
xfeed_2021 0 1 tie_x0
xfeed_2022 0 1 tie_x0
xfeed_2023 0 1 tie_x0
xfeed_2024 0 1 tie_x0
xfeed_2025 0 1 tie_x0
xfeed_2026 0 1 tie_x0
xfeed_2027 0 1 tie_x0
xfeed_2028 0 1 tie_x0
xfeed_2029 0 1 tie_x0
xfeed_6349 0 1 tie_x0
xfeed_6348 0 1 tie_x0
xfeed_6347 0 1 tie_x0
xfeed_6346 0 1 tie_x0
xfeed_6345 0 1 tie_x0
xfeed_6344 0 1 tie_x0
xfeed_6343 0 1 tie_x0
xfeed_6342 0 1 tie_x0
xfeed_6341 0 1 tie_x0
xfeed_6340 0 1 tie_x0
xfeed_5819 0 1 tie_x0
xfeed_5818 0 1 tie_x0
xfeed_5817 0 1 tie_x0
xfeed_5816 0 1 tie_x0
xfeed_5815 0 1 tie_x0
xfeed_5814 0 1 tie_x0
xfeed_5813 0 1 tie_x0
xfeed_5812 0 1 tie_x0
xfeed_5811 0 1 tie_x0
xfeed_5810 0 1 tie_x0
xfeed_1500 0 1 tie_x0
xfeed_1501 0 1 tie_x0
xfeed_1502 0 1 tie_x0
xfeed_1503 0 1 tie_x0
xfeed_1504 0 1 tie_x0
xfeed_1505 0 1 tie_x0
xfeed_1506 0 1 tie_x0
xfeed_1507 0 1 tie_x0
xfeed_1508 0 1 tie_x0
xfeed_1509 0 1 tie_x0
xfeed_2030 0 1 tie_x0
xfeed_2031 0 1 tie_x0
xfeed_2032 0 1 tie_x0
xfeed_2033 0 1 tie_x0
xfeed_2034 0 1 tie_x0
xfeed_2035 0 1 tie_x0
xfeed_2036 0 1 tie_x0
xfeed_2037 0 1 tie_x0
xfeed_2038 0 1 tie_x0
xfeed_2039 0 1 tie_x0
xfeed_6359 0 1 tie_x0
xfeed_6358 0 1 tie_x0
xfeed_6357 0 1 tie_x0
xfeed_6356 0 1 tie_x0
xfeed_6355 0 1 tie_x0
xfeed_6354 0 1 tie_x0
xfeed_6353 0 1 tie_x0
xfeed_6352 0 1 tie_x0
xfeed_6351 0 1 tie_x0
xfeed_6350 0 1 tie_x0
xfeed_5829 0 1 tie_x0
xfeed_5828 0 1 tie_x0
xfeed_5827 0 1 tie_x0
xfeed_5826 0 1 tie_x0
xfeed_5825 0 1 tie_x0
xfeed_5824 0 1 tie_x0
xfeed_5823 0 1 tie_x0
xfeed_5822 0 1 tie_x0
xfeed_5821 0 1 tie_x0
xfeed_5820 0 1 tie_x0
xsubckt_124_nxr2_x1 0 1 155 160 157 nxr2_x1
xfeed_1510 0 1 tie_x0
xfeed_1511 0 1 tie_x0
xfeed_1512 0 1 tie_x0
xfeed_1513 0 1 tie_x0
xfeed_1514 0 1 tie_x0
xfeed_1515 0 1 tie_x0
xfeed_1516 0 1 tie_x0
xfeed_1517 0 1 tie_x0
xfeed_1518 0 1 tie_x0
xfeed_1519 0 1 tie_x0
xfeed_2040 0 1 tie_x0
xfeed_2041 0 1 tie_x0
xfeed_2042 0 1 tie_x0
xfeed_2043 0 1 tie_x0
xfeed_2044 0 1 tie_x0
xfeed_2045 0 1 tie_x0
xfeed_2046 0 1 tie_x0
xfeed_2047 0 1 tie_x0
xfeed_2048 0 1 tie_x0
xfeed_2049 0 1 tie_x0
xfeed_6369 0 1 tie_x0
xfeed_6368 0 1 tie_x0
xfeed_6367 0 1 tie_x0
xfeed_6366 0 1 tie_x0
xfeed_6365 0 1 tie_x0
xfeed_6364 0 1 tie_x0
xfeed_6363 0 1 tie_x0
xfeed_6362 0 1 tie_x0
xfeed_6361 0 1 tie_x0
xfeed_6360 0 1 tie_x0
xfeed_5839 0 1 tie_x0
xfeed_5838 0 1 tie_x0
xfeed_5837 0 1 tie_x0
xfeed_5836 0 1 tie_x0
xfeed_5835 0 1 tie_x0
xfeed_5834 0 1 tie_x0
xfeed_5833 0 1 tie_x0
xfeed_5832 0 1 tie_x0
xfeed_5831 0 1 tie_x0
xfeed_5830 0 1 tie_x0
xfeed_1520 0 1 tie_x0
xfeed_1521 0 1 tie_x0
xfeed_1522 0 1 tie_x0
xfeed_1523 0 1 tie_x0
xfeed_1524 0 1 tie_x0
xfeed_1525 0 1 tie_x0
xfeed_1526 0 1 tie_x0
xfeed_1527 0 1 tie_x0
xfeed_1528 0 1 tie_x0
xfeed_1529 0 1 tie_x0
xfeed_2050 0 1 tie_x0
xfeed_2051 0 1 tie_x0
xfeed_2052 0 1 tie_x0
xfeed_2053 0 1 tie_x0
xfeed_2054 0 1 rowend_x0
xfeed_2055 0 1 tie_x0
xfeed_2056 0 1 tie_x0
xfeed_2057 0 1 tie_x0
xfeed_2058 0 1 tie_x0
xfeed_2059 0 1 tie_x0
xfeed_6379 0 1 tie_x0
xfeed_6378 0 1 tie_x0
xfeed_6377 0 1 tie_x0
xfeed_6376 0 1 tie_x0
xfeed_6375 0 1 tie_x0
xfeed_6374 0 1 tie_x0
xfeed_6373 0 1 tie_x0
xfeed_6372 0 1 tie_x0
xfeed_6371 0 1 tie_x0
xfeed_6370 0 1 tie_x0
xfeed_5849 0 1 tie_x0
xfeed_5848 0 1 tie_x0
xfeed_5847 0 1 tie_x0
xfeed_5846 0 1 tie_x0
xfeed_5845 0 1 tie_x0
xfeed_5844 0 1 tie_x0
xfeed_5843 0 1 tie_x0
xfeed_5842 0 1 tie_x0
xfeed_5841 0 1 tie_x0
xfeed_5840 0 1 tie_x0
xfeed_1530 0 1 tie_x0
xfeed_1531 0 1 tie_x0
xfeed_1532 0 1 tie_x0
xfeed_1533 0 1 tie_x0
xfeed_1534 0 1 tie_x0
xfeed_1535 0 1 tie_x0
xfeed_1536 0 1 tie_x0
xfeed_1537 0 1 tie_x0
xfeed_1538 0 1 tie_x0
xfeed_1539 0 1 tie_x0
xfeed_2060 0 1 tie_x0
xfeed_2061 0 1 tie_x0
xfeed_2062 0 1 tie_x0
xfeed_2063 0 1 tie_x0
xfeed_2064 0 1 tie_x0
xfeed_2065 0 1 tie_x0
xfeed_2066 0 1 tie_x0
xfeed_2067 0 1 tie_x0
xfeed_2068 0 1 tie_x0
xfeed_2069 0 1 tie_x0
xsubckt_11_mx2_x2 0 1 228 9 126 2 mx2_x2
xfeed_6389 0 1 tie_x0
xfeed_6388 0 1 tie_x0
xfeed_6387 0 1 tie_x0
xfeed_6386 0 1 tie_x0
xfeed_6385 0 1 tie_x0
xfeed_6384 0 1 tie_x0
xfeed_6383 0 1 tie_x0
xfeed_6382 0 1 tie_x0
xfeed_6381 0 1 tie_x0
xfeed_6380 0 1 tie_x0
xfeed_5859 0 1 tie_x0
xfeed_5858 0 1 tie_x0
xfeed_5857 0 1 tie_x0
xfeed_5856 0 1 tie_x0
xfeed_5855 0 1 tie_x0
xfeed_5854 0 1 tie_x0
xfeed_5853 0 1 tie_x0
xfeed_5852 0 1 tie_x0
xfeed_5851 0 1 tie_x0
xfeed_5850 0 1 tie_x0
xsubckt_85_ao22_x2 0 1 188 192 190 204 ao22_x2
xfeed_1540 0 1 tie_x0
xfeed_1541 0 1 tie_x0
xfeed_1542 0 1 tie_x0
xfeed_1543 0 1 tie_x0
xfeed_1544 0 1 tie_x0
xfeed_1545 0 1 tie_x0
xfeed_1546 0 1 tie_x0
xfeed_1547 0 1 tie_x0
xfeed_1548 0 1 rowend_x0
xfeed_1549 0 1 tie_x0
xfeed_2070 0 1 tie_x0
xfeed_2071 0 1 tie_x0
xfeed_2072 0 1 tie_x0
xfeed_2073 0 1 tie_x0
xfeed_2074 0 1 tie_x0
xfeed_2075 0 1 tie_x0
xfeed_2076 0 1 tie_x0
xfeed_2077 0 1 tie_x0
xfeed_2078 0 1 tie_x0
xfeed_2079 0 1 tie_x0
xfeed_7009 0 1 tie_x0
xfeed_7008 0 1 tie_x0
xfeed_7007 0 1 tie_x0
xfeed_7006 0 1 tie_x0
xfeed_7005 0 1 tie_x0
xfeed_7004 0 1 tie_x0
xfeed_7003 0 1 tie_x0
xfeed_7002 0 1 tie_x0
xfeed_7001 0 1 tie_x0
xfeed_7000 0 1 tie_x0
xfeed_6399 0 1 tie_x0
xfeed_6398 0 1 tie_x0
xfeed_6397 0 1 tie_x0
xfeed_6396 0 1 tie_x0
xfeed_6395 0 1 tie_x0
xfeed_6394 0 1 tie_x0
xfeed_6393 0 1 tie_x0
xfeed_6392 0 1 tie_x0
xfeed_6391 0 1 tie_x0
xfeed_6390 0 1 tie_x0
xfeed_5869 0 1 tie_x0
xfeed_5868 0 1 tie_x0
xfeed_5867 0 1 tie_x0
xfeed_5866 0 1 tie_x0
xfeed_5865 0 1 tie_x0
xfeed_5864 0 1 tie_x0
xfeed_5863 0 1 tie_x0
xfeed_5862 0 1 tie_x0
xfeed_5861 0 1 tie_x0
xfeed_5860 0 1 tie_x0
xsubckt_51_na2_x1 0 1 88 6 2 na2_x1
xfeed_1550 0 1 tie_x0
xfeed_1551 0 1 tie_x0
xfeed_1552 0 1 tie_x0
xfeed_1553 0 1 tie_x0
xfeed_1554 0 1 tie_x0
xfeed_1555 0 1 tie_x0
xfeed_1556 0 1 tie_x0
xfeed_1557 0 1 tie_x0
xfeed_1558 0 1 tie_x0
xfeed_1559 0 1 tie_x0
xfeed_2080 0 1 tie_x0
xfeed_2081 0 1 tie_x0
xfeed_2082 0 1 tie_x0
xfeed_2083 0 1 tie_x0
xfeed_2084 0 1 tie_x0
xfeed_2085 0 1 tie_x0
xfeed_2086 0 1 tie_x0
xfeed_2087 0 1 tie_x0
xfeed_2088 0 1 tie_x0
xfeed_2089 0 1 tie_x0
xfeed_7019 0 1 tie_x0
xfeed_7018 0 1 tie_x0
xfeed_7017 0 1 tie_x0
xfeed_7016 0 1 tie_x0
xfeed_7015 0 1 tie_x0
xfeed_7014 0 1 tie_x0
xfeed_7013 0 1 tie_x0
xfeed_7012 0 1 tie_x0
xfeed_7011 0 1 tie_x0
xfeed_7010 0 1 tie_x0
xfeed_5876 0 1 tie_x0
xfeed_5875 0 1 tie_x0
xfeed_5874 0 1 tie_x0
xfeed_5873 0 1 tie_x0
xfeed_5872 0 1 tie_x0
xfeed_5871 0 1 tie_x0
xfeed_5870 0 1 tie_x0
xsubckt_153_sff1_x4 0 1 5 224 66 sff1_x4
xspare_feed_100 0 1 rowend_x0
xspare_feed_101 0 1 tie_x0
xspare_feed_102 0 1 rowend_x0
xspare_feed_103 0 1 rowend_x0
xspare_feed_104 0 1 tie_x0
xspare_feed_105 0 1 rowend_x0
xspare_feed_106 0 1 tie_x0
xspare_feed_107 0 1 rowend_x0
xspare_feed_108 0 1 rowend_x0
xspare_feed_109 0 1 tie_x0
xfeed_1560 0 1 tie_x0
xfeed_1561 0 1 tie_x0
xfeed_1562 0 1 tie_x0
xfeed_1563 0 1 tie_x0
xfeed_1564 0 1 tie_x0
xfeed_1565 0 1 tie_x0
xfeed_1566 0 1 tie_x0
xfeed_1567 0 1 tie_x0
xfeed_1568 0 1 tie_x0
xfeed_1569 0 1 tie_x0
xfeed_2090 0 1 tie_x0
xfeed_2091 0 1 tie_x0
xfeed_2092 0 1 tie_x0
xfeed_2093 0 1 tie_x0
xfeed_2094 0 1 tie_x0
xfeed_2095 0 1 tie_x0
xfeed_2096 0 1 tie_x0
xfeed_2097 0 1 tie_x0
xfeed_2098 0 1 tie_x0
xfeed_2099 0 1 tie_x0
xfeed_5879 0 1 tie_x0
xfeed_5878 0 1 tie_x0
xfeed_5877 0 1 tie_x0
xsubckt_149_sff1_x4 0 1 9 228 24 sff1_x4
xfeed_7029 0 1 tie_x0
xfeed_7028 0 1 tie_x0
xfeed_7027 0 1 tie_x0
xfeed_7026 0 1 tie_x0
xfeed_7025 0 1 tie_x0
xfeed_7024 0 1 tie_x0
xfeed_7023 0 1 tie_x0
xfeed_7022 0 1 tie_x0
xfeed_7021 0 1 tie_x0
xfeed_7020 0 1 tie_x0
xfeed_5883 0 1 tie_x0
xfeed_5882 0 1 tie_x0
xfeed_5881 0 1 tie_x0
xfeed_5880 0 1 tie_x0
xspare_feed_110 0 1 rowend_x0
xspare_feed_111 0 1 tie_x0
xspare_feed_112 0 1 rowend_x0
xspare_feed_113 0 1 rowend_x0
xspare_feed_114 0 1 tie_x0
xspare_feed_115 0 1 rowend_x0
xspare_feed_116 0 1 tie_x0
xspare_feed_117 0 1 rowend_x0
xspare_feed_118 0 1 rowend_x0
xspare_feed_119 0 1 tie_x0
xfeed_1570 0 1 tie_x0
xfeed_1571 0 1 tie_x0
xfeed_1572 0 1 tie_x0
xfeed_1573 0 1 tie_x0
xfeed_1574 0 1 tie_x0
xfeed_1575 0 1 tie_x0
xfeed_1576 0 1 tie_x0
xfeed_1577 0 1 tie_x0
xfeed_1578 0 1 tie_x0
xfeed_1579 0 1 tie_x0
xfeed_5889 0 1 tie_x0
xfeed_5888 0 1 tie_x0
xfeed_5887 0 1 tie_x0
xfeed_5886 0 1 tie_x0
xfeed_5885 0 1 tie_x0
xfeed_5884 0 1 tie_x0
xfeed_7039 0 1 tie_x0
xfeed_7038 0 1 tie_x0
xfeed_7037 0 1 tie_x0
xfeed_7036 0 1 tie_x0
xfeed_7035 0 1 tie_x0
xfeed_7034 0 1 tie_x0
xfeed_7033 0 1 tie_x0
xfeed_7032 0 1 tie_x0
xfeed_7031 0 1 tie_x0
xfeed_7030 0 1 tie_x0
xfeed_6509 0 1 tie_x0
xfeed_6508 0 1 tie_x0
xfeed_6507 0 1 tie_x0
xfeed_6506 0 1 tie_x0
xfeed_6505 0 1 tie_x0
xfeed_6504 0 1 tie_x0
xfeed_6503 0 1 tie_x0
xfeed_6502 0 1 tie_x0
xfeed_6501 0 1 tie_x0
xfeed_6500 0 1 tie_x0
xfeed_5890 0 1 tie_x0
xspare_feed_120 0 1 rowend_x0
xspare_feed_121 0 1 tie_x0
xspare_feed_122 0 1 rowend_x0
xspare_feed_123 0 1 rowend_x0
xspare_feed_124 0 1 tie_x0
xspare_feed_125 0 1 rowend_x0
xspare_feed_126 0 1 tie_x0
xspare_feed_127 0 1 rowend_x0
xspare_feed_128 0 1 rowend_x0
xspare_feed_129 0 1 tie_x0
xfeed_1580 0 1 tie_x0
xfeed_1581 0 1 tie_x0
xfeed_1582 0 1 tie_x0
xfeed_1583 0 1 tie_x0
xfeed_1584 0 1 tie_x0
xfeed_1585 0 1 tie_x0
xfeed_1586 0 1 tie_x0
xfeed_1587 0 1 tie_x0
xfeed_1588 0 1 tie_x0
xfeed_1589 0 1 tie_x0
xfeed_5899 0 1 tie_x0
xfeed_5898 0 1 tie_x0
xfeed_5897 0 1 tie_x0
xfeed_5896 0 1 tie_x0
xfeed_5895 0 1 tie_x0
xfeed_5894 0 1 tie_x0
xfeed_5893 0 1 tie_x0
xfeed_5892 0 1 tie_x0
xfeed_5891 0 1 rowend_x0
xfeed_7049 0 1 tie_x0
xfeed_7048 0 1 tie_x0
xfeed_7047 0 1 tie_x0
xfeed_7046 0 1 tie_x0
xfeed_7045 0 1 tie_x0
xfeed_7044 0 1 tie_x0
xfeed_7043 0 1 tie_x0
xfeed_7042 0 1 tie_x0
xfeed_7041 0 1 tie_x0
xfeed_7040 0 1 tie_x0
xfeed_6519 0 1 tie_x0
xfeed_6518 0 1 tie_x0
xfeed_6517 0 1 tie_x0
xfeed_6516 0 1 tie_x0
xfeed_6515 0 1 tie_x0
xfeed_6514 0 1 tie_x0
xfeed_6513 0 1 tie_x0
xfeed_6512 0 1 tie_x0
xfeed_6511 0 1 tie_x0
xfeed_6510 0 1 tie_x0
xfeed_2209 0 1 tie_x0
xfeed_2208 0 1 tie_x0
xfeed_2207 0 1 tie_x0
xfeed_2206 0 1 tie_x0
xfeed_2205 0 1 tie_x0
xfeed_2204 0 1 tie_x0
xfeed_2203 0 1 tie_x0
xfeed_2202 0 1 tie_x0
xfeed_2201 0 1 tie_x0
xfeed_2200 0 1 rowend_x0
xspare_feed_130 0 1 rowend_x0
xspare_feed_131 0 1 tie_x0
xspare_feed_132 0 1 rowend_x0
xspare_feed_133 0 1 rowend_x0
xspare_feed_134 0 1 tie_x0
xspare_feed_135 0 1 rowend_x0
xspare_feed_136 0 1 tie_x0
xspare_feed_137 0 1 rowend_x0
xspare_feed_138 0 1 rowend_x0
xspare_feed_139 0 1 tie_x0
xfeed_1590 0 1 tie_x0
xfeed_1591 0 1 tie_x0
xfeed_1592 0 1 tie_x0
xfeed_1593 0 1 tie_x0
xfeed_1594 0 1 tie_x0
xfeed_1595 0 1 tie_x0
xfeed_1596 0 1 rowend_x0
xfeed_1597 0 1 tie_x0
xfeed_1598 0 1 tie_x0
xfeed_1599 0 1 tie_x0
xfeed_7059 0 1 tie_x0
xfeed_7058 0 1 tie_x0
xfeed_7057 0 1 tie_x0
xfeed_7056 0 1 tie_x0
xfeed_7055 0 1 tie_x0
xfeed_7054 0 1 tie_x0
xfeed_7053 0 1 tie_x0
xfeed_7052 0 1 tie_x0
xfeed_7051 0 1 tie_x0
xfeed_7050 0 1 tie_x0
xfeed_6529 0 1 tie_x0
xfeed_6528 0 1 tie_x0
xfeed_6527 0 1 tie_x0
xfeed_6526 0 1 tie_x0
xfeed_6525 0 1 tie_x0
xfeed_6524 0 1 tie_x0
xfeed_6523 0 1 tie_x0
xfeed_6522 0 1 tie_x0
xfeed_6521 0 1 tie_x0
xfeed_6520 0 1 tie_x0
xfeed_2219 0 1 tie_x0
xfeed_2218 0 1 tie_x0
xfeed_2217 0 1 tie_x0
xfeed_2216 0 1 tie_x0
xfeed_2215 0 1 tie_x0
xfeed_2214 0 1 tie_x0
xfeed_2213 0 1 tie_x0
xfeed_2212 0 1 tie_x0
xfeed_2211 0 1 tie_x0
xfeed_2210 0 1 tie_x0
xspare_feed_140 0 1 rowend_x0
xspare_feed_141 0 1 tie_x0
xspare_feed_142 0 1 rowend_x0
xspare_feed_143 0 1 rowend_x0
xspare_feed_144 0 1 tie_x0
xspare_feed_145 0 1 rowend_x0
xspare_feed_146 0 1 tie_x0
xspare_feed_147 0 1 rowend_x0
xspare_feed_148 0 1 rowend_x0
xspare_feed_149 0 1 tie_x0
xfeed_7069 0 1 tie_x0
xfeed_7068 0 1 tie_x0
xfeed_7067 0 1 tie_x0
xfeed_7066 0 1 tie_x0
xfeed_7065 0 1 tie_x0
xfeed_7064 0 1 tie_x0
xfeed_7063 0 1 tie_x0
xfeed_7062 0 1 tie_x0
xfeed_7061 0 1 tie_x0
xfeed_7060 0 1 tie_x0
xfeed_6539 0 1 tie_x0
xfeed_6538 0 1 tie_x0
xfeed_6537 0 1 tie_x0
xfeed_6536 0 1 tie_x0
xfeed_6535 0 1 tie_x0
xfeed_6534 0 1 tie_x0
xfeed_6533 0 1 tie_x0
xfeed_6532 0 1 tie_x0
xfeed_6531 0 1 tie_x0
xfeed_6530 0 1 tie_x0
xfeed_2229 0 1 tie_x0
xfeed_2228 0 1 tie_x0
xfeed_2227 0 1 tie_x0
xfeed_2226 0 1 tie_x0
xfeed_2225 0 1 tie_x0
xfeed_2224 0 1 tie_x0
xfeed_2223 0 1 tie_x0
xfeed_2222 0 1 tie_x0
xfeed_2221 0 1 tie_x0
xfeed_2220 0 1 tie_x0
xspare_feed_150 0 1 rowend_x0
xspare_feed_151 0 1 tie_x0
xspare_feed_152 0 1 rowend_x0
xspare_feed_153 0 1 rowend_x0
xspare_feed_154 0 1 tie_x0
xspare_feed_155 0 1 rowend_x0
xspare_feed_156 0 1 tie_x0
xspare_feed_157 0 1 rowend_x0
xspare_feed_158 0 1 rowend_x0
xspare_feed_159 0 1 tie_x0
xfeed_209 0 1 tie_x0
xfeed_208 0 1 tie_x0
xfeed_207 0 1 tie_x0
xfeed_206 0 1 tie_x0
xfeed_205 0 1 tie_x0
xfeed_204 0 1 tie_x0
xfeed_203 0 1 tie_x0
xfeed_202 0 1 tie_x0
xfeed_201 0 1 tie_x0
xfeed_200 0 1 tie_x0
xfeed_7079 0 1 tie_x0
xfeed_7078 0 1 tie_x0
xfeed_7077 0 1 tie_x0
xfeed_7076 0 1 tie_x0
xfeed_7075 0 1 tie_x0
xfeed_7074 0 1 tie_x0
xfeed_7073 0 1 tie_x0
xfeed_7072 0 1 tie_x0
xfeed_7071 0 1 tie_x0
xfeed_7070 0 1 tie_x0
xfeed_6549 0 1 tie_x0
xfeed_6548 0 1 tie_x0
xfeed_6547 0 1 tie_x0
xfeed_6546 0 1 tie_x0
xfeed_6545 0 1 tie_x0
xfeed_6544 0 1 rowend_x0
xfeed_6543 0 1 tie_x0
xfeed_6542 0 1 tie_x0
xfeed_6541 0 1 tie_x0
xfeed_6540 0 1 tie_x0
xfeed_2239 0 1 tie_x0
xfeed_2238 0 1 tie_x0
xfeed_2237 0 1 tie_x0
xfeed_2236 0 1 tie_x0
xfeed_2235 0 1 tie_x0
xfeed_2234 0 1 tie_x0
xfeed_2233 0 1 tie_x0
xfeed_2232 0 1 tie_x0
xfeed_2231 0 1 tie_x0
xfeed_2230 0 1 tie_x0
xspare_feed_160 0 1 rowend_x0
xspare_feed_161 0 1 tie_x0
xspare_feed_162 0 1 rowend_x0
xspare_feed_163 0 1 rowend_x0
xspare_feed_164 0 1 tie_x0
xspare_feed_165 0 1 rowend_x0
xspare_feed_166 0 1 tie_x0
xspare_feed_167 0 1 rowend_x0
xspare_feed_168 0 1 rowend_x0
xspare_feed_169 0 1 tie_x0
xfeed_1700 0 1 tie_x0
xfeed_1701 0 1 tie_x0
xfeed_1702 0 1 tie_x0
xfeed_1703 0 1 tie_x0
xfeed_1704 0 1 tie_x0
xfeed_1705 0 1 tie_x0
xfeed_1706 0 1 tie_x0
xfeed_1707 0 1 tie_x0
xfeed_1708 0 1 tie_x0
xfeed_1709 0 1 tie_x0
xfeed_219 0 1 tie_x0
xfeed_218 0 1 tie_x0
xfeed_217 0 1 tie_x0
xfeed_216 0 1 tie_x0
xfeed_215 0 1 tie_x0
xfeed_214 0 1 tie_x0
xfeed_213 0 1 tie_x0
xfeed_212 0 1 tie_x0
xfeed_211 0 1 tie_x0
xfeed_210 0 1 tie_x0
xfeed_7089 0 1 tie_x0
xfeed_7088 0 1 tie_x0
xfeed_7087 0 1 tie_x0
xfeed_7086 0 1 tie_x0
xfeed_7085 0 1 tie_x0
xfeed_7084 0 1 tie_x0
xfeed_7083 0 1 tie_x0
xfeed_7082 0 1 tie_x0
xfeed_7081 0 1 tie_x0
xfeed_7080 0 1 tie_x0
xfeed_6559 0 1 tie_x0
xfeed_6558 0 1 tie_x0
xfeed_6557 0 1 tie_x0
xfeed_6556 0 1 tie_x0
xfeed_6555 0 1 tie_x0
xfeed_6554 0 1 tie_x0
xfeed_6553 0 1 tie_x0
xfeed_6552 0 1 tie_x0
xfeed_6551 0 1 tie_x0
xfeed_6550 0 1 tie_x0
xfeed_2249 0 1 tie_x0
xfeed_2248 0 1 tie_x0
xfeed_2247 0 1 tie_x0
xfeed_2246 0 1 tie_x0
xfeed_2245 0 1 tie_x0
xfeed_2244 0 1 tie_x0
xfeed_2243 0 1 tie_x0
xfeed_2242 0 1 tie_x0
xfeed_2241 0 1 tie_x0
xfeed_2240 0 1 tie_x0
xspare_feed_170 0 1 rowend_x0
xspare_feed_171 0 1 tie_x0
xspare_feed_172 0 1 rowend_x0
xspare_feed_173 0 1 rowend_x0
xspare_feed_174 0 1 tie_x0
xspare_feed_175 0 1 rowend_x0
xspare_feed_176 0 1 tie_x0
xfeed_1710 0 1 tie_x0
xfeed_1711 0 1 tie_x0
xfeed_1712 0 1 tie_x0
xfeed_1713 0 1 tie_x0
xfeed_1714 0 1 tie_x0
xfeed_1715 0 1 tie_x0
xfeed_1716 0 1 tie_x0
xfeed_1717 0 1 tie_x0
xfeed_1718 0 1 tie_x0
xfeed_1719 0 1 tie_x0
xfeed_229 0 1 tie_x0
xfeed_228 0 1 tie_x0
xfeed_227 0 1 tie_x0
xfeed_226 0 1 tie_x0
xfeed_225 0 1 tie_x0
xfeed_224 0 1 tie_x0
xfeed_223 0 1 tie_x0
xfeed_222 0 1 tie_x0
xfeed_221 0 1 tie_x0
xfeed_220 0 1 tie_x0
xspare_feed_177 0 1 rowend_x0
xspare_feed_178 0 1 rowend_x0
xspare_feed_179 0 1 tie_x0
xfeed_7099 0 1 tie_x0
xfeed_7098 0 1 tie_x0
xfeed_7097 0 1 tie_x0
xfeed_7096 0 1 tie_x0
xfeed_7095 0 1 tie_x0
xfeed_7094 0 1 tie_x0
xfeed_7093 0 1 tie_x0
xfeed_7092 0 1 tie_x0
xfeed_7091 0 1 tie_x0
xfeed_7090 0 1 tie_x0
xfeed_6569 0 1 tie_x0
xfeed_6568 0 1 tie_x0
xfeed_6567 0 1 tie_x0
xfeed_6566 0 1 tie_x0
xfeed_6565 0 1 tie_x0
xfeed_6564 0 1 tie_x0
xfeed_6563 0 1 tie_x0
xfeed_6562 0 1 tie_x0
xfeed_6561 0 1 tie_x0
xfeed_6560 0 1 tie_x0
xfeed_2259 0 1 tie_x0
xfeed_2258 0 1 tie_x0
xfeed_2257 0 1 tie_x0
xfeed_2256 0 1 tie_x0
xfeed_2255 0 1 tie_x0
xfeed_2254 0 1 tie_x0
xfeed_2253 0 1 tie_x0
xfeed_2252 0 1 tie_x0
xfeed_2251 0 1 rowend_x0
xfeed_2250 0 1 tie_x0
xspare_feed_180 0 1 rowend_x0
xspare_feed_181 0 1 tie_x0
xspare_feed_182 0 1 rowend_x0
xspare_feed_183 0 1 rowend_x0
xfeed_1720 0 1 tie_x0
xfeed_1721 0 1 tie_x0
xfeed_1722 0 1 rowend_x0
xfeed_1723 0 1 tie_x0
xfeed_1724 0 1 tie_x0
xfeed_1725 0 1 tie_x0
xfeed_1726 0 1 tie_x0
xfeed_1727 0 1 tie_x0
xfeed_1728 0 1 tie_x0
xfeed_1729 0 1 tie_x0
xfeed_239 0 1 tie_x0
xfeed_238 0 1 tie_x0
xfeed_237 0 1 tie_x0
xfeed_236 0 1 tie_x0
xfeed_235 0 1 tie_x0
xfeed_234 0 1 tie_x0
xfeed_233 0 1 tie_x0
xfeed_232 0 1 tie_x0
xfeed_231 0 1 tie_x0
xfeed_230 0 1 tie_x0
xsubckt_15_na4_x1 0 1 122 18 13 17 12 na4_x1
xspare_feed_184 0 1 tie_x0
xspare_feed_185 0 1 rowend_x0
xspare_feed_186 0 1 tie_x0
xspare_feed_187 0 1 rowend_x0
xspare_feed_188 0 1 rowend_x0
xspare_feed_189 0 1 tie_x0
xfeed_6576 0 1 tie_x0
xfeed_6575 0 1 tie_x0
xfeed_6574 0 1 tie_x0
xfeed_6573 0 1 tie_x0
xfeed_6572 0 1 tie_x0
xfeed_6571 0 1 tie_x0
xfeed_6570 0 1 tie_x0
xfeed_2269 0 1 tie_x0
xfeed_2268 0 1 tie_x0
xfeed_2267 0 1 tie_x0
xfeed_2266 0 1 tie_x0
xfeed_2265 0 1 tie_x0
xfeed_2264 0 1 tie_x0
xfeed_2263 0 1 tie_x0
xfeed_2262 0 1 tie_x0
xfeed_2261 0 1 tie_x0
xfeed_2260 0 1 tie_x0
xsubckt_22_mx2_x2 0 1 227 8 116 2 mx2_x2
xspare_feed_190 0 1 rowend_x0
xfeed_1730 0 1 tie_x0
xfeed_1731 0 1 tie_x0
xfeed_1732 0 1 tie_x0
xfeed_1733 0 1 tie_x0
xfeed_1734 0 1 tie_x0
xfeed_1735 0 1 tie_x0
xfeed_1736 0 1 tie_x0
xfeed_1737 0 1 tie_x0
xfeed_6579 0 1 tie_x0
xfeed_6578 0 1 tie_x0
xfeed_6577 0 1 tie_x0
xfeed_249 0 1 tie_x0
xfeed_248 0 1 tie_x0
xfeed_247 0 1 tie_x0
xfeed_246 0 1 tie_x0
xfeed_245 0 1 tie_x0
xfeed_244 0 1 tie_x0
xfeed_243 0 1 tie_x0
xfeed_242 0 1 tie_x0
xfeed_241 0 1 tie_x0
xfeed_240 0 1 tie_x0
xspare_feed_191 0 1 tie_x0
xspare_feed_192 0 1 rowend_x0
xspare_feed_193 0 1 rowend_x0
xspare_feed_194 0 1 tie_x0
xspare_feed_195 0 1 rowend_x0
xspare_feed_196 0 1 tie_x0
xspare_feed_197 0 1 rowend_x0
xspare_feed_198 0 1 rowend_x0
xspare_feed_199 0 1 tie_x0
xfeed_0 0 1 tie_x0
xfeed_1738 0 1 tie_x0
xfeed_1739 0 1 tie_x0
xfeed_6583 0 1 tie_x0
xfeed_6582 0 1 tie_x0
xfeed_6581 0 1 tie_x0
xfeed_6580 0 1 tie_x0
xfeed_2279 0 1 tie_x0
xfeed_2278 0 1 tie_x0
xfeed_2277 0 1 tie_x0
xfeed_2276 0 1 tie_x0
xfeed_2275 0 1 tie_x0
xfeed_2274 0 1 tie_x0
xfeed_2273 0 1 tie_x0
xfeed_2272 0 1 tie_x0
xfeed_2271 0 1 tie_x0
xfeed_2270 0 1 tie_x0
xfeed_1 0 1 tie_x0
xfeed_2 0 1 tie_x0
xfeed_3 0 1 tie_x0
xfeed_4 0 1 tie_x0
xfeed_5 0 1 tie_x0
xfeed_6 0 1 tie_x0
xfeed_7 0 1 tie_x0
xfeed_8 0 1 tie_x0
xfeed_9 0 1 tie_x0
xfeed_1740 0 1 tie_x0
xfeed_1741 0 1 tie_x0
xfeed_1742 0 1 rowend_x0
xfeed_1743 0 1 tie_x0
xfeed_1744 0 1 tie_x0
xfeed_6589 0 1 tie_x0
xfeed_6588 0 1 tie_x0
xfeed_6587 0 1 tie_x0
xfeed_6586 0 1 tie_x0
xfeed_6585 0 1 tie_x0
xfeed_6584 0 1 tie_x0
xfeed_259 0 1 tie_x0
xfeed_258 0 1 tie_x0
xfeed_257 0 1 tie_x0
xfeed_256 0 1 tie_x0
xfeed_255 0 1 tie_x0
xfeed_254 0 1 tie_x0
xfeed_253 0 1 tie_x0
xfeed_252 0 1 tie_x0
xfeed_251 0 1 tie_x0
xfeed_250 0 1 tie_x0
xfeed_1745 0 1 tie_x0
xfeed_1746 0 1 tie_x0
xfeed_1747 0 1 tie_x0
xfeed_1748 0 1 tie_x0
xfeed_1749 0 1 tie_x0
xfeed_7209 0 1 tie_x0
xfeed_7208 0 1 tie_x0
xfeed_7207 0 1 tie_x0
xfeed_7206 0 1 tie_x0
xfeed_7205 0 1 tie_x0
xfeed_7204 0 1 tie_x0
xfeed_7203 0 1 tie_x0
xfeed_7202 0 1 tie_x0
xfeed_7201 0 1 tie_x0
xfeed_7200 0 1 tie_x0
xfeed_6590 0 1 tie_x0
xfeed_2289 0 1 tie_x0
xfeed_2288 0 1 tie_x0
xfeed_2287 0 1 tie_x0
xfeed_2286 0 1 tie_x0
xfeed_2285 0 1 tie_x0
xfeed_2284 0 1 tie_x0
xfeed_2283 0 1 tie_x0
xfeed_2282 0 1 tie_x0
xfeed_2281 0 1 tie_x0
xfeed_2280 0 1 tie_x0
xfeed_1750 0 1 tie_x0
xfeed_1751 0 1 tie_x0
xfeed_6599 0 1 tie_x0
xfeed_6598 0 1 tie_x0
xfeed_6597 0 1 tie_x0
xfeed_6596 0 1 tie_x0
xfeed_6595 0 1 tie_x0
xfeed_6594 0 1 tie_x0
xfeed_6593 0 1 tie_x0
xfeed_6592 0 1 tie_x0
xfeed_6591 0 1 tie_x0
xfeed_269 0 1 tie_x0
xfeed_268 0 1 tie_x0
xfeed_267 0 1 tie_x0
xfeed_266 0 1 tie_x0
xfeed_265 0 1 tie_x0
xfeed_264 0 1 tie_x0
xfeed_263 0 1 tie_x0
xfeed_262 0 1 tie_x0
xfeed_261 0 1 tie_x0
xfeed_260 0 1 tie_x0
xfeed_1752 0 1 tie_x0
xfeed_1753 0 1 tie_x0
xfeed_1754 0 1 tie_x0
xfeed_1755 0 1 tie_x0
xfeed_1756 0 1 tie_x0
xfeed_1757 0 1 tie_x0
xfeed_1758 0 1 tie_x0
xfeed_1759 0 1 tie_x0
xfeed_7219 0 1 tie_x0
xfeed_7218 0 1 tie_x0
xfeed_7217 0 1 tie_x0
xfeed_7216 0 1 tie_x0
xfeed_7215 0 1 tie_x0
xfeed_7214 0 1 rowend_x0
xfeed_7213 0 1 tie_x0
xfeed_7212 0 1 tie_x0
xfeed_7211 0 1 tie_x0
xfeed_7210 0 1 tie_x0
xfeed_2297 0 1 tie_x0
xfeed_2296 0 1 tie_x0
xfeed_2295 0 1 tie_x0
xfeed_2294 0 1 tie_x0
xfeed_2293 0 1 tie_x0
xfeed_2292 0 1 tie_x0
xfeed_2291 0 1 tie_x0
xfeed_2290 0 1 tie_x0
xsubckt_122_xr2_x4 0 1 157 77 6 xr2_x4
xfeed_2299 0 1 tie_x0
xfeed_2298 0 1 tie_x0
xfeed_279 0 1 tie_x0
xfeed_278 0 1 tie_x0
xfeed_277 0 1 tie_x0
xfeed_276 0 1 tie_x0
xfeed_275 0 1 tie_x0
xfeed_274 0 1 tie_x0
xfeed_273 0 1 tie_x0
xfeed_272 0 1 tie_x0
xfeed_271 0 1 tie_x0
xfeed_270 0 1 tie_x0
xfeed_1760 0 1 tie_x0
xfeed_1761 0 1 tie_x0
xfeed_1762 0 1 tie_x0
xfeed_1763 0 1 tie_x0
xfeed_1764 0 1 tie_x0
xfeed_1765 0 1 tie_x0
xfeed_1766 0 1 tie_x0
xfeed_1767 0 1 rowend_x0
xfeed_1768 0 1 tie_x0
xfeed_1769 0 1 tie_x0
xfeed_7229 0 1 tie_x0
xfeed_7228 0 1 tie_x0
xfeed_7227 0 1 tie_x0
xfeed_7226 0 1 tie_x0
xfeed_7225 0 1 tie_x0
xfeed_7224 0 1 tie_x0
xfeed_7223 0 1 tie_x0
xfeed_7222 0 1 tie_x0
xfeed_7221 0 1 tie_x0
xfeed_7220 0 1 tie_x0
xfeed_289 0 1 tie_x0
xfeed_288 0 1 tie_x0
xfeed_287 0 1 tie_x0
xfeed_286 0 1 tie_x0
xfeed_285 0 1 tie_x0
xfeed_284 0 1 tie_x0
xfeed_283 0 1 tie_x0
xfeed_282 0 1 tie_x0
xfeed_281 0 1 tie_x0
xfeed_280 0 1 tie_x0
xfeed_1770 0 1 tie_x0
xfeed_1771 0 1 tie_x0
xfeed_1772 0 1 tie_x0
xfeed_1773 0 1 tie_x0
xfeed_1774 0 1 tie_x0
xfeed_1775 0 1 tie_x0
xfeed_1776 0 1 tie_x0
xfeed_1777 0 1 tie_x0
xfeed_1778 0 1 tie_x0
xfeed_1779 0 1 tie_x0
xfeed_7239 0 1 tie_x0
xfeed_7238 0 1 tie_x0
xfeed_7237 0 1 tie_x0
xfeed_7236 0 1 tie_x0
xfeed_7235 0 1 tie_x0
xfeed_7234 0 1 tie_x0
xfeed_7233 0 1 tie_x0
xfeed_7232 0 1 tie_x0
xfeed_7231 0 1 tie_x0
xfeed_7230 0 1 tie_x0
xfeed_6709 0 1 tie_x0
xfeed_6708 0 1 tie_x0
xfeed_6707 0 1 tie_x0
xfeed_6706 0 1 tie_x0
xfeed_6705 0 1 tie_x0
xfeed_6704 0 1 tie_x0
xfeed_6703 0 1 tie_x0
xfeed_6702 0 1 tie_x0
xfeed_6701 0 1 tie_x0
xfeed_6700 0 1 tie_x0
xfeed_299 0 1 tie_x0
xfeed_298 0 1 tie_x0
xfeed_297 0 1 tie_x0
xfeed_296 0 1 tie_x0
xfeed_295 0 1 tie_x0
xfeed_294 0 1 tie_x0
xfeed_293 0 1 tie_x0
xfeed_292 0 1 tie_x0
xfeed_291 0 1 tie_x0
xfeed_290 0 1 tie_x0
xspare_buffer_16 0 1 31 71 buf_x8
xspare_buffer_12 0 1 44 71 buf_x8
xfeed_1780 0 1 tie_x0
xfeed_1781 0 1 tie_x0
xfeed_1782 0 1 tie_x0
xfeed_1783 0 1 tie_x0
xfeed_1784 0 1 tie_x0
xfeed_1785 0 1 tie_x0
xfeed_1786 0 1 tie_x0
xfeed_1787 0 1 tie_x0
xfeed_1788 0 1 tie_x0
xfeed_1789 0 1 tie_x0
xfeed_7249 0 1 tie_x0
xfeed_7248 0 1 tie_x0
xfeed_7247 0 1 tie_x0
xfeed_7246 0 1 tie_x0
xfeed_7245 0 1 tie_x0
xfeed_7244 0 1 tie_x0
xfeed_7243 0 1 tie_x0
xfeed_7242 0 1 tie_x0
xfeed_7241 0 1 tie_x0
xfeed_7240 0 1 tie_x0
xfeed_6716 0 1 tie_x0
xfeed_6715 0 1 tie_x0
xfeed_6714 0 1 tie_x0
xfeed_6713 0 1 tie_x0
xfeed_6712 0 1 tie_x0
xfeed_6711 0 1 tie_x0
xfeed_6710 0 1 tie_x0
xfeed_2409 0 1 tie_x0
xfeed_2408 0 1 tie_x0
xfeed_2407 0 1 tie_x0
xfeed_2406 0 1 tie_x0
xfeed_2405 0 1 tie_x0
xfeed_2404 0 1 tie_x0
xfeed_2403 0 1 tie_x0
xfeed_2402 0 1 tie_x0
xfeed_2401 0 1 tie_x0
xfeed_2400 0 1 tie_x0
xsubckt_43_na3_x1 0 1 95 101 99 98 na3_x1
xsubckt_116_a2_x2 0 1 218 131 163 a2_x2
xfeed_6719 0 1 tie_x0
xfeed_6718 0 1 tie_x0
xfeed_6717 0 1 tie_x0
xspare_buffer_29 0 1 62 70 buf_x8
xspare_buffer_28 0 1 63 70 buf_x8
xspare_buffer_26 0 1 64 70 buf_x8
xspare_buffer_25 0 1 65 70 buf_x8
xspare_buffer_24 0 1 66 70 buf_x8
xspare_buffer_22 0 1 67 70 buf_x8
xspare_buffer_21 0 1 68 70 buf_x8
xspare_buffer_20 0 1 69 70 buf_x8
xfeed_1790 0 1 tie_x0
xfeed_1791 0 1 tie_x0
xfeed_1792 0 1 tie_x0
xfeed_1793 0 1 tie_x0
xfeed_1794 0 1 tie_x0
xfeed_1795 0 1 tie_x0
xfeed_1796 0 1 tie_x0
xfeed_1797 0 1 tie_x0
xfeed_1798 0 1 tie_x0
xfeed_1799 0 1 tie_x0
xfeed_7259 0 1 tie_x0
xfeed_7258 0 1 tie_x0
xfeed_7257 0 1 tie_x0
xfeed_7256 0 1 tie_x0
xfeed_7255 0 1 tie_x0
xfeed_7254 0 1 tie_x0
xfeed_7253 0 1 tie_x0
xfeed_7252 0 1 tie_x0
xfeed_7251 0 1 tie_x0
xfeed_7250 0 1 tie_x0
xfeed_6723 0 1 tie_x0
xfeed_6722 0 1 tie_x0
xfeed_6721 0 1 tie_x0
xfeed_6720 0 1 tie_x0
xfeed_2419 0 1 tie_x0
xfeed_2418 0 1 tie_x0
xfeed_2417 0 1 tie_x0
xfeed_2416 0 1 tie_x0
xfeed_2415 0 1 tie_x0
xfeed_2414 0 1 tie_x0
xfeed_2413 0 1 tie_x0
xfeed_2412 0 1 tie_x0
xfeed_2411 0 1 tie_x0
xfeed_2410 0 1 tie_x0
xfeed_6729 0 1 tie_x0
xfeed_6728 0 1 tie_x0
xfeed_6727 0 1 tie_x0
xfeed_6726 0 1 tie_x0
xfeed_6725 0 1 tie_x0
xfeed_6724 0 1 tie_x0
xspare_buffer_37 0 1 55 57 buf_x8
xspare_buffer_36 0 1 56 57 buf_x8
xspare_buffer_34 0 1 58 70 buf_x8
xspare_buffer_33 0 1 59 70 buf_x8
xspare_buffer_32 0 1 60 70 buf_x8
xspare_buffer_30 0 1 61 70 buf_x8
xfeed_7269 0 1 tie_x0
xfeed_7268 0 1 tie_x0
xfeed_7267 0 1 tie_x0
xfeed_7266 0 1 tie_x0
xfeed_7265 0 1 tie_x0
xfeed_7264 0 1 tie_x0
xfeed_7263 0 1 tie_x0
xfeed_7262 0 1 tie_x0
xfeed_7261 0 1 tie_x0
xfeed_7260 0 1 tie_x0
xfeed_6730 0 1 tie_x0
xfeed_2429 0 1 tie_x0
xfeed_2428 0 1 tie_x0
xfeed_2427 0 1 tie_x0
xfeed_2426 0 1 tie_x0
xfeed_2425 0 1 tie_x0
xfeed_2424 0 1 tie_x0
xfeed_2423 0 1 tie_x0
xfeed_2422 0 1 tie_x0
xfeed_2421 0 1 tie_x0
xfeed_2420 0 1 tie_x0
xspare_buffer_38 0 1 54 57 buf_x8
.ends mac_cts_r
