* tie_diff_w2
* tie_diff_w2
.subckt tie_diff_w2 vdd vss

.ends tie_diff_w2
