* BulkConn_10000WNoUp
.subckt BulkConn_10000WNoUp vdd vss iovdd iovss

.ends BulkConn_10000WNoUp
