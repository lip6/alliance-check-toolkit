* GateDecode
.subckt GateDecode vdd vss iovdd core en ngate pgate
Xtieinst vdd vss tie
Xen_inv vdd vss en en_n inv_x1
Xngate_nor vdd vss ngate_core core en_n nor2_x1
Xngate_levelup vdd iovdd vss ngate_core ngate LevelUp
Xpgate_nand vdd vss pgate_core core en nand2_x1
Xpgate_levelup vdd iovdd vss pgate_core pgate LevelUp
.ends GateDecode
