* nand3_x0
* nand3_x0
.subckt nand3_x0 vdd vss nq i0 i1 i2
Mn0 vss i0 int0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp0 vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
Mn1 int0 i1 int1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp1 nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
Mn2 int1 i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp2 vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
.ends nand3_x0
