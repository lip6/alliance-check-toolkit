-- no model for nexor2_x0
