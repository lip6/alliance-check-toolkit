-- no model for and3_x1
