* Spice description of buf_x2
* Spice driver version 1688526619
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:38

* INTERF i q vdd vss 


.subckt buf_x2 3 2 1 4 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i
* NET 4 = vss
Mtr_00004 2 5 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00003 1 3 5 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00002 4 3 5 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.51U AS=0.1224P AD=0.1224P PS=1.5U PD=1.5U 
Mtr_00001 2 5 4 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C5 1 4 1.17336e-15
C4 2 4 2.15173e-15
C3 3 4 2.41133e-15
C2 4 4 1.17336e-15
C1 5 4 1.31956e-15
.ends buf_x2

