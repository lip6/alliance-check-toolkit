* Spice description of an12_x1
* Spice driver version -952934629
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:32

* INTERF i0 i1 q vdd vss 


.subckt an12_x1 4 2 6 1 5 
* NET 1 = vdd
* NET 2 = i1
* NET 4 = i0
* NET 5 = vss
* NET 6 = q
Mtr_00006 3 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 1 3 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00004 1 4 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00003 3 2 5 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 5 3 6 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 6 4 5 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C6 1 5 1.41822e-15
C5 2 5 2.06462e-15
C4 3 5 1.75845e-15
C3 4 5 1.8384e-15
C2 5 5 1.98312e-15
C1 6 5 2.27334e-15
.ends an12_x1

