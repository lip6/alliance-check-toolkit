* Spice description of a2_x4
* Spice driver version -86868197
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:28

* INTERF i0 i1 q vdd vss 


.subckt a2_x4 4 3 2 1 7 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i1
* NET 4 = i0
* NET 7 = vss
Mtr_00008 1 6 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 2 6 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 1 3 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00005 6 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00004 7 6 2 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 2 6 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 7 3 5 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 5 4 6 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C7 1 7 2.66231e-15
C6 2 7 1.17884e-15
C5 3 7 2.52998e-15
C4 4 7 1.70287e-15
C2 6 7 2.19688e-15
C1 7 7 1.92431e-15
.ends a2_x4

