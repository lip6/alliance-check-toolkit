-- no model for nand3_x0
