* Spice description of na2_x4
* Spice driver version -2002718949
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:49

* INTERF i0 i1 nq vdd vss 


.subckt na2_x4 6 5 3 1 4 
* NET 1 = vdd
* NET 3 = nq
* NET 4 = vss
* NET 5 = i1
* NET 6 = i0
Mtr_00010 1 5 8 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00009 8 6 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00008 3 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 1 2 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 2 8 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00005 4 5 7 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00004 7 6 8 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00003 3 2 4 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00002 2 8 4 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.93U AS=0.2232P AD=0.2232P PS=2.35U PD=2.35U 
Mtr_00001 4 2 3 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
C8 1 4 2.22964e-15
C7 2 4 2.01418e-15
C6 3 4 1.79621e-15
C5 4 4 2.20855e-15
C4 5 4 1.79868e-15
C3 6 4 1.78955e-15
C1 8 4 2.63736e-15
.ends na2_x4

