-- no model for nand2_x1
