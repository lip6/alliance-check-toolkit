* nand2_x1
.subckt nand2_x1 vdd vss nq i0 i1
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
Mi1_nmos _net0 i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
.ends nand2_x1
