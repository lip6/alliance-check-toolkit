* and21nor_x1
* and21nor_x1
.subckt and21nor_x1 vdd vss nq i0 i1 i2
Mi0_nmos vss i0 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi0_pmos _net0 i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
Mi1_nmos _net1 i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi1_pmos vdd i1 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
Mi2_nmos nq i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi2_pmos _net0 i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
.ends and21nor_x1
