sky130_fd_sc_hd__inv_4_chain 10 inv_4_hitas with slope 
*
* from
* top_sky130_fd_sc_hd__inv_4_chain.spi
* ngspice simulation
* 

*****************

.TEMP 25

******************
******************
* BSIM4 transistor model parameters for ngspice
*
* nfet_01v8
*.include sky130_fd_pr__nfet_01v8__mismatch.corner.spice
*.include sky130_fd_pr__nfet_01v8__tt.corner.spice
* pfet_01v8_hvt
*.include sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
*.include sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice

*******************************

*******************************
*Simulation conditions

Vground evss 0 0
Vsupply evdd 0 DC 1.8

******************
* circuit model
* include circuit netlist
.INCLUDE sky130_fd_sc_hd__inv_4_chain.spi
*****************

*****************
* Circuit Instantiation
*.subckt sky130_fd_sc_hd__inv_4_chain in out vdd gnd
* 10 inverters
Xinv_4_chain in out evdd evss sky130_fd_sc_hd__inv_4_chain



.end

