-- no model for IOPadIOVdd
