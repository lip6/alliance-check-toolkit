* Filler400
.subckt Filler400 vss vdd iovss iovdd
Xbulkconn vdd vss iovdd iovss BulkConn_400WNoUp
.ends Filler400
