* nor4_x0
* nor4_x0
.subckt nor4_x0 vdd vss nq i0 i1 i2 i3
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi0_pmos vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi1_pmos _net0 i1 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi2_nmos vss i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi2_pmos _net1 i2 _net2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi3_nmos nq i3 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi3_pmos _net2 i3 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends nor4_x0
