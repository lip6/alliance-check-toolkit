-- no model for or2_x1
