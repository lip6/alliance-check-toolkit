* Spice description of nd2abv0x05
* Spice driver version -8806629
* Date ( dd/mm/yyyy hh:mm:ss ): 23/06/2024 at 14:07:17

* INTERF a b vdd vss z 


.subckt nd2abv0x05 2 5 1 6 7 
* NET 1 = vdd
* NET 2 = a
* NET 3 = an
* NET 4 = 08
* NET 5 = b
* NET 6 = vss
* NET 7 = z
* NET 8 = bn
M03 1 5 8 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.9U AS=0.333P AD=0.333P PS=2.55U PD=2.55U 
M07 7 8 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.9U AS=0.333P AD=0.333P PS=2.55U PD=2.55U 
M05 1 3 7 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.9U AS=0.333P AD=0.333P PS=2.55U PD=2.55U 
M01 3 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.9U AS=0.333P AD=0.333P PS=2.55U PD=2.55U 
M04 6 5 8 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.45U AS=0.1665P AD=0.1665P PS=1.65U PD=1.65U 
M08 4 8 7 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.2775P AD=0.2775P PS=2.25U PD=2.25U 
M06 6 3 4 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.2775P AD=0.2775P PS=2.25U PD=2.25U 
M02 3 2 6 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.45U AS=0.1665P AD=0.1665P PS=1.65U PD=1.65U 
C8 1 6 2.59971e-15
C7 2 6 8.98131e-16
C6 3 6 1.46816e-15
C4 5 6 1.19538e-15
C3 6 6 2.64363e-15
C2 7 6 1.54618e-15
C1 8 6 1.51773e-15
.ends nd2abv0x05

