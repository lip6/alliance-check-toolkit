-- no model for inv_x2
