-- no model for inv_x1
