* DP8TArray_16X16
.subckt DP8TArray_16X16 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_16X8
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X8
.ends DP8TArray_16X16
