-- no model for nand4_x1
