* diode_sf
.param
+ sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult=7.9012e-01 
+ sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult=9.1728e-01 
+ sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult=7.0406e-01 
+ sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult=0.69 
+ sky130_fd_pr__nfet_01v8__ajunction_mult=0.7739
+ sky130_fd_pr__nfet_01v8__pjunction_mult=0.79336
+ sky130_fd_pr__pfet_01v8__ajunction_mult=1.0909
+ sky130_fd_pr__pfet_01v8__pjunction_mult=1.096
