* powmid_x0
.subckt powmid_x0 vss vdd

.ends powmid_x0
