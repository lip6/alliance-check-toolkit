* Spice description of noa2a2a23_x1
* Spice driver version 2096709403
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:09

* INTERF i0 i1 i2 i3 i4 i5 nq vdd vss 


.subckt noa2a2a23_x1 4 5 7 8 10 11 12 1 14 
* NET 1 = vdd
* NET 4 = i0
* NET 5 = i1
* NET 7 = i2
* NET 8 = i3
* NET 10 = i4
* NET 11 = i5
* NET 12 = nq
* NET 14 = vss
Mtr_00012 1 4 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 2 5 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 2 8 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 3 10 12 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 12 11 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 3 7 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 14 4 6 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 6 5 12 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 14 7 9 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 9 8 12 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 12 10 13 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 13 11 14 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C14 1 14 3.12982e-15
C13 2 14 7.71835e-16
C12 3 14 7.92919e-16
C11 4 14 1.39425e-15
C10 5 14 1.39425e-15
C8 7 14 1.63156e-15
C7 8 14 1.5886e-15
C5 10 14 1.52203e-15
C4 11 14 1.4764e-15
C3 12 14 2.64749e-15
C1 14 14 2.78018e-15
.ends noa2a2a23_x1

