* BulkConn_400WNoUp
* BulkConn_400WNoUp
.subckt BulkConn_400WNoUp vdd vss iovdd iovss

.ends BulkConn_400WNoUp
