* Corner
* Corner
.subckt Corner vss vdd iovss iovdd

.ends Corner
