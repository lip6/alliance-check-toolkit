* GuardRing_N17368W8096HTF
.subckt GuardRing_N17368W8096HTF conn

.ends GuardRing_N17368W8096HTF
