* Spice description of inv_x8
* Spice driver version -1171701989
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:43

* INTERF i nq vdd vss 


.subckt inv_x8 3 5 1 4 
* NET 1 = vdd
* NET 3 = i
* NET 4 = vss
* NET 5 = nq
Mtr_00008 5 3 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 1 3 5 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 2 3 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 1 3 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00004 5 3 4 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 4 3 5 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 2 3 4 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 4 3 2 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C5 1 4 3.10868e-15
C4 2 4 1.17884e-15
C3 3 4 3.54572e-15
C2 4 4 2.29468e-15
C1 5 4 2.33414e-15
.ends inv_x8

