* Spice description of tie_x0
* Spice driver version -1553649893
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:30:04

* INTERF vdd vss 


.subckt tie_x0 1 2 
* NET 1 = vdd
* NET 2 = vss
C2 1 2 1.44526e-15
C1 2 2 1.21917e-15
.ends tie_x0

