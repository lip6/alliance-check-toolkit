../rtl/inc16.vhdl