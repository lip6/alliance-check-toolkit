* DP8TArray_32X32
.subckt DP8TArray_32X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_32X16
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X16
.ends DP8TArray_32X32
