* Spice description of zero_x0
* Spice driver version 76410651
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:46

* INTERF nq vdd vss 


.subckt zero_x0 3 1 2 
* NET 1 = vdd
* NET 2 = vss
* NET 3 = nq
Mtr_00001 3 1 2 2 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C3 1 2 2.28992e-15
C2 2 2 1.4282e-15
C1 3 2 1.99727e-15
.ends zero_x0

