* Spice description of nxr2_x4
* Spice driver version -1548132581
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:19

* INTERF i0 i1 nq vdd vss 


.subckt nxr2_x4 9 5 3 2 10 
* NET 2 = vdd
* NET 3 = nq
* NET 5 = i1
* NET 9 = i0
* NET 10 = vss
Mtr_00016 2 7 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00015 3 7 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00014 2 5 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 1 11 7 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 1 9 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 7 4 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 4 5 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00009 2 9 11 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00008 10 7 3 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00007 3 7 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00006 4 5 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00005 10 9 11 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00004 8 11 7 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 10 4 8 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 7 5 6 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 6 9 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C11 1 10 5.28612e-16
C10 2 10 4.30428e-15
C9 3 10 2.15173e-15
C8 4 10 1.92318e-15
C7 5 10 2.78088e-15
C5 7 10 3.28518e-15
C3 9 10 2.54824e-15
C2 10 10 3.49027e-15
C1 11 10 1.51574e-15
.ends nxr2_x4

