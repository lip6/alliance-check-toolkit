* nsnrlatch_x0
* nsnrlatch_x0
.subckt nsnrlatch_x0 vdd vss nset nrst q nq
Mnset_nmos q nset _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnset_pmos vdd nset q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnq_nmos _net0 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnq_pmos q q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mq_nmos vss q _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mq_pmos vdd q nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnrst_nmos _net1 nset nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnrst_pmos nq nset vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nsnrlatch_x0
