../adder.vhdl