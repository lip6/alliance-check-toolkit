* Spice description of nmx3_x1
* Spice driver version -728613093
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:59

* INTERF cmd0 cmd1 i0 i1 i2 nq vdd vss 


.subckt nmx3_x1 7 16 6 8 13 14 5 18 
* NET 5 = vdd
* NET 6 = i0
* NET 7 = cmd0
* NET 8 = i1
* NET 13 = i2
* NET 14 = nq
* NET 16 = cmd1
* NET 18 = vss
Mtr_00018 5 9 4 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00017 4 8 2 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00016 12 16 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00015 3 13 4 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00014 14 16 3 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00013 2 12 14 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00012 1 7 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00011 14 6 1 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00010 5 7 9 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00009 10 9 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00008 12 16 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.68U AS=0.1632P AD=0.1632P PS=1.84U PD=1.84U 
Mtr_00007 18 7 9 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.68U AS=0.1632P AD=0.1632P PS=1.84U PD=1.84U 
Mtr_00006 14 12 15 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00005 15 13 17 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00004 14 6 10 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00003 18 7 17 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00002 17 8 11 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00001 11 16 14 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
C15 4 18 8.63043e-16
C14 5 18 3.66092e-15
C13 6 18 1.36556e-15
C12 7 18 2.01198e-15
C11 8 18 1.14216e-15
C10 9 18 1.84566e-15
C7 12 18 1.92755e-15
C6 13 18 9.62699e-16
C5 14 18 3.71747e-15
C3 16 18 2.15016e-15
C2 17 18 8.02238e-16
C1 18 18 3.6212e-15
.ends nmx3_x1

