*
* sky130_fd_sc_hd__inv_4_3.spi
* 

* sky130_fd_sc_hd__inv_4
*.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y

.INCLUDE sky130_fd_sc_hd__inv_4.spice

.subckt sky130_fd_sc_hd__inv_4_3 in out vdd gnd
Xa in gnd gnd vdd vdd n1   sky130_fd_sc_hd__inv_4
Xb n1 gnd gnd vdd vdd n2   sky130_fd_sc_hd__inv_4
Xc n2 gnd gnd vdd vdd out  sky130_fd_sc_hd__inv_4
.ends sky130_fd_sc_hd__inv_4_3


