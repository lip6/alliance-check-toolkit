* Spice description of arlet6502_cts_r_transistors_ihp
* Spice driver version 66370477
* Date ( dd/mm/yyyy hh:mm:ss ): 30/09/2024 at 15:11:36

* INTERF a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] a[9] a[10] a[11] a[12] 
* INTERF a[13] a[14] a[15] clk di[0] di[1] di[2] di[3] di[4] di[5] di[6] 
* INTERF di[7] do[0] do[1] do[2] do[3] do[4] do[5] do[6] do[7] irq nmi rdy 
* INTERF reset vdd vss we 


.subckt arlet6502_cts_r_transistors_ihp 3441 2148 2281 5601 3866 5146 4490 4083 3281 8768 8741 8716 8688 8665 8646 8617 4311 8585 8566 7928 7071 6701 6410 6234 4305 2939 1876 1118 943 7826 6975 6138 5341 4751 2187 4158 3158 8552 8787 1215 
* NET 55 = subckt_1650_sff1_x4.sff_s
* NET 59 = subckt_1650_sff1_x4.sff_m
* NET 61 = subckt_1650_sff1_x4.ckr
* NET 63 = subckt_1650_sff1_x4.nckr
* NET 67 = subckt_1620_sff1_x4.sff_s
* NET 71 = subckt_1620_sff1_x4.sff_m
* NET 73 = subckt_1620_sff1_x4.ckr
* NET 74 = subckt_1620_sff1_x4.nckr
* NET 75 = abc_11867_auto_rtlil_cc_2608_muxgate_11610
* NET 82 = subckt_1634_sff1_x4.sff_s
* NET 86 = subckt_1634_sff1_x4.sff_m
* NET 89 = subckt_1634_sff1_x4.ckr
* NET 90 = subckt_1634_sff1_x4.nckr
* NET 94 = subckt_1622_sff1_x4.sff_s
* NET 97 = subckt_1622_sff1_x4.sff_m
* NET 99 = subckt_1622_sff1_x4.ckr
* NET 101 = subckt_1622_sff1_x4.nckr
* NET 103 = subckt_1649_sff1_x4.sff_s
* NET 106 = subckt_1649_sff1_x4.sff_m
* NET 111 = subckt_1649_sff1_x4.ckr
* NET 112 = subckt_1649_sff1_x4.nckr
* NET 115 = subckt_1619_sff1_x4.sff_s
* NET 119 = subckt_1619_sff1_x4.sff_m
* NET 121 = subckt_1619_sff1_x4.ckr
* NET 123 = subckt_1619_sff1_x4.nckr
* NET 125 = subckt_1633_sff1_x4.sff_s
* NET 128 = subckt_1633_sff1_x4.sff_m
* NET 133 = subckt_1633_sff1_x4.ckr
* NET 134 = subckt_1633_sff1_x4.nckr
* NET 137 = subckt_1618_sff1_x4.sff_s
* NET 142 = subckt_1618_sff1_x4.sff_m
* NET 143 = subckt_1618_sff1_x4.ckr
* NET 145 = subckt_1618_sff1_x4.nckr
* NET 148 = subckt_1621_sff1_x4.sff_s
* NET 152 = subckt_1621_sff1_x4.sff_m
* NET 154 = subckt_1621_sff1_x4.ckr
* NET 156 = subckt_1621_sff1_x4.nckr
* NET 168 = abc_11867_new_n485
* NET 175 = abc_11867_new_n872
* NET 177 = abc_11867_new_n873
* NET 179 = abc_11867_new_n875
* NET 181 = abc_11867_new_n868
* NET 185 = abc_11867_new_n428
* NET 190 = abc_11867_new_n473
* NET 193 = abc_11867_new_n430_hfns_2
* NET 195 = abc_11867_new_n430
* NET 198 = abc_11867_new_n431
* NET 248 = subckt_1653_sff1_x4.sff_s
* NET 253 = subckt_1653_sff1_x4.sff_m
* NET 256 = subckt_1653_sff1_x4.ckr
* NET 257 = subckt_1653_sff1_x4.nckr
* NET 259 = abc_11867_auto_rtlil_cc_2608_muxgate_11658
* NET 264 = subckt_1623_sff1_x4.sff_s
* NET 269 = subckt_1623_sff1_x4.sff_m
* NET 271 = subckt_1623_sff1_x4.ckr
* NET 273 = subckt_1623_sff1_x4.nckr
* NET 274 = mos6502_axys_2_3
* NET 276 = mos6502_axys_3_3
* NET 281 = subckt_1652_sff1_x4.sff_s
* NET 285 = subckt_1652_sff1_x4.sff_m
* NET 288 = subckt_1652_sff1_x4.ckr
* NET 290 = subckt_1652_sff1_x4.nckr
* NET 291 = abc_11867_auto_rtlil_cc_2608_muxgate_11662
* NET 297 = subckt_1636_sff1_x4.sff_s
* NET 301 = subckt_1636_sff1_x4.sff_m
* NET 304 = subckt_1636_sff1_x4.ckr
* NET 306 = subckt_1636_sff1_x4.nckr
* NET 307 = abc_11867_auto_rtlil_cc_2608_muxgate_11656
* NET 313 = abc_11867_auto_rtlil_cc_2608_muxgate_11608
* NET 318 = subckt_1648_sff1_x4.sff_s
* NET 322 = subckt_1648_sff1_x4.sff_m
* NET 326 = subckt_1648_sff1_x4.nckr
* NET 327 = subckt_1648_sff1_x4.ckr
* NET 328 = abc_11867_auto_rtlil_cc_2608_muxgate_11654
* NET 333 = abc_11867_auto_rtlil_cc_2608_muxgate_11606
* NET 338 = abc_11867_auto_rtlil_cc_2608_muxgate_11612
* NET 349 = subckt_1632_sff1_x4.sff_s
* NET 354 = subckt_1632_sff1_x4.sff_m
* NET 356 = abc_11867_auto_rtlil_cc_2608_muxgate_11622
* NET 358 = subckt_1632_sff1_x4.ckr
* NET 359 = subckt_1632_sff1_x4.nckr
* NET 360 = abc_11867_new_n1410
* NET 363 = abc_11867_new_n1411
* NET 369 = abc_11867_new_n640
* NET 372 = abc_11867_new_n476
* NET 374 = abc_11867_new_n864
* NET 378 = abc_11867_new_n877
* NET 382 = abc_11867_new_n871
* NET 388 = abc_11867_new_n878
* NET 391 = abc_11867_new_n862
* NET 396 = abc_11867_new_n471
* NET 398 = abc_11867_new_n471_hfns_3
* NET 415 = abc_11867_new_n608
* NET 416 = abc_11867_new_n431_hfns_2
* NET 418 = abc_11867_new_n482
* NET 492 = abc_11867_new_n1424
* NET 498 = abc_11867_new_n521
* NET 499 = abc_11867_new_n522
* NET 502 = abc_11867_auto_rtlil_cc_2608_muxgate_11664
* NET 510 = subckt_1624_sff1_x4.sff_s
* NET 512 = subckt_1624_sff1_x4.sff_m
* NET 515 = subckt_1624_sff1_x4.ckr
* NET 516 = subckt_1624_sff1_x4.nckr
* NET 517 = abc_11867_auto_rtlil_cc_2608_muxgate_11616
* NET 524 = subckt_1637_sff1_x4.sff_s
* NET 528 = subckt_1637_sff1_x4.sff_m
* NET 530 = subckt_1637_sff1_x4.ckr
* NET 531 = subckt_1637_sff1_x4.nckr
* NET 532 = mos6502_axys_0_3
* NET 534 = abc_11867_auto_rtlil_cc_2608_muxgate_11626
* NET 538 = mos6502_axys_2_5
* NET 542 = mos6502_axys_3_5
* NET 543 = abc_11867_auto_rtlil_cc_2608_muxgate_11614
* NET 548 = mos6502_axys_0_5
* NET 550 = abc_11867_auto_rtlil_cc_2608_muxgate_11630
* NET 554 = mos6502_axys_3_2
* NET 555 = mos6502_axys_2_2
* NET 559 = abc_11867_auto_rtlil_cc_2608_muxgate_11624
* NET 560 = mos6502_axys_0_2
* NET 571 = subckt_1617_sff1_x4.sff_s
* NET 575 = subckt_1617_sff1_x4.sff_m
* NET 576 = subckt_1617_sff1_x4.ckr
* NET 578 = subckt_1617_sff1_x4.nckr
* NET 581 = subckt_1651_sff1_x4.sff_s
* NET 584 = subckt_1651_sff1_x4.sff_m
* NET 587 = subckt_1651_sff1_x4.ckr
* NET 588 = subckt_1651_sff1_x4.nckr
* NET 591 = subckt_1635_sff1_x4.sff_s
* NET 594 = subckt_1635_sff1_x4.sff_m
* NET 597 = subckt_1635_sff1_x4.ckr
* NET 598 = subckt_1635_sff1_x4.nckr
* NET 599 = abc_11867_new_n1421
* NET 602 = abc_11867_new_n639
* NET 608 = abc_11867_new_n1426
* NET 609 = abc_11867_new_n856
* NET 612 = abc_11867_new_n865
* NET 613 = abc_11867_new_n874
* NET 614 = abc_11867_new_n867
* NET 616 = abc_11867_new_n876
* NET 621 = abc_11867_new_n473_hfns_3
* NET 625 = abc_11867_new_n525
* NET 628 = abc_11867_new_n608_hfns_2
* NET 632 = abc_11867_new_n478
* NET 638 = abc_11867_new_n426
* NET 680 = abc_11867_auto_rtlil_cc_2608_muxgate_11620
* NET 684 = abc_11867_new_n1425
* NET 699 = subckt_1654_sff1_x4.sff_s
* NET 700 = subckt_1654_sff1_x4.sff_m
* NET 706 = subckt_1654_sff1_x4.nckr
* NET 707 = subckt_1654_sff1_x4.ckr
* NET 708 = abc_11867_auto_rtlil_cc_2608_muxgate_11666
* NET 715 = abc_11867_auto_rtlil_cc_2608_muxgate_11618
* NET 720 = mos6502_axys_3_6
* NET 721 = mos6502_axys_2_6
* NET 726 = mos6502_axys_0_6
* NET 728 = abc_11867_auto_rtlil_cc_2608_muxgate_11632
* NET 736 = subckt_1644_sff1_x4.sff_s
* NET 737 = subckt_1644_sff1_x4.sff_m
* NET 745 = subckt_1644_sff1_x4.nckr
* NET 746 = subckt_1644_sff1_x4.ckr
* NET 751 = subckt_1631_sff1_x4.sff_s
* NET 752 = subckt_1631_sff1_x4.sff_m
* NET 759 = subckt_1631_sff1_x4.ckr
* NET 761 = subckt_1631_sff1_x4.nckr
* NET 764 = mos6502_axys_3_1
* NET 765 = mos6502_axys_2_1
* NET 767 = mos6502_axys_0_1
* NET 777 = abc_11867_auto_rtlil_cc_2608_muxgate_11628
* NET 779 = abc_11867_new_n1148
* NET 783 = abc_11867_new_n1427
* NET 786 = abc_11867_new_n1418
* NET 792 = abc_11867_new_n1409
* NET 793 = abc_11867_new_n1414
* NET 794 = abc_11867_new_n1412
* NET 795 = abc_11867_new_n1413
* NET 800 = abc_11867_new_n654
* NET 802 = abc_11867_new_n1407
* NET 805 = abc_11867_new_n863
* NET 807 = abc_11867_new_n860
* NET 815 = abc_11867_new_n475
* NET 817 = abc_11867_new_n490
* NET 824 = abc_11867_new_n518
* NET 827 = abc_11867_new_n516
* NET 831 = abc_11867_new_n478_hfns_3
* NET 835 = abc_11867_new_n514_hfns_2
* NET 836 = abc_11867_new_n514
* NET 911 = subckt_1642_sff1_x4.sff_s
* NET 914 = subckt_1642_sff1_x4.sff_m
* NET 918 = subckt_1642_sff1_x4.ckr
* NET 919 = subckt_1642_sff1_x4.nckr
* NET 920 = abc_11867_auto_rtlil_cc_2608_muxgate_11642
* NET 925 = mos6502_axys_3_7
* NET 926 = mos6502_axys_2_7
* NET 931 = mos6502_axys_0_7
* NET 933 = subckt_1638_sff1_x4.sff_s
* NET 935 = subckt_1638_sff1_x4.sff_m
* NET 937 = abc_11867_auto_rtlil_cc_2608_muxgate_11634
* NET 940 = subckt_1638_sff1_x4.nckr
* NET 941 = subckt_1638_sff1_x4.ckr
* NET 943 = do[3]
* NET 944 = abc_11867_auto_rtlil_cc_2608_muxgate_11646
* NET 951 = subckt_1641_sff1_x4.sff_s
* NET 955 = subckt_1641_sff1_x4.sff_m
* NET 956 = subckt_1641_sff1_x4.ckr
* NET 958 = subckt_1641_sff1_x4.nckr
* NET 959 = mos6502_axys_1_2
* NET 960 = abc_11867_auto_rtlil_cc_2608_muxgate_11640
* NET 967 = subckt_1647_sff1_x4.sff_s
* NET 971 = subckt_1647_sff1_x4.sff_m
* NET 972 = subckt_1647_sff1_x4.ckr
* NET 974 = subckt_1647_sff1_x4.nckr
* NET 975 = abc_11867_auto_rtlil_cc_2608_muxgate_11652
* NET 980 = abc_11867_auto_rtlil_cc_2608_muxgate_11604
* NET 983 = abc_11867_new_n1103
* NET 986 = abc_11867_auto_rtlil_cc_2608_muxgate_11660
* NET 988 = abc_11867_new_n1166
* NET 992 = mos6502_axys_3_4
* NET 993 = mos6502_axys_2_4
* NET 994 = mos6502_axys_0_4
* NET 1001 = subckt_1643_sff1_x4.sff_s
* NET 1004 = subckt_1643_sff1_x4.sff_m
* NET 1005 = subckt_1643_sff1_x4.ckr
* NET 1007 = subckt_1643_sff1_x4.nckr
* NET 1009 = abc_11867_new_n383
* NET 1011 = abc_11867_new_n479
* NET 1013 = abc_11867_new_n1417
* NET 1015 = abc_11867_new_n429
* NET 1016 = abc_11867_new_n500
* NET 1019 = abc_11867_new_n1423
* NET 1020 = abc_11867_new_n859
* NET 1021 = abc_11867_new_n858
* NET 1030 = abc_11867_new_n641
* NET 1034 = abc_11867_new_n638
* NET 1037 = abc_11867_new_n527
* NET 1044 = abc_11867_new_n426_hfns_2
* NET 1046 = abc_11867_new_n482_hfns_2
* NET 1076 = subckt_1645_sff1_x4.sff_s
* NET 1080 = subckt_1645_sff1_x4.sff_m
* NET 1084 = subckt_1645_sff1_x4.ckr
* NET 1085 = subckt_1645_sff1_x4.nckr
* NET 1092 = mos6502_axys_1_3
* NET 1095 = spare_buffer_82.q
* NET 1100 = abc_11867_new_n909
* NET 1105 = mos6502_axys_1_5
* NET 1113 = abc_11867_new_n901
* NET 1114 = abc_11867_new_n900
* NET 1116 = abc_11867_new_n902
* NET 1118 = do[2]
* NET 1119 = abc_11867_new_n991
* NET 1121 = spare_buffer_78.q
* NET 1123 = abc_11867_new_n881
* NET 1124 = mos6502_axys_3_0
* NET 1125 = mos6502_axys_2_0
* NET 1127 = mos6502_axys_0_0
* NET 1128 = abc_11867_new_n882
* NET 1129 = abc_11867_new_n883
* NET 1135 = abc_11867_new_n916
* NET 1138 = abc_11867_new_n915
* NET 1140 = mos6502_axys_1_4
* NET 1141 = abc_11867_auto_rtlil_cc_2608_muxgate_11644
* NET 1147 = abc_11867_new_n1415
* NET 1149 = abc_11867_new_n1420
* NET 1151 = abc_11867_new_n1419
* NET 1154 = abc_11867_new_n600
* NET 1159 = abc_11867_new_n1467
* NET 1166 = spare_buffer_66.q
* NET 1173 = abc_11867_new_n475_hfns_3
* NET 1180 = abc_11867_new_n490_hfns_2
* NET 1189 = abc_11867_new_n606
* NET 1193 = abc_11867_new_n605
* NET 1199 = spare_buffer_62.q
* NET 1201 = abc_11867_new_n665
* NET 1202 = abc_11867_new_n664
* NET 1203 = mos6502_state[2]
* NET 1204 = subckt_1627_sff1_x4.sff_s
* NET 1210 = subckt_1627_sff1_x4.sff_m
* NET 1212 = subckt_1627_sff1_x4.ckr
* NET 1214 = subckt_1627_sff1_x4.nckr
* NET 1215 = we
* NET 1280 = mos6502_axys_1_7
* NET 1281 = subckt_1646_sff1_x4.sff_s
* NET 1286 = abc_11867_auto_rtlil_cc_2608_muxgate_11650
* NET 1288 = subckt_1646_sff1_x4.sff_m
* NET 1290 = subckt_1646_sff1_x4.ckr
* NET 1291 = subckt_1646_sff1_x4.nckr
* NET 1292 = abc_11867_auto_rtlil_cc_2608_muxgate_11648
* NET 1297 = mos6502_axys_1_6
* NET 1300 = spare_buffer_81.q
* NET 1302 = clk_root_tr_tr_0
* NET 1308 = abc_11867_new_n1792
* NET 1309 = abc_11867_new_n1796
* NET 1310 = abc_11867_new_n1830
* NET 1318 = abc_11867_new_n1829
* NET 1323 = abc_11867_new_n1817
* NET 1325 = abc_11867_new_n1821
* NET 1333 = abc_11867_new_n1854
* NET 1335 = spare_buffer_77.q
* NET 1338 = abc_11867_new_n917
* NET 1339 = abc_11867_new_n914
* NET 1347 = subckt_1640_sff1_x4.sff_s
* NET 1350 = subckt_1640_sff1_x4.sff_m
* NET 1355 = subckt_1640_sff1_x4.ckr
* NET 1356 = subckt_1640_sff1_x4.nckr
* NET 1358 = abc_11867_new_n1465
* NET 1362 = abc_11867_new_n1468
* NET 1363 = abc_11867_new_n663
* NET 1364 = abc_11867_new_n1466
* NET 1365 = spare_buffer_65.q
* NET 1367 = clk_root_tl_tr_0
* NET 1369 = abc_11867_new_n380
* NET 1372 = abc_11867_new_n599
* NET 1373 = abc_11867_new_n602
* NET 1381 = abc_11867_new_n659
* NET 1382 = abc_11867_new_n660
* NET 1386 = spare_buffer_61.q
* NET 1390 = mos6502_state[0]
* NET 1391 = subckt_1625_sff1_x4.sff_s
* NET 1394 = subckt_1625_sff1_x4.sff_m
* NET 1399 = subckt_1625_sff1_x4.ckr
* NET 1400 = subckt_1625_sff1_x4.nckr
* NET 1447 = abc_11867_new_n1807
* NET 1455 = abc_11867_new_n1806
* NET 1456 = abc_11867_new_n1804
* NET 1462 = abc_11867_new_n907
* NET 1463 = abc_11867_new_n908
* NET 1476 = abc_11867_new_n1816
* NET 1477 = abc_11867_new_n1831
* NET 1479 = abc_11867_new_n1855
* NET 1487 = abc_11867_new_n1851
* NET 1489 = abc_11867_new_n1853
* NET 1496 = abc_11867_new_n1684
* NET 1498 = abc_11867_new_n1874
* NET 1505 = mos6502_axys_1_0
* NET 1506 = subckt_1639_sff1_x4.sff_s
* NET 1509 = subckt_1639_sff1_x4.sff_m
* NET 1513 = abc_11867_auto_rtlil_cc_2608_muxgate_11636
* NET 1516 = clk_root_tr_tl_0
* NET 1517 = subckt_1639_sff1_x4.ckr
* NET 1518 = subckt_1639_sff1_x4.nckr
* NET 1521 = abc_11867_auto_rtlil_cc_2608_muxgate_11638
* NET 1522 = mos6502_axys_1_1
* NET 1525 = abc_11867_new_n1157
* NET 1535 = abc_11867_new_n1434
* NET 1537 = abc_11867_new_n1668
* NET 1538 = abc_11867_new_n1422
* NET 1539 = abc_11867_new_n1408
* NET 1546 = abc_11867_new_n766
* NET 1552 = abc_11867_new_n604
* NET 1553 = abc_11867_new_n656
* NET 1558 = abc_11867_new_n857
* NET 1564 = abc_11867_new_n690
* NET 1566 = abc_11867_new_n689
* NET 1567 = mos6502_state[5]
* NET 1568 = subckt_1630_sff1_x4.sff_s
* NET 1574 = subckt_1630_sff1_x4.sff_m
* NET 1576 = subckt_1630_sff1_x4.ckr
* NET 1578 = subckt_1630_sff1_x4.nckr
* NET 1586 = abc_11867_new_n738
* NET 1590 = abc_11867_new_n657
* NET 1591 = abc_11867_new_n735
* NET 1592 = abc_11867_new_n736
* NET 1596 = abc_11867_new_n729
* NET 1599 = abc_11867_new_n666
* NET 1602 = abc_11867_new_n726
* NET 1641 = abc_11867_new_n658
* NET 1702 = abc_11867_new_n1811
* NET 1706 = abc_11867_new_n1809
* NET 1709 = abc_11867_new_n1801
* NET 1710 = abc_11867_new_n1808
* NET 1712 = abc_11867_new_n1805
* NET 1716 = abc_11867_new_n1797
* NET 1717 = abc_11867_new_n1803
* NET 1722 = abc_11867_new_n1802
* NET 1723 = abc_11867_new_n1836
* NET 1725 = abc_11867_new_n1840
* NET 1729 = abc_11867_new_n1839
* NET 1732 = abc_11867_new_n1827
* NET 1737 = abc_11867_new_n1856
* NET 1738 = abc_11867_new_n1860
* NET 1741 = abc_11867_new_n1849
* NET 1744 = abc_11867_new_n1852
* NET 1747 = abc_11867_new_n1876
* NET 1753 = abc_11867_new_n895
* NET 1755 = abc_11867_new_n1846
* NET 1757 = abc_11867_new_n893
* NET 1758 = abc_11867_new_n894
* NET 1760 = abc_11867_new_n485_hfns_4
* NET 1763 = abc_11867_new_n951
* NET 1765 = abc_11867_new_n966
* NET 1766 = abc_11867_new_n965
* NET 1768 = abc_11867_new_n768
* NET 1769 = abc_11867_new_n855
* NET 1771 = abc_11867_new_n1667
* NET 1772 = abc_11867_new_n598
* NET 1777 = abc_11867_new_n775
* NET 1781 = abc_11867_new_n567
* NET 1783 = abc_11867_new_n603
* NET 1790 = abc_11867_new_n645
* NET 1791 = abc_11867_new_n644
* NET 1793 = abc_11867_new_n661
* NET 1794 = abc_11867_new_n825
* NET 1795 = abc_11867_new_n823
* NET 1798 = abc_11867_new_n652
* NET 1805 = subckt_1628_sff1_x4.sff_s
* NET 1809 = subckt_1628_sff1_x4.sff_m
* NET 1811 = subckt_1628_sff1_x4.nckr
* NET 1812 = subckt_1628_sff1_x4.ckr
* NET 1862 = abc_11867_new_n1826
* NET 1870 = abc_11867_new_n578
* NET 1876 = do[1]
* NET 1879 = abc_11867_new_n1815
* NET 1882 = abc_11867_new_n1813
* NET 1883 = abc_11867_new_n1812
* NET 1886 = abc_11867_new_n1810
* NET 1890 = abc_11867_new_n1800
* NET 1897 = abc_11867_new_n1890
* NET 1898 = abc_11867_new_n1889
* NET 1901 = abc_11867_new_n1841
* NET 1902 = abc_11867_new_n1838
* NET 1907 = abc_11867_new_n1825
* NET 1910 = abc_11867_new_n1861
* NET 1911 = abc_11867_new_n1888
* NET 1914 = abc_11867_new_n1833
* NET 1915 = abc_11867_new_n1822
* NET 1916 = abc_11867_new_n1828
* NET 1917 = abc_11867_new_n1832
* NET 1922 = abc_11867_new_n1773
* NET 1923 = abc_11867_new_n1857
* NET 1924 = abc_11867_new_n1886
* NET 1926 = abc_11867_new_n1858
* NET 1928 = abc_11867_new_n1850
* NET 1931 = abc_11867_new_n1859
* NET 1937 = abc_11867_new_n1875
* NET 1945 = abc_11867_new_n1872
* NET 1946 = abc_11867_new_n1873
* NET 1951 = abc_11867_new_n1842
* NET 1952 = abc_11867_new_n1845
* NET 1954 = abc_11867_new_n983
* NET 1956 = abc_11867_new_n1681
* NET 1959 = abc_11867_new_n1678
* NET 1966 = abc_11867_new_n1662
* NET 1967 = abc_11867_new_n1661
* NET 1972 = abc_11867_new_n1436
* NET 1973 = abc_11867_new_n1441
* NET 1975 = abc_11867_new_n1435
* NET 1976 = abc_11867_new_n1437
* NET 1977 = abc_11867_new_n484
* NET 1978 = abc_11867_new_n509
* NET 1980 = abc_11867_new_n517
* NET 1988 = abc_11867_new_n613
* NET 1992 = abc_11867_new_n691
* NET 1995 = abc_11867_new_n642
* NET 1996 = abc_11867_new_n649
* NET 1997 = abc_11867_new_n519
* NET 1998 = abc_11867_new_n831
* NET 1999 = abc_11867_new_n830
* NET 2000 = abc_11867_new_n829
* NET 2008 = abc_11867_new_n580
* NET 2015 = abc_11867_new_n763
* NET 2016 = abc_11867_new_n662
* NET 2017 = abc_11867_new_n562
* NET 2020 = subckt_1656_sff1_x4.sff_s
* NET 2021 = subckt_1656_sff1_x4.sff_m
* NET 2026 = subckt_1656_sff1_x4.ckr
* NET 2028 = clk_root_tl_tl_0
* NET 2029 = subckt_1656_sff1_x4.nckr
* NET 2101 = abc_11867_new_n1769
* NET 2103 = abc_11867_new_n1814
* NET 2105 = abc_11867_new_n1891
* NET 2107 = abc_11867_new_n1893
* NET 2108 = abc_11867_new_n1898
* NET 2117 = abc_11867_new_n1887
* NET 2119 = abc_11867_new_n1835
* NET 2120 = abc_11867_new_n1837
* NET 2121 = abc_11867_new_n1791
* NET 2122 = abc_11867_new_n1834
* NET 2127 = abc_11867_new_n1798
* NET 2128 = abc_11867_new_n1885
* NET 2129 = abc_11867_new_n1881
* NET 2133 = abc_11867_new_n1878
* NET 2137 = abc_11867_new_n1863
* NET 2138 = abc_11867_new_n1867
* NET 2139 = abc_11867_new_n1869
* NET 2145 = abc_11867_new_n356
* NET 2148 = a[1]
* NET 2151 = abc_11867_new_n503
* NET 2153 = abc_11867_new_n1688
* NET 2155 = abc_11867_new_n1689
* NET 2157 = abc_11867_new_n1663
* NET 2159 = abc_11867_new_n524
* NET 2160 = abc_11867_new_n625
* NET 2161 = abc_11867_new_n565
* NET 2170 = abc_11867_new_n646
* NET 2171 = abc_11867_new_n650
* NET 2172 = abc_11867_new_n832
* NET 2173 = abc_11867_new_n824
* NET 2174 = abc_11867_new_n523
* NET 2176 = abc_11867_new_n549
* NET 2178 = abc_11867_new_n724
* NET 2179 = abc_11867_new_n730
* NET 2180 = abc_11867_new_n725
* NET 2182 = abc_11867_new_n651
* NET 2183 = abc_11867_new_n667
* NET 2185 = abc_11867_new_n737
* NET 2187 = nmi
* NET 2189 = mos6502_nmi_1
* NET 2191 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[2]
* NET 2192 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[3]
* NET 2235 = abc_11867_new_n1728
* NET 2245 = abc_11867_new_n1760
* NET 2247 = abc_11867_new_n942
* NET 2248 = abc_11867_new_n943
* NET 2251 = abc_11867_new_n935
* NET 2252 = abc_11867_new_n936
* NET 2255 = abc_11867_new_n1799
* NET 2260 = abc_11867_new_n1669
* NET 2263 = abc_11867_new_n1871
* NET 2267 = abc_11867_new_n1879
* NET 2268 = abc_11867_new_n1877
* NET 2270 = abc_11867_new_n1870
* NET 2272 = abc_11867_new_n1880
* NET 2273 = abc_11867_new_n884
* NET 2274 = abc_11867_new_n880
* NET 2277 = abc_11867_new_n1848
* NET 2281 = a[2]
* NET 2284 = abc_11867_new_n1104
* NET 2290 = subckt_1717_sff1_x4.sff_s
* NET 2293 = abc_11867_auto_rtlil_cc_2608_muxgate_11782
* NET 2297 = subckt_1717_sff1_x4.sff_m
* NET 2299 = subckt_1717_sff1_x4.ckr
* NET 2300 = subckt_1717_sff1_x4.nckr
* NET 2301 = abc_11867_new_n1442
* NET 2302 = abc_11867_new_n1429
* NET 2305 = abc_11867_new_n615
* NET 2307 = abc_11867_new_n1687
* NET 2315 = abc_11867_new_n614
* NET 2318 = abc_11867_new_n493
* NET 2320 = abc_11867_new_n1433
* NET 2321 = abc_11867_new_n1431
* NET 2325 = abc_11867_new_n1439
* NET 2328 = abc_11867_new_n1438
* NET 2334 = abc_11867_new_n530
* NET 2337 = abc_11867_new_n583
* NET 2343 = abc_11867_new_n581
* NET 2344 = abc_11867_new_n584
* NET 2346 = abc_11867_new_n607
* NET 2350 = abc_11867_new_n526
* NET 2354 = abc_11867_new_n552
* NET 2359 = abc_11867_new_n553
* NET 2362 = subckt_1626_sff1_x4.sff_s
* NET 2364 = subckt_1626_sff1_x4.sff_m
* NET 2370 = subckt_1626_sff1_x4.ckr
* NET 2371 = subckt_1626_sff1_x4.nckr
* NET 2372 = abc_11867_new_n790
* NET 2374 = abc_11867_new_n781
* NET 2376 = abc_11867_new_n816
* NET 2471 = abc_11867_new_n1766
* NET 2476 = abc_11867_new_n1761
* NET 2481 = abc_11867_new_n1725
* NET 2482 = abc_11867_new_n1765
* NET 2498 = abc_11867_new_n1774
* NET 2499 = abc_11867_new_n1751
* NET 2500 = abc_11867_new_n1750
* NET 2501 = abc_11867_new_n1747
* NET 2504 = abc_11867_new_n927
* NET 2505 = abc_11867_new_n926
* NET 2508 = abc_11867_new_n1824
* NET 2509 = abc_11867_new_n1710
* NET 2511 = abc_11867_new_n1712
* NET 2515 = abc_11867_new_n1926
* NET 2517 = abc_11867_new_n1884
* NET 2518 = abc_11867_new_n1925
* NET 2521 = subckt_1718_sff1_x4.sff_s
* NET 2524 = subckt_1718_sff1_x4.sff_m
* NET 2527 = abc_11867_auto_rtlil_cc_2608_muxgate_11784
* NET 2530 = subckt_1718_sff1_x4.ckr
* NET 2531 = subckt_1718_sff1_x4.nckr
* NET 2532 = abc_11867_new_n841
* NET 2535 = abc_11867_new_n845
* NET 2537 = abc_11867_new_n1679
* NET 2542 = abc_11867_new_n579
* NET 2548 = abc_11867_new_n958
* NET 2550 = abc_11867_new_n960
* NET 2551 = abc_11867_new_n1430
* NET 2555 = abc_11867_new_n1440
* NET 2559 = abc_11867_new_n569
* NET 2563 = abc_11867_new_n774
* NET 2564 = abc_11867_new_n777
* NET 2566 = mos6502_state[1]
* NET 2567 = abc_11867_new_n621
* NET 2569 = abc_11867_new_n620
* NET 2570 = abc_11867_new_n616
* NET 2571 = abc_11867_new_n551
* NET 2572 = abc_11867_new_n563
* NET 2573 = abc_11867_new_n809
* NET 2576 = abc_11867_new_n810
* NET 2578 = abc_11867_new_n566
* NET 2579 = abc_11867_new_n571
* NET 2582 = abc_11867_new_n668
* NET 2584 = abc_11867_new_n528
* NET 2586 = abc_11867_new_n508
* NET 2587 = abc_11867_new_n623
* NET 2588 = abc_11867_new_n820
* NET 2589 = abc_11867_new_n529
* NET 2591 = abc_11867_new_n669
* NET 2592 = abc_11867_new_n554
* NET 2593 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[0]
* NET 2596 = abc_11867_new_n815
* NET 2639 = abc_11867_new_n1763
* NET 2644 = abc_11867_new_n1767
* NET 2645 = abc_11867_new_n1762
* NET 2648 = abc_11867_new_n1756
* NET 2659 = abc_11867_new_n1738
* NET 2662 = abc_11867_new_n1785
* NET 2664 = abc_11867_new_n1759
* NET 2666 = abc_11867_new_n1784
* NET 2670 = abc_11867_new_n1783
* NET 2671 = abc_11867_new_n1786
* NET 2672 = abc_11867_new_n1789
* NET 2675 = abc_11867_new_n1788
* NET 2678 = abc_11867_new_n1780
* NET 2682 = abc_11867_new_n1782
* NET 2685 = abc_11867_new_n1787
* NET 2693 = subckt_1750_sff1_x4.sff_s
* NET 2699 = abc_11867_auto_rtlil_cc_2608_muxgate_11848
* NET 2701 = subckt_1750_sff1_x4.sff_m
* NET 2703 = subckt_1750_sff1_x4.ckr
* NET 2704 = subckt_1750_sff1_x4.nckr
* NET 2706 = abc_11867_new_n1924
* NET 2707 = abc_11867_new_n1883
* NET 2711 = abc_11867_new_n1882
* NET 2715 = abc_11867_new_n1703
* NET 2718 = abc_11867_new_n1126
* NET 2723 = abc_11867_new_n848
* NET 2727 = abc_11867_new_n956
* NET 2732 = abc_11867_new_n957
* NET 2734 = abc_11867_new_n1102
* NET 2743 = abc_11867_new_n1432
* NET 2745 = abc_11867_new_n1100
* NET 2746 = abc_11867_new_n1101
* NET 2748 = abc_11867_new_n767
* NET 2749 = abc_11867_new_n769
* NET 2754 = abc_11867_new_n850
* NET 2756 = abc_11867_new_n612
* NET 2760 = abc_11867_new_n570
* NET 2763 = abc_11867_new_n806
* NET 2764 = abc_11867_new_n653
* NET 2769 = abc_11867_new_n776
* NET 2771 = abc_11867_new_n834
* NET 2772 = abc_11867_new_n833
* NET 2773 = abc_11867_new_n835
* NET 2775 = abc_11867_new_n622
* NET 2776 = abc_11867_new_n817
* NET 2781 = abc_11867_new_n555
* NET 2782 = abc_11867_new_n573
* NET 2783 = abc_11867_new_n593
* NET 2784 = abc_11867_new_n505
* NET 2787 = abc_11867_new_n592
* NET 2789 = abc_11867_new_n634
* NET 2795 = abc_11867_new_n811
* NET 2798 = abc_11867_new_n803
* NET 2803 = abc_11867_new_n733
* NET 2805 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[1]
* NET 2847 = abc_11867_new_n807
* NET 2884 = abc_11867_new_n967
* NET 2887 = abc_11867_new_n962
* NET 2890 = abc_11867_new_n427
* NET 2897 = abc_11867_new_n837
* NET 2898 = abc_11867_new_n788
* NET 2904 = abc_11867_new_n1903
* NET 2906 = abc_11867_new_n1768
* NET 2907 = abc_11867_new_n1902
* NET 2910 = abc_11867_new_n1790
* NET 2911 = abc_11867_new_n1901
* NET 2920 = abc_11867_new_n1737
* NET 2922 = abc_11867_new_n1764
* NET 2923 = abc_11867_new_n1757
* NET 2926 = abc_11867_new_n1779
* NET 2927 = abc_11867_new_n1776
* NET 2930 = abc_11867_new_n1781
* NET 2931 = abc_11867_new_n1777
* NET 2933 = abc_11867_new_n1778
* NET 2934 = abc_11867_new_n1775
* NET 2936 = abc_11867_new_n1715
* NET 2937 = abc_11867_new_n1847
* NET 2938 = abc_11867_new_n885
* NET 2939 = do[0]
* NET 2940 = abc_11867_new_n847
* NET 2942 = abc_11867_new_n1701
* NET 2944 = abc_11867_new_n1704
* NET 2945 = abc_11867_new_n1706
* NET 2947 = abc_11867_new_n1707
* NET 2949 = abc_11867_new_n1648
* NET 2958 = abc_11867_new_n770
* NET 2960 = abc_11867_new_n487
* NET 2961 = abc_11867_new_n381
* NET 2962 = abc_11867_new_n488
* NET 2963 = abc_11867_new_n477
* NET 2964 = abc_11867_new_n853
* NET 2965 = abc_11867_new_n852
* NET 2966 = abc_11867_new_n851
* NET 2968 = abc_11867_new_n771
* NET 2972 = abc_11867_new_n778
* NET 2974 = abc_11867_new_n861
* NET 2976 = abc_11867_new_n870
* NET 2978 = abc_11867_new_n779
* NET 2979 = abc_11867_new_n772
* NET 2981 = abc_11867_new_n780
* NET 2983 = abc_11867_new_n550
* NET 2986 = mos6502_state[4]
* NET 2988 = subckt_1629_sff1_x4.sff_s
* NET 2992 = subckt_1629_sff1_x4.sff_m
* NET 2994 = subckt_1629_sff1_x4.ckr
* NET 2995 = subckt_1629_sff1_x4.nckr
* NET 2997 = abc_11867_new_n800
* NET 2998 = abc_11867_new_n556
* NET 2999 = abc_11867_new_n572
* NET 3000 = abc_11867_new_n574
* NET 3001 = abc_11867_new_n560
* NET 3005 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[5]
* NET 3006 = abc_11867_new_n632
* NET 3007 = abc_11867_new_n635
* NET 3009 = abc_11867_new_n789
* NET 3011 = abc_11867_new_n818
* NET 3012 = abc_11867_new_n819
* NET 3015 = abc_11867_new_n814
* NET 3048 = abc_11867_new_n515
* NET 3049 = abc_11867_new_n700
* NET 3055 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[4]
* NET 3058 = abc_11867_new_n808
* NET 3061 = abc_11867_new_n826
* NET 3065 = abc_11867_new_n1739
* NET 3066 = abc_11867_new_n1729
* NET 3073 = abc_11867_new_n1734
* NET 3076 = spare_buffer_74.q
* NET 3078 = abc_11867_new_n1713
* NET 3082 = abc_11867_new_n1709
* NET 3083 = abc_11867_new_n1702
* NET 3085 = abc_11867_new_n1742
* NET 3090 = abc_11867_new_n1758
* NET 3092 = abc_11867_new_n1755
* NET 3095 = abc_11867_new_n1754
* NET 3100 = abc_11867_new_n1752
* NET 3102 = abc_11867_new_n1753
* NET 3106 = abc_11867_new_n1731
* NET 3110 = abc_11867_new_n1819
* NET 3113 = spare_buffer_70.q
* NET 3120 = abc_11867_new_n961
* NET 3121 = abc_11867_new_n1045
* NET 3125 = abc_11867_new_n1044
* NET 3126 = abc_11867_new_n1041
* NET 3133 = abc_11867_new_n491
* NET 3136 = abc_11867_new_n382
* NET 3137 = abc_11867_new_n483
* NET 3141 = abc_11867_new_n1659
* NET 3144 = abc_11867_new_n959
* NET 3148 = spare_buffer_58.q
* NET 3150 = abc_11867_new_n1428
* NET 3154 = abc_11867_new_n590
* NET 3156 = abc_11867_new_n591
* NET 3158 = reset
* NET 3160 = abc_11867_new_n495
* NET 3163 = abc_11867_new_n836
* NET 3164 = abc_11867_new_n506
* NET 3165 = abc_11867_new_n655
* NET 3170 = abc_11867_new_n797
* NET 3171 = abc_11867_new_n798
* NET 3172 = spare_buffer_54.q
* NET 3175 = abc_11867_new_n827
* NET 3178 = abc_11867_new_n731
* NET 3180 = abc_11867_new_n732
* NET 3181 = abc_11867_new_n792
* NET 3246 = abc_11867_new_n1743
* NET 3247 = abc_11867_new_n1744
* NET 3251 = spare_buffer_73.q
* NET 3254 = abc_11867_new_n1682
* NET 3257 = abc_11867_new_n1683
* NET 3258 = abc_11867_new_n1696
* NET 3261 = abc_11867_new_n1649
* NET 3262 = abc_11867_new_n1862
* NET 3265 = abc_11867_new_n1014
* NET 3266 = abc_11867_new_n1771
* NET 3269 = abc_11867_new_n1823
* NET 3271 = abc_11867_new_n1866
* NET 3273 = abc_11867_new_n1820
* NET 3274 = abc_11867_new_n955
* NET 3275 = abc_11867_new_n1868
* NET 3276 = spare_buffer_69.q
* NET 3278 = clk_root_tr_0
* NET 3280 = abc_11867_new_n1046
* NET 3281 = a[8]
* NET 3285 = abc_11867_new_n952
* NET 3288 = abc_11867_new_n950
* NET 3289 = abc_11867_new_n972
* NET 3290 = abc_11867_new_n1042
* NET 3291 = abc_11867_new_n1039
* NET 3294 = abc_11867_new_n575
* NET 3295 = abc_11867_new_n499
* NET 3297 = abc_11867_new_n486
* NET 3300 = abc_11867_new_n520
* NET 3302 = spare_buffer_57.q
* NET 3305 = abc_11867_new_n701
* NET 3307 = abc_11867_new_n489
* NET 3310 = abc_11867_new_n511
* NET 3314 = abc_11867_new_n504
* NET 3315 = abc_11867_new_n510
* NET 3317 = abc_11867_new_n597
* NET 3318 = abc_11867_new_n711
* NET 3320 = abc_11867_new_n428_hfns_5
* NET 3324 = abc_11867_new_n513
* NET 3325 = abc_11867_new_n512
* NET 3326 = abc_11867_new_n561
* NET 3327 = spare_buffer_53.q
* NET 3329 = clk_root_tl_bl_0
* NET 3330 = clk_root_tl_0
* NET 3333 = abc_11867_new_n426_hfns_1
* NET 3334 = abc_11867_new_n739
* NET 3335 = abc_11867_new_n762
* NET 3338 = abc_11867_new_n716
* NET 3341 = abc_11867_new_n802
* NET 3342 = abc_11867_new_n813
* NET 3343 = abc_11867_new_n812
* NET 3388 = abc_11867_new_n1912
* NET 3389 = abc_11867_new_n1723
* NET 3390 = abc_11867_new_n1909
* NET 3392 = abc_11867_new_n1911
* NET 3395 = abc_11867_new_n1717
* NET 3396 = abc_11867_new_n1724
* NET 3398 = abc_11867_new_n1718
* NET 3400 = abc_11867_new_n1692
* NET 3405 = abc_11867_new_n1697
* NET 3411 = abc_11867_new_n1699
* NET 3414 = abc_11867_new_n1650
* NET 3415 = abc_11867_new_n1698
* NET 3429 = abc_11867_new_n1686
* NET 3433 = abc_11867_new_n1772
* NET 3441 = a[0]
* NET 3445 = abc_11867_new_n1865
* NET 3448 = subckt_1724_sff1_x4.sff_s
* NET 3452 = abc_11867_auto_rtlil_cc_2608_muxgate_11796
* NET 3455 = subckt_1724_sff1_x4.sff_m
* NET 3458 = subckt_1724_sff1_x4.ckr
* NET 3459 = subckt_1724_sff1_x4.nckr
* NET 3460 = abc_11867_new_n954
* NET 3462 = abc_11867_new_n953
* NET 3463 = abc_11867_new_n949
* NET 3467 = abc_11867_new_n968
* NET 3469 = abc_11867_new_n918
* NET 3471 = abc_11867_new_n846
* NET 3472 = abc_11867_new_n849
* NET 3478 = abc_11867_new_n1705
* NET 3479 = abc_11867_new_n1708
* NET 3482 = abc_11867_new_n1666
* NET 3484 = abc_11867_new_n1664
* NET 3485 = abc_11867_new_n1660
* NET 3490 = abc_11867_new_n473_hfns_2
* NET 3493 = abc_11867_new_n637
* NET 3494 = abc_11867_new_n643
* NET 3498 = abc_11867_new_n740
* NET 3502 = abc_11867_new_n588
* NET 3509 = abc_11867_new_n773
* NET 3512 = abc_11867_new_n709
* NET 3516 = abc_11867_new_n596
* NET 3519 = abc_11867_new_n713
* NET 3525 = abc_11867_new_n715
* NET 3526 = abc_11867_new_n714
* NET 3527 = abc_11867_new_n702
* NET 3531 = abc_11867_new_n471_hfns_0
* NET 3535 = abc_11867_new_n839
* NET 3538 = abc_11867_new_n787
* NET 3539 = abc_11867_new_n838
* NET 3541 = abc_11867_new_n786
* NET 3544 = abc_11867_new_n694
* NET 3546 = abc_11867_new_n720
* NET 3547 = abc_11867_new_n717
* NET 3551 = abc_11867_new_n683
* NET 3552 = abc_11867_new_n801
* NET 3553 = abc_11867_new_n799
* NET 3637 = abc_11867_new_n1665
* NET 3639 = abc_11867_new_n1900
* NET 3641 = abc_11867_new_n1905
* NET 3644 = abc_11867_new_n1740
* NET 3646 = abc_11867_new_n1741
* NET 3648 = abc_11867_new_n1745
* NET 3650 = abc_11867_new_n1920
* NET 3651 = abc_11867_new_n1913
* NET 3652 = abc_11867_new_n1897
* NET 3654 = abc_11867_new_n1716
* NET 3655 = abc_11867_new_n1711
* NET 3657 = abc_11867_new_n1714
* NET 3658 = abc_11867_new_n1693
* NET 3660 = abc_11867_new_n1676
* NET 3662 = abc_11867_new_n1735
* NET 3665 = abc_11867_new_n1736
* NET 3666 = abc_11867_new_n1732
* NET 3668 = abc_11867_new_n1733
* NET 3670 = abc_11867_new_n1695
* NET 3671 = abc_11867_new_n1694
* NET 3672 = abc_11867_new_n1685
* NET 3673 = abc_11867_new_n1680
* NET 3676 = abc_11867_new_n1691
* NET 3677 = abc_11867_new_n1690
* NET 3678 = abc_11867_new_n1416
* NET 3680 = abc_11867_new_n1118
* NET 3685 = abc_11867_new_n1730
* NET 3688 = subckt_1716_sff1_x4.sff_s
* NET 3691 = subckt_1716_sff1_x4.sff_m
* NET 3693 = abc_11867_auto_rtlil_cc_2608_muxgate_11780
* NET 3695 = subckt_1716_sff1_x4.ckr
* NET 3696 = subckt_1716_sff1_x4.nckr
* NET 3698 = subckt_1720_sff1_x4.sff_s
* NET 3703 = subckt_1720_sff1_x4.sff_m
* NET 3705 = clk_root_tr_bl_0
* NET 3706 = subckt_1720_sff1_x4.ckr
* NET 3707 = subckt_1720_sff1_x4.nckr
* NET 3709 = abc_11867_new_n1110
* NET 3716 = abc_11867_new_n647
* NET 3717 = abc_11867_new_n609
* NET 3718 = abc_11867_new_n924
* NET 3721 = abc_11867_new_n923
* NET 3723 = abc_11867_new_n1043
* NET 3730 = subckt_1715_sff1_x4.sff_s
* NET 3733 = subckt_1715_sff1_x4.sff_m
* NET 3735 = abc_11867_auto_rtlil_cc_2608_muxgate_11778
* NET 3736 = subckt_1715_sff1_x4.ckr
* NET 3738 = subckt_1715_sff1_x4.nckr
* NET 3744 = abc_11867_new_n474
* NET 3745 = abc_11867_new_n636
* NET 3749 = abc_11867_new_n589
* NET 3750 = mos6502_backwards
* NET 3753 = abc_11867_new_n475_hfns_1
* NET 3755 = abc_11867_new_n1175
* NET 3759 = abc_11867_new_n502
* NET 3761 = abc_11867_new_n712
* NET 3762 = abc_11867_new_n710
* NET 3763 = abc_11867_new_n703
* NET 3765 = abc_11867_new_n785
* NET 3767 = abc_11867_new_n475_hfns_2
* NET 3771 = abc_11867_new_n704
* NET 3772 = abc_11867_new_n822
* NET 3773 = abc_11867_new_n796
* NET 3775 = abc_11867_new_n794
* NET 3776 = abc_11867_new_n795
* NET 3809 = abc_11867_new_n1931
* NET 3811 = abc_11867_new_n1933
* NET 3812 = abc_11867_new_n1932
* NET 3814 = abc_11867_new_n1908
* NET 3822 = abc_11867_new_n1906
* NET 3824 = abc_11867_new_n1910
* NET 3825 = abc_11867_new_n1907
* NET 3826 = abc_11867_new_n1904
* NET 3827 = abc_11867_new_n1746
* NET 3828 = abc_11867_new_n1720
* NET 3832 = abc_11867_new_n1700
* NET 3835 = abc_11867_new_n1914
* NET 3838 = abc_11867_new_n1670
* NET 3840 = abc_11867_new_n999
* NET 3843 = abc_11867_new_n1124
* NET 3846 = abc_11867_new_n1022
* NET 3849 = abc_11867_new_n1132
* NET 3854 = abc_11867_new_n1794
* NET 3857 = abc_11867_new_n1795
* NET 3860 = abc_11867_new_n353
* NET 3861 = abc_11867_new_n954_hfns_2
* NET 3863 = abc_11867_auto_rtlil_cc_2608_muxgate_11788
* NET 3866 = a[4]
* NET 3872 = abc_11867_new_n928
* NET 3874 = abc_11867_new_n933
* NET 3875 = abc_11867_new_n931
* NET 3880 = abc_11867_new_n932
* NET 3881 = abc_11867_new_n930
* NET 3884 = abc_11867_new_n921
* NET 3885 = abc_11867_new_n843
* NET 3897 = abc_11867_new_n727
* NET 3898 = abc_11867_new_n482_hfns_1
* NET 3903 = abc_11867_new_n974
* NET 3912 = abc_11867_new_n624
* NET 3915 = abc_11867_new_n564
* NET 3920 = subckt_1655_sff1_x4.sff_s
* NET 3925 = subckt_1655_sff1_x4.sff_m
* NET 3927 = abc_11867_auto_rtlil_cc_2608_muxgate_11670
* NET 3929 = subckt_1655_sff1_x4.ckr
* NET 3930 = subckt_1655_sff1_x4.nckr
* NET 3931 = abc_11867_new_n498
* NET 3936 = abc_11867_new_n501
* NET 3942 = abc_11867_new_n568
* NET 3944 = abc_11867_new_n594
* NET 3946 = abc_11867_new_n492
* NET 3950 = abc_11867_new_n783
* NET 3956 = abc_11867_new_n473_hfns_0
* NET 3960 = abc_11867_new_n514_hfns_1
* NET 3964 = abc_11867_new_n471_hfns_1
* NET 3968 = abc_11867_new_n693
* NET 3969 = abc_11867_new_n692
* NET 3972 = abc_11867_new_n684
* NET 3973 = abc_11867_new_n686
* NET 3977 = abc_11867_new_n679
* NET 3978 = abc_11867_new_n671
* NET 3979 = abc_11867_new_n678
* NET 4027 = abc_11867_new_n765
* NET 4040 = abc_11867_new_n352
* NET 4046 = abc_11867_new_n386
* NET 4049 = subckt_1754_sff1_x4.sff_s
* NET 4050 = subckt_1754_sff1_x4.ckr
* NET 4053 = subckt_1754_sff1_x4.sff_m
* NET 4055 = abc_11867_auto_rtlil_cc_2608_muxgate_11856
* NET 4057 = clk_root_tr_br_0
* NET 4058 = subckt_1754_sff1_x4.nckr
* NET 4059 = abc_11867_new_n1921
* NET 4061 = abc_11867_new_n1922
* NET 4062 = abc_11867_new_n1919
* NET 4064 = abc_11867_new_n1894
* NET 4065 = abc_11867_new_n1918
* NET 4068 = abc_11867_new_n1140
* NET 4073 = abc_11867_new_n1146
* NET 4075 = abc_11867_new_n610
* NET 4079 = abc_11867_new_n1030
* NET 4083 = a[7]
* NET 4085 = abc_11867_new_n1015
* NET 4087 = abc_11867_new_n1020
* NET 4088 = abc_11867_new_n981
* NET 4090 = abc_11867_new_n976
* NET 4092 = abc_11867_new_n1012
* NET 4095 = abc_11867_new_n1007
* NET 4096 = abc_11867_new_n1864
* NET 4099 = abc_11867_new_n1040
* NET 4103 = abc_11867_new_n922
* NET 4105 = abc_11867_new_n929
* NET 4108 = abc_11867_new_n887
* NET 4109 = abc_11867_new_n482_hfns_0
* NET 4111 = abc_11867_new_n608_hfns_1
* NET 4114 = subckt_1699_sff1_x4.sff_s
* NET 4115 = subckt_1699_sff1_x4.ckr
* NET 4118 = subckt_1699_sff1_x4.sff_m
* NET 4121 = clk_root_tl_br_0
* NET 4122 = subckt_1699_sff1_x4.nckr
* NET 4123 = abc_11867_auto_rtlil_cc_2608_muxgate_11746
* NET 4126 = abc_11867_new_n1338
* NET 4127 = abc_11867_new_n1337
* NET 4132 = abc_11867_new_n496
* NET 4135 = abc_11867_new_n494
* NET 4138 = abc_11867_new_n869
* NET 4139 = abc_11867_new_n426_hfns_0
* NET 4140 = abc_11867_new_n784
* NET 4142 = abc_11867_new_n497
* NET 4143 = abc_11867_new_n630
* NET 4144 = abc_11867_new_n626
* NET 4147 = abc_11867_new_n531
* NET 4148 = abc_11867_new_n548
* NET 4152 = abc_11867_new_n699
* NET 4153 = abc_11867_new_n682
* NET 4154 = abc_11867_new_n680
* NET 4157 = abc_11867_new_n533
* NET 4158 = rdy
* NET 4205 = subckt_1749_sff1_x4.sff_m
* NET 4206 = abc_11867_auto_rtlil_cc_2608_muxgate_11846
* NET 4210 = subckt_1758_sff1_x4.sff_m
* NET 4213 = subckt_1723_sff1_x4.sff_m
* NET 4215 = abc_11867_auto_rtlil_cc_2608_muxgate_11794
* NET 4217 = abc_11867_new_n1339
* NET 4225 = subckt_1685_sff1_x4.sff_m
* NET 4229 = subckt_1686_sff1_x4.sff_m
* NET 4230 = abc_11867_new_n805
* NET 4235 = subckt_1684_sff1_x4.sff_m
* NET 4237 = abc_11867_new_n793
* NET 4238 = subckt_1749_sff1_x4.sff_s
* NET 4243 = subckt_1749_sff1_x4.ckr
* NET 4244 = subckt_1749_sff1_x4.nckr
* NET 4247 = abc_11867_new_n1916
* NET 4250 = subckt_1758_sff1_x4.sff_s
* NET 4255 = subckt_1758_sff1_x4.ckr
* NET 4256 = subckt_1758_sff1_x4.nckr
* NET 4258 = abc_11867_new_n1895
* NET 4268 = subckt_1723_sff1_x4.sff_s
* NET 4275 = subckt_1723_sff1_x4.ckr
* NET 4276 = subckt_1723_sff1_x4.nckr
* NET 4279 = abc_11867_new_n1116
* NET 4281 = abc_11867_new_n1117
* NET 4285 = abc_11867_new_n1038
* NET 4286 = abc_11867_new_n891
* NET 4289 = abc_11867_new_n348
* NET 4292 = abc_11867_new_n1469
* NET 4295 = abc_11867_new_n1551
* NET 4299 = abc_11867_new_n968_hfns_2
* NET 4300 = abc_11867_new_n428_hfns_0
* NET 4302 = abc_11867_new_n1552
* NET 4305 = di[7]
* NET 4306 = subckt_101_nmx2_x1.q
* NET 4311 = clk
* NET 4313 = abc_11867_new_n920
* NET 4318 = abc_11867_new_n919
* NET 4319 = abc_11867_new_n357
* NET 4320 = abc_11867_new_n1464
* NET 4321 = abc_11867_new_n1461
* NET 4324 = abc_11867_new_n1654
* NET 4327 = abc_11867_new_n1647
* NET 4328 = abc_11867_new_n1653
* NET 4330 = abc_11867_new_n1658
* NET 4334 = abc_11867_new_n1652
* NET 4338 = abc_11867_new_n1393
* NET 4339 = abc_11867_new_n1400
* NET 4342 = abc_11867_new_n1394
* NET 4346 = abc_11867_new_n866
* NET 4349 = subckt_1685_sff1_x4.sff_s
* NET 4350 = mos6502_src_reg[0]
* NET 4355 = subckt_1685_sff1_x4.ckr
* NET 4356 = subckt_1685_sff1_x4.nckr
* NET 4357 = subckt_1686_sff1_x4.sff_s
* NET 4358 = mos6502_src_reg[1]
* NET 4362 = subckt_1686_sff1_x4.ckr
* NET 4364 = subckt_1686_sff1_x4.nckr
* NET 4367 = subckt_1684_sff1_x4.sff_s
* NET 4371 = subckt_1684_sff1_x4.ckr
* NET 4373 = subckt_1684_sff1_x4.nckr
* NET 4374 = rdy_hfns_4
* NET 4459 = subckt_1755_sff1_x4.sff_s
* NET 4462 = subckt_1755_sff1_x4.sff_m
* NET 4464 = abc_11867_auto_rtlil_cc_2608_muxgate_11858
* NET 4466 = subckt_1755_sff1_x4.ckr
* NET 4467 = subckt_1755_sff1_x4.nckr
* NET 4469 = abc_11867_new_n1899
* NET 4471 = abc_11867_auto_rtlil_cc_2608_muxgate_11864
* NET 4472 = subckt_1615_nmx2_x1.q
* NET 4473 = abc_11867_new_n336
* NET 4476 = abc_11867_new_n1121
* NET 4479 = abc_11867_new_n1120
* NET 4481 = abc_11867_new_n1123
* NET 4483 = abc_11867_new_n1122
* NET 4485 = abc_11867_new_n1115
* NET 4487 = abc_11867_new_n1113
* NET 4488 = abc_11867_new_n1112
* NET 4490 = a[6]
* NET 4498 = abc_11867_new_n1108
* NET 4499 = abc_11867_new_n1106
* NET 4501 = mos6502_abl[0]
* NET 4502 = abc_11867_new_n333
* NET 4503 = abc_11867_new_n1481
* NET 4508 = subckt_1732_sff1_x4.sff_s
* NET 4511 = subckt_1732_sff1_x4.sff_m
* NET 4514 = subckt_1732_sff1_x4.ckr
* NET 4515 = subckt_1732_sff1_x4.nckr
* NET 4516 = abc_11867_auto_rtlil_cc_2608_muxgate_11812
* NET 4518 = abc_11867_new_n1470
* NET 4519 = abc_11867_new_n1483
* NET 4520 = abc_11867_new_n1482
* NET 4522 = mos6502_abh[0]
* NET 4523 = abc_11867_new_n1553
* NET 4526 = abc_11867_new_n1109
* NET 4527 = abc_11867_new_n1107
* NET 4529 = abc_11867_new_n648
* NET 4530 = abc_11867_new_n611
* NET 4532 = abc_11867_new_n631
* NET 4533 = abc_11867_new_n595
* NET 4536 = abc_11867_new_n608_hfns_0
* NET 4538 = abc_11867_new_n888
* NET 4539 = abc_11867_new_n1497
* NET 4541 = abc_11867_new_n619
* NET 4545 = subckt_1689_sff1_x4.sff_s
* NET 4548 = subckt_1689_sff1_x4.sff_m
* NET 4550 = subckt_1689_sff1_x4.ckr
* NET 4552 = subckt_1689_sff1_x4.nckr
* NET 4553 = abc_11867_new_n331
* NET 4554 = abc_11867_auto_rtlil_cc_2608_muxgate_11740
* NET 4557 = abc_11867_new_n363
* NET 4558 = abc_11867_new_n324
* NET 4562 = abc_11867_new_n1401
* NET 4563 = abc_11867_new_n328
* NET 4564 = abc_11867_new_n1398
* NET 4565 = abc_11867_new_n1366
* NET 4567 = subckt_1709_sff1_x4.sff_s
* NET 4572 = subckt_1709_sff1_x4.sff_m
* NET 4573 = abc_11867_auto_rtlil_cc_2608_muxgate_11768
* NET 4575 = subckt_1709_sff1_x4.ckr
* NET 4576 = subckt_1709_sff1_x4.nckr
* NET 4577 = abc_11867_new_n475_hfns_0
* NET 4579 = abc_11867_new_n1181
* NET 4580 = abc_11867_new_n387
* NET 4583 = mos6502_index_y
* NET 4584 = abc_11867_auto_rtlil_cc_2608_muxgate_11728
* NET 4590 = subckt_1687_sff1_x4.sff_s
* NET 4593 = subckt_1687_sff1_x4.sff_m
* NET 4597 = subckt_1687_sff1_x4.nckr
* NET 4598 = subckt_1687_sff1_x4.ckr
* NET 4646 = abc_11867_new_n1722
* NET 4650 = subckt_1752_sff1_x4.sff_s
* NET 4652 = subckt_1752_sff1_x4.sff_m
* NET 4658 = subckt_1752_sff1_x4.ckr
* NET 4659 = subckt_1752_sff1_x4.nckr
* NET 4660 = abc_11867_auto_rtlil_cc_2608_muxgate_11852
* NET 4662 = abc_11867_new_n1896
* NET 4667 = subckt_1751_sff1_x4.sff_s
* NET 4670 = subckt_1751_sff1_x4.sff_m
* NET 4673 = abc_11867_auto_rtlil_cc_2608_muxgate_11850
* NET 4676 = subckt_1751_sff1_x4.ckr
* NET 4677 = subckt_1751_sff1_x4.nckr
* NET 4679 = subckt_1722_sff1_x4.sff_s
* NET 4682 = subckt_1722_sff1_x4.sff_m
* NET 4683 = abc_11867_auto_rtlil_cc_2608_muxgate_11792
* NET 4688 = subckt_1722_sff1_x4.ckr
* NET 4689 = subckt_1722_sff1_x4.nckr
* NET 4690 = abc_11867_new_n1036
* NET 4693 = abc_11867_new_n1675
* NET 4697 = abc_11867_new_n423
* NET 4700 = abc_11867_new_n905
* NET 4703 = abc_11867_new_n980
* NET 4706 = abc_11867_new_n1460
* NET 4712 = abc_11867_new_n890
* NET 4714 = abc_11867_new_n1480
* NET 4715 = mos6502_pc[0]
* NET 4718 = abc_11867_new_n1485
* NET 4720 = abc_11867_new_n1498
* NET 4723 = abc_11867_new_n422
* NET 4727 = mos6502_dihold[7]
* NET 4728 = subckt_1697_sff1_x4.sff_s
* NET 4731 = subckt_1697_sff1_x4.sff_m
* NET 4735 = subckt_1697_sff1_x4.ckr
* NET 4737 = subckt_1697_sff1_x4.nckr
* NET 4744 = abc_11867_new_n903
* NET 4747 = mos6502_nmi_edge
* NET 4748 = abc_11867_new_n1488
* NET 4750 = abc_11867_new_n728
* NET 4751 = irq
* NET 4754 = mos6502_i
* NET 4755 = abc_11867_new_n434
* NET 4758 = mos6502_res
* NET 4759 = abc_11867_new_n323
* NET 4768 = abc_11867_new_n1099
* NET 4773 = abc_11867_new_n1657
* NET 4776 = subckt_1713_sff1_x4.sff_s
* NET 4778 = abc_11867_auto_rtlil_cc_2608_muxgate_11776
* NET 4781 = subckt_1713_sff1_x4.sff_m
* NET 4785 = subckt_1713_sff1_x4.ckr
* NET 4786 = subckt_1713_sff1_x4.nckr
* NET 4787 = abc_11867_new_n1392
* NET 4788 = abc_11867_new_n1399
* NET 4789 = abc_11867_new_n1404
* NET 4791 = abc_11867_new_n1368
* NET 4792 = abc_11867_new_n617
* NET 4795 = abc_11867_new_n1651
* NET 4799 = abc_11867_new_n347
* NET 4801 = subckt_1682_sff1_x4.sff_s
* NET 4805 = subckt_1682_sff1_x4.sff_m
* NET 4809 = subckt_1682_sff1_x4.nckr
* NET 4810 = subckt_1682_sff1_x4.ckr
* NET 4811 = subckt_1661_sff1_x4.sff_s
* NET 4816 = subckt_1661_sff1_x4.sff_m
* NET 4820 = subckt_1661_sff1_x4.ckr
* NET 4821 = subckt_1661_sff1_x4.nckr
* NET 4822 = abc_11867_new_n1300
* NET 4823 = abc_11867_auto_rtlil_cc_2608_muxgate_11732
* NET 4826 = abc_11867_new_n688
* NET 4830 = abc_11867_new_n1181_hfns_2
* NET 4832 = abc_11867_auto_rtlil_cc_2608_muxgate_11734
* NET 4833 = mos6502_dst_reg[0]
* NET 4839 = abc_11867_new_n723
* NET 4927 = abc_11867_new_n1143
* NET 4928 = abc_11867_new_n341
* NET 4929 = abc_11867_new_n335
* NET 4934 = abc_11867_new_n1142
* NET 4935 = abc_11867_new_n1145
* NET 4937 = abc_11867_new_n1144
* NET 4941 = abc_11867_new_n1139
* NET 4943 = mos6502_alu_hc
* NET 4944 = abc_11867_new_n1114
* NET 4947 = abc_11867_new_n1131
* NET 4949 = abc_11867_new_n1035
* NET 4951 = abc_11867_new_n1033
* NET 4952 = abc_11867_new_n1034
* NET 4955 = abc_11867_new_n1031
* NET 4957 = abc_11867_new_n355
* NET 4961 = abc_11867_new_n979
* NET 4963 = abc_11867_new_n368
* NET 4965 = abc_11867_new_n1674
* NET 4966 = abc_11867_new_n1673
* NET 4968 = abc_11867_new_n997
* NET 4971 = abc_11867_new_n977
* NET 4973 = abc_11867_new_n1500
* NET 4974 = abc_11867_new_n1499
* NET 4977 = mos6502_abl[2]
* NET 4978 = abc_11867_new_n1496
* NET 4979 = abc_11867_new_n989
* NET 4984 = abc_11867_new_n587
* NET 4985 = abc_11867_new_n1471
* NET 4986 = abc_11867_new_n577
* NET 4987 = abc_11867_new_n1474
* NET 4988 = abc_11867_new_n585
* NET 4990 = abc_11867_new_n1489
* NET 4997 = abc_11867_new_n1377
* NET 4999 = abc_11867_new_n481
* NET 5002 = subckt_1677_sff1_x4.sff_s
* NET 5005 = subckt_1677_sff1_x4.sff_m
* NET 5007 = subckt_1677_sff1_x4.ckr
* NET 5009 = subckt_1677_sff1_x4.nckr
* NET 5010 = abc_11867_new_n969
* NET 5011 = abc_11867_new_n1098
* NET 5013 = abc_11867_new_n473_hfns_1
* NET 5014 = abc_11867_new_n1655
* NET 5015 = abc_11867_new_n1403
* NET 5023 = abc_11867_new_n1367
* NET 5031 = abc_11867_new_n1365
* NET 5033 = abc_11867_new_n385
* NET 5035 = abc_11867_auto_rtlil_cc_2608_muxgate_11724
* NET 5036 = mos6502_write_back
* NET 5041 = abc_11867_new_n1363
* NET 5042 = abc_11867_new_n344
* NET 5043 = abc_11867_new_n764
* NET 5044 = abc_11867_new_n782
* NET 5046 = abc_11867_new_n514_hfns_0
* NET 5048 = abc_11867_new_n384
* NET 5050 = subckt_1666_sff1_x4.sff_s
* NET 5053 = subckt_1666_sff1_x4.sff_m
* NET 5057 = subckt_1666_sff1_x4.ckr
* NET 5058 = subckt_1666_sff1_x4.nckr
* NET 5059 = abc_11867_new_n719
* NET 5112 = abc_11867_new_n1917
* NET 5119 = abc_11867_new_n1136
* NET 5124 = abc_11867_new_n1138
* NET 5127 = abc_11867_new_n1134
* NET 5130 = abc_11867_new_n1130
* NET 5137 = abc_11867_new_n1129
* NET 5139 = abc_11867_new_n1128
* NET 5142 = abc_11867_new_n1032
* NET 5143 = abc_11867_new_n375
* NET 5146 = a[5]
* NET 5150 = abc_11867_new_n1727
* NET 5153 = abc_11867_new_n996
* NET 5160 = abc_11867_new_n904
* NET 5161 = abc_11867_new_n992
* NET 5162 = abc_11867_new_n350
* NET 5166 = abc_11867_new_n1484
* NET 5169 = abc_11867_new_n1478
* NET 5170 = abc_11867_new_n1490
* NET 5171 = abc_11867_new_n1491
* NET 5173 = abc_11867_new_n984
* NET 5174 = abc_11867_new_n349
* NET 5176 = abc_11867_new_n1554
* NET 5179 = abc_11867_new_n988
* NET 5180 = abc_11867_new_n985
* NET 5183 = abc_11867_new_n1844
* NET 5186 = abc_11867_new_n944
* NET 5188 = mos6502_abl[1]
* NET 5189 = abc_11867_new_n947
* NET 5192 = abc_11867_new_n471_hfns_2
* NET 5196 = abc_11867_new_n945
* NET 5198 = subckt_1711_sff1_x4.sff_s
* NET 5205 = subckt_1711_sff1_x4.sff_m
* NET 5207 = subckt_1711_sff1_x4.ckr
* NET 5208 = subckt_1711_sff1_x4.nckr
* NET 5209 = abc_11867_new_n1351
* NET 5212 = abc_11867_new_n1378
* NET 5214 = abc_11867_new_n879
* NET 5215 = abc_11867_new_n1375
* NET 5216 = abc_11867_new_n1379
* NET 5218 = abc_11867_new_n1376
* NET 5220 = mos6502_op[2]
* NET 5221 = subckt_1672_sff1_x4.sff_s
* NET 5228 = subckt_1672_sff1_x4.sff_m
* NET 5229 = subckt_1672_sff1_x4.ckr
* NET 5231 = abc_11867_new_n329
* NET 5232 = subckt_1672_sff1_x4.nckr
* NET 5237 = abc_11867_new_n1402
* NET 5243 = abc_11867_new_n1364
* NET 5244 = abc_11867_new_n1397
* NET 5245 = subckt_1041_nmx2_x1.q
* NET 5246 = abc_11867_new_n1395
* NET 5250 = subckt_1674_sff1_x4.sff_s
* NET 5255 = subckt_1674_sff1_x4.sff_m
* NET 5258 = subckt_1674_sff1_x4.ckr
* NET 5259 = subckt_1674_sff1_x4.nckr
* NET 5260 = abc_11867_new_n1298
* NET 5261 = abc_11867_auto_rtlil_cc_2608_muxgate_11730
* NET 5263 = mos6502_php
* NET 5265 = abc_11867_new_n1185
* NET 5267 = abc_11867_auto_rtlil_cc_2608_muxgate_11680
* NET 5269 = abc_11867_new_n757
* NET 5270 = mos6502_cli
* NET 5272 = abc_11867_new_n1204
* NET 5274 = abc_11867_auto_rtlil_cc_2608_muxgate_11690
* NET 5275 = abc_11867_new_n1207
* NET 5279 = abc_11867_new_n633
* NET 5280 = abc_11867_new_n532
* NET 5284 = mos6502_sei
* NET 5285 = subckt_1667_sff1_x4.sff_s
* NET 5290 = subckt_1667_sff1_x4.sff_m
* NET 5292 = abc_11867_auto_rtlil_cc_2608_muxgate_11692
* NET 5294 = subckt_1667_sff1_x4.ckr
* NET 5295 = subckt_1667_sff1_x4.nckr
* NET 5341 = do[7]
* NET 5363 = abc_11867_new_n376
* NET 5365 = abc_11867_new_n325
* NET 5371 = abc_11867_new_n1915
* NET 5377 = subckt_1756_sff1_x4.sff_s
* NET 5378 = subckt_1756_sff1_x4.ckr
* NET 5381 = subckt_1756_sff1_x4.sff_m
* NET 5383 = abc_11867_auto_rtlil_cc_2608_muxgate_11860
* NET 5385 = subckt_1756_sff1_x4.nckr
* NET 5386 = spare_buffer_50.q
* NET 5388 = abc_11867_new_n1005
* NET 5390 = abc_11867_new_n1028
* NET 5396 = subckt_1721_sff1_x4.sff_s
* NET 5398 = subckt_1721_sff1_x4.ckr
* NET 5400 = subckt_1721_sff1_x4.sff_m
* NET 5402 = abc_11867_auto_rtlil_cc_2608_muxgate_11790
* NET 5405 = subckt_1721_sff1_x4.nckr
* NET 5406 = abc_11867_new_n1749
* NET 5408 = abc_11867_new_n1671
* NET 5411 = abc_11867_new_n993
* NET 5412 = abc_11867_new_n912
* NET 5415 = mos6502_adj_bcd
* NET 5416 = subckt_1714_sff1_x4.sff_s
* NET 5418 = subckt_1714_sff1_x4.ckr
* NET 5420 = subckt_1714_sff1_x4.sff_m
* NET 5424 = subckt_1714_sff1_x4.nckr
* NET 5426 = abc_11867_new_n1555
* NET 5427 = abc_11867_new_n1493
* NET 5428 = abc_11867_new_n359
* NET 5430 = spare_buffer_46.q
* NET 5432 = abc_11867_new_n1550
* NET 5434 = abc_11867_new_n987
* NET 5436 = abc_11867_new_n369
* NET 5438 = abc_11867_new_n1476
* NET 5440 = mos6502_alu_out[0]
* NET 5445 = abc_11867_new_n910
* NET 5446 = abc_11867_new_n432
* NET 5450 = subckt_1712_sff1_x4.sff_s
* NET 5453 = subckt_1712_sff1_x4.ckr
* NET 5455 = subckt_1712_sff1_x4.sff_m
* NET 5456 = subckt_1712_sff1_x4.nckr
* NET 5459 = abc_11867_auto_rtlil_cc_2608_muxgate_11772
* NET 5460 = abc_11867_new_n1381
* NET 5461 = abc_11867_new_n1380
* NET 5465 = abc_11867_new_n431_hfns_1
* NET 5466 = mos6502_adc_bcd
* NET 5467 = spare_buffer_34.q
* NET 5469 = abc_11867_new_n1264
* NET 5470 = mos6502_state[3]
* NET 5471 = abc_11867_new_n430_hfns_0
* NET 5474 = subckt_1675_sff1_x4.sff_s
* NET 5476 = subckt_1675_sff1_x4.ckr
* NET 5478 = subckt_1675_sff1_x4.sff_m
* NET 5482 = subckt_1675_sff1_x4.nckr
* NET 5484 = abc_11867_new_n1396
* NET 5488 = subckt_1662_sff1_x4.sff_s
* NET 5489 = subckt_1662_sff1_x4.ckr
* NET 5493 = subckt_1662_sff1_x4.sff_m
* NET 5495 = subckt_1662_sff1_x4.nckr
* NET 5496 = abc_11867_auto_rtlil_cc_2608_muxgate_11706
* NET 5498 = mos6502_rotate
* NET 5505 = abc_11867_new_n1205
* NET 5506 = spare_buffer_30.q
* NET 5508 = abc_11867_new_n697
* NET 5510 = abc_11867_new_n761
* NET 5542 = subckt_1757_sff1_x4.sff_m
* NET 5543 = abc_11867_auto_rtlil_cc_2608_muxgate_11862
* NET 5547 = subckt_1719_sff1_x4.sff_m
* NET 5548 = abc_11867_new_n1487
* NET 5551 = abc_11867_new_n937
* NET 5554 = abc_11867_new_n1265
* NET 5555 = abc_11867_auto_rtlil_cc_2608_muxgate_11714
* NET 5557 = abc_11867_new_n1463
* NET 5562 = abc_11867_new_n431_hfns_0
* NET 5563 = abc_11867_new_n430_hfns_1
* NET 5565 = mos6502_clc
* NET 5569 = subckt_1663_sff1_x4.sff_m
* NET 5572 = subckt_1757_sff1_x4.sff_s
* NET 5577 = subckt_1757_sff1_x4.ckr
* NET 5578 = subckt_1757_sff1_x4.nckr
* NET 5580 = abc_11867_new_n1677
* NET 5586 = abc_11867_new_n1137
* NET 5587 = abc_11867_new_n1135
* NET 5590 = spare_buffer_49.q
* NET 5593 = subckt_1719_sff1_x4.sff_s
* NET 5598 = subckt_1719_sff1_x4.ckr
* NET 5599 = subckt_1719_sff1_x4.nckr
* NET 5600 = abc_11867_auto_rtlil_cc_2608_muxgate_11786
* NET 5601 = a[3]
* NET 5606 = abc_11867_new_n1019
* NET 5609 = abc_11867_new_n1016
* NET 5611 = abc_11867_new_n995
* NET 5612 = abc_11867_new_n370
* NET 5619 = abc_11867_new_n911
* NET 5624 = abc_11867_new_n898
* NET 5625 = abc_11867_new_n897
* NET 5628 = spare_buffer_45.q
* NET 5631 = abc_11867_new_n1818
* NET 5634 = abc_11867_new_n940
* NET 5637 = abc_11867_new_n1387
* NET 5638 = abc_11867_new_n1388
* NET 5641 = abc_11867_new_n938
* NET 5643 = abc_11867_new_n886
* NET 5644 = abc_11867_new_n618
* NET 5645 = abc_11867_new_n896
* NET 5647 = abc_11867_flatten_mos6502_0_adj_bcd_0_0
* NET 5651 = abc_11867_auto_rtlil_cc_2608_muxgate_11774
* NET 5656 = abc_11867_new_n1383
* NET 5660 = abc_11867_new_n1390
* NET 5662 = abc_11867_new_n1389
* NET 5666 = abc_11867_new_n1355
* NET 5668 = abc_11867_new_n1352
* NET 5669 = abc_11867_new_n1350
* NET 5673 = spare_buffer_33.q
* NET 5676 = mos6502_shift_right
* NET 5677 = abc_11867_auto_rtlil_cc_2608_muxgate_11708
* NET 5683 = abc_11867_new_n1190
* NET 5684 = abc_11867_new_n1187
* NET 5685 = abc_11867_auto_rtlil_cc_2608_muxgate_11682
* NET 5687 = subckt_1663_sff1_x4.sff_s
* NET 5692 = subckt_1663_sff1_x4.nckr
* NET 5693 = subckt_1663_sff1_x4.ckr
* NET 5694 = spare_buffer_29.q
* NET 5702 = abc_11867_new_n681
* NET 5703 = abc_11867_new_n677
* NET 5776 = abc_11867_new_n842
* NET 5785 = abc_11867_new_n1719
* NET 5789 = abc_11867_new_n1357
* NET 5790 = mos6502_alu_co
* NET 5795 = subckt_1753_sff1_x4.sff_s
* NET 5798 = subckt_1753_sff1_x4.sff_m
* NET 5801 = subckt_1753_sff1_x4.ckr
* NET 5802 = subckt_1753_sff1_x4.nckr
* NET 5803 = abc_11867_new_n1027
* NET 5805 = abc_11867_new_n1000
* NET 5810 = abc_11867_new_n351
* NET 5812 = abc_11867_new_n1023
* NET 5817 = abc_11867_new_n354
* NET 5818 = abc_11867_new_n1024
* NET 5822 = abc_11867_new_n1010
* NET 5824 = abc_11867_new_n1011
* NET 5826 = mos6502_pc[1]
* NET 5828 = subckt_1733_sff1_x4.sff_s
* NET 5831 = subckt_1733_sff1_x4.sff_m
* NET 5833 = abc_11867_auto_rtlil_cc_2608_muxgate_11814
* NET 5835 = clk_root_br_tl_0
* NET 5836 = subckt_1733_sff1_x4.ckr
* NET 5837 = subckt_1733_sff1_x4.nckr
* NET 5841 = abc_11867_new_n946
* NET 5843 = abc_11867_new_n889
* NET 5844 = abc_11867_new_n844
* NET 5848 = abc_11867_new_n939
* NET 5849 = abc_11867_new_n619_hfns_2
* NET 5851 = mos6502_alu_out[2]
* NET 5853 = abc_11867_new_n432_hfns_2
* NET 5856 = abc_11867_new_n1356
* NET 5864 = abc_11867_new_n1385
* NET 5865 = abc_11867_new_n1384
* NET 5870 = mos6502_c
* NET 5872 = mos6502_n
* NET 5877 = abc_11867_new_n1386
* NET 5879 = subckt_1679_sff1_x4.sff_s
* NET 5882 = subckt_1679_sff1_x4.sff_m
* NET 5886 = subckt_1679_sff1_x4.ckr
* NET 5887 = subckt_1679_sff1_x4.nckr
* NET 5888 = abc_11867_new_n1274
* NET 5889 = abc_11867_auto_rtlil_cc_2608_muxgate_11718
* NET 5890 = abc_11867_new_n1268
* NET 5891 = abc_11867_new_n1263
* NET 5892 = abc_11867_new_n1266
* NET 5893 = abc_11867_new_n1656
* NET 5895 = abc_11867_new_n1221
* NET 5898 = subckt_1660_sff1_x4.sff_s
* NET 5903 = subckt_1660_sff1_x4.sff_m
* NET 5905 = subckt_1660_sff1_x4.ckr
* NET 5906 = subckt_1660_sff1_x4.nckr
* NET 5907 = mos6502_sec
* NET 5908 = abc_11867_new_n1192
* NET 5910 = abc_11867_auto_rtlil_cc_2608_muxgate_11684
* NET 5911 = abc_11867_new_n1195
* NET 5912 = abc_11867_new_n1297
* NET 5914 = abc_11867_new_n1208
* NET 5915 = abc_11867_new_n756
* NET 5916 = abc_11867_new_n698
* NET 5917 = abc_11867_new_n687
* NET 5919 = abc_11867_new_n758
* NET 5920 = abc_11867_new_n746
* NET 5922 = abc_11867_new_n722
* NET 5957 = abc_11867_new_n748
* NET 5958 = mos6502_alu_ai7
* NET 5960 = subckt_1759_sff1_x4.sff_s
* NET 5965 = subckt_1759_sff1_x4.sff_m
* NET 5966 = abc_11867_auto_rtlil_cc_2608_muxgate_11866
* NET 5968 = subckt_1759_sff1_x4.ckr
* NET 5970 = subckt_1759_sff1_x4.nckr
* NET 5974 = abc_11867_new_n1358
* NET 5976 = abc_11867_auto_rtlil_cc_2608_muxgate_11854
* NET 5978 = abc_11867_new_n1892
* NET 5984 = subckt_97_nmx2_x1.q
* NET 5985 = abc_11867_new_n1026
* NET 5988 = abc_11867_new_n374
* NET 5989 = abc_11867_new_n1001
* NET 5990 = abc_11867_new_n1004
* NET 5993 = abc_11867_new_n1018
* NET 5996 = abc_11867_new_n373
* NET 5998 = mos6502_abl[7]
* NET 6000 = mos6502_abl[3]
* NET 6005 = mos6502_abl[4]
* NET 6006 = abc_11867_new_n372
* NET 6007 = abc_11867_new_n586
* NET 6008 = abc_11867_new_n1008
* NET 6021 = abc_11867_new_n428_hfns_3
* NET 6022 = mos6502_alu_out[5]
* NET 6026 = abc_11867_new_n428_hfns_4
* NET 6027 = mos6502_alu_out[4]
* NET 6029 = abc_11867_new_n485_hfns_1
* NET 6032 = abc_11867_new_n1576
* NET 6037 = abc_11867_new_n490_hfns_1
* NET 6040 = abc_11867_new_n478_hfns_2
* NET 6043 = abc_11867_new_n485_hfns_3
* NET 6048 = subckt_1708_sff1_x4.sff_s
* NET 6052 = abc_11867_auto_rtlil_cc_2608_muxgate_11764
* NET 6055 = subckt_1708_sff1_x4.sff_m
* NET 6057 = subckt_1708_sff1_x4.ckr
* NET 6059 = subckt_1708_sff1_x4.nckr
* NET 6060 = mos6502_z
* NET 6062 = mos6502_v
* NET 6072 = mos6502_adc_sbc
* NET 6073 = abc_11867_new_n1354
* NET 6075 = abc_11867_new_n1371
* NET 6077 = abc_11867_new_n433
* NET 6078 = subckt_1048_nmx2_x1.q
* NET 6080 = subckt_1670_sff1_x4.sff_s
* NET 6082 = subckt_1670_sff1_x4.sff_m
* NET 6088 = subckt_1670_sff1_x4.ckr
* NET 6089 = subckt_1670_sff1_x4.nckr
* NET 6092 = abc_11867_new_n708
* NET 6095 = abc_11867_new_n358
* NET 6104 = abc_11867_new_n1182
* NET 6106 = abc_11867_auto_rtlil_cc_2608_muxgate_11678
* NET 6107 = abc_11867_new_n676
* NET 6109 = abc_11867_new_n1210
* NET 6111 = abc_11867_new_n557
* NET 6115 = abc_11867_new_n1183
* NET 6118 = abc_11867_new_n760
* NET 6123 = abc_11867_new_n759
* NET 6125 = abc_11867_new_n1291
* NET 6128 = abc_11867_new_n718
* NET 6132 = abc_11867_new_n747
* NET 6134 = abc_11867_new_n744
* NET 6136 = abc_11867_new_n628
* NET 6138 = do[6]
* NET 6223 = mos6502_alu_bi7
* NET 6226 = subckt_1748_sff1_x4.sff_s
* NET 6227 = abc_11867_auto_rtlil_cc_2608_muxgate_11844
* NET 6229 = subckt_1748_sff1_x4.sff_m
* NET 6230 = subckt_1748_sff1_x4.ckr
* NET 6232 = clk_root_br_tr_0
* NET 6233 = subckt_1748_sff1_x4.nckr
* NET 6234 = di[6]
* NET 6235 = abc_11867_new_n1025
* NET 6238 = abc_11867_new_n419
* NET 6241 = abc_11867_new_n1017
* NET 6242 = abc_11867_new_n415
* NET 6245 = abc_11867_new_n1003
* NET 6246 = abc_11867_new_n973
* NET 6247 = abc_11867_new_n371
* NET 6250 = mos6502_abl[6]
* NET 6251 = mos6502_abl[5]
* NET 6252 = abc_11867_new_n1540
* NET 6254 = abc_11867_new_n619_hfns_1
* NET 6255 = abc_11867_new_n1506
* NET 6257 = abc_11867_new_n1514
* NET 6259 = abc_11867_new_n1726
* NET 6262 = abc_11867_new_n1748
* NET 6265 = abc_11867_new_n1770
* NET 6268 = abc_11867_new_n1793
* NET 6271 = mos6502_alu_out[7]
* NET 6272 = abc_11867_new_n432_hfns_1
* NET 6273 = abc_11867_new_n1575
* NET 6275 = abc_11867_new_n1843
* NET 6276 = abc_11867_new_n1672
* NET 6279 = abc_11867_new_n334
* NET 6281 = abc_11867_new_n1577
* NET 6282 = abc_11867_new_n478_hfns_0
* NET 6283 = mos6502_alu_out[1]
* NET 6284 = abc_11867_new_n428_hfns_1
* NET 6285 = abc_11867_new_n490_hfns_0
* NET 6286 = abc_11867_new_n485_hfns_2
* NET 6287 = abc_11867_new_n1057
* NET 6288 = abc_11867_new_n337
* NET 6290 = mos6502_alu_out[6]
* NET 6291 = abc_11867_new_n1360
* NET 6292 = abc_11867_new_n1353
* NET 6293 = abc_11867_new_n1359
* NET 6294 = abc_11867_new_n1361
* NET 6296 = abc_11867_new_n705
* NET 6298 = abc_11867_new_n707
* NET 6299 = abc_11867_new_n706
* NET 6303 = abc_11867_new_n1373
* NET 6307 = abc_11867_new_n582
* NET 6309 = abc_11867_new_n1372
* NET 6311 = mos6502_alu_out[3]
* NET 6312 = abc_11867_new_n326
* NET 6316 = mos6502_plp
* NET 6319 = abc_11867_new_n1370
* NET 6320 = abc_11867_new_n1267
* NET 6323 = abc_11867_auto_rtlil_cc_2608_muxgate_11698
* NET 6324 = mos6502_op[0]
* NET 6332 = subckt_1669_sff1_x4.sff_s
* NET 6335 = subckt_1669_sff1_x4.sff_m
* NET 6336 = subckt_1669_sff1_x4.ckr
* NET 6338 = subckt_1669_sff1_x4.nckr
* NET 6339 = mos6502_inc
* NET 6342 = subckt_1680_sff1_x4.sff_s
* NET 6345 = subckt_1680_sff1_x4.sff_m
* NET 6347 = abc_11867_auto_rtlil_cc_2608_muxgate_11720
* NET 6349 = subckt_1680_sff1_x4.ckr
* NET 6350 = subckt_1680_sff1_x4.nckr
* NET 6352 = mos6502_clv
* NET 6353 = subckt_1668_sff1_x4.sff_s
* NET 6356 = subckt_1668_sff1_x4.sff_m
* NET 6358 = abc_11867_auto_rtlil_cc_2608_muxgate_11694
* NET 6361 = clk_root_bl_tl_0
* NET 6362 = subckt_1668_sff1_x4.ckr
* NET 6363 = subckt_1668_sff1_x4.nckr
* NET 6364 = abc_11867_new_n1214
* NET 6365 = abc_11867_new_n470
* NET 6368 = abc_11867_new_n1296
* NET 6370 = abc_11867_new_n458
* NET 6372 = abc_11867_new_n750
* NET 6373 = abc_11867_new_n547
* NET 6374 = abc_11867_new_n749
* NET 6376 = abc_11867_new_n459
* NET 6377 = abc_11867_new_n457
* NET 6378 = abc_11867_new_n439
* NET 6408 = abc_11867_new_n1541
* NET 6410 = di[5]
* NET 6413 = subckt_93_nmx2_x1.q
* NET 6415 = abc_11867_new_n418
* NET 6417 = abc_11867_new_n1507
* NET 6420 = abc_11867_new_n414
* NET 6422 = abc_11867_new_n1531
* NET 6426 = abc_11867_new_n1522
* NET 6428 = abc_11867_new_n1009
* NET 6432 = abc_11867_new_n1092
* NET 6433 = abc_11867_new_n343
* NET 6438 = abc_11867_new_n1639
* NET 6439 = abc_11867_new_n1638
* NET 6446 = abc_11867_new_n1601
* NET 6447 = abc_11867_new_n1602
* NET 6453 = abc_11867_new_n1588
* NET 6455 = abc_11867_new_n1589
* NET 6458 = abc_11867_new_n1590
* NET 6462 = abc_11867_new_n1050
* NET 6466 = mos6502_d
* NET 6467 = subckt_1710_sff1_x4.sff_s
* NET 6473 = abc_11867_auto_rtlil_cc_2608_muxgate_11770
* NET 6474 = subckt_1710_sff1_x4.sff_m
* NET 6476 = subckt_1710_sff1_x4.ckr
* NET 6478 = subckt_1710_sff1_x4.nckr
* NET 6479 = subckt_1658_sff1_x4.sff_s
* NET 6485 = subckt_1658_sff1_x4.sff_m
* NET 6487 = subckt_1658_sff1_x4.ckr
* NET 6489 = abc_11867_new_n332
* NET 6490 = subckt_1658_sff1_x4.nckr
* NET 6492 = subckt_1673_sff1_x4.sff_s
* NET 6494 = subckt_1673_sff1_x4.sff_m
* NET 6500 = subckt_1673_sff1_x4.nckr
* NET 6501 = subckt_1673_sff1_x4.ckr
* NET 6502 = subckt_1676_sff1_x4.sff_s
* NET 6507 = subckt_1676_sff1_x4.sff_m
* NET 6511 = subckt_1676_sff1_x4.ckr
* NET 6512 = clk_root_bl_tr_0
* NET 6513 = subckt_1676_sff1_x4.nckr
* NET 6514 = mos6502_bit_ins
* NET 6515 = abc_11867_auto_rtlil_cc_2608_muxgate_11696
* NET 6526 = abc_11867_new_n1257
* NET 6530 = abc_11867_new_n559
* NET 6537 = abc_11867_new_n804
* NET 6541 = abc_11867_new_n558
* NET 6543 = abc_11867_new_n754
* NET 6548 = abc_11867_new_n1315
* NET 6549 = abc_11867_new_n1314
* NET 6553 = abc_11867_new_n1313
* NET 6632 = abc_11867_new_n411
* NET 6633 = abc_11867_new_n410
* NET 6635 = abc_11867_new_n1640
* NET 6637 = abc_11867_new_n1600
* NET 6644 = abc_11867_new_n441
* NET 6648 = abc_11867_auto_rtlil_cc_2608_muxgate_11674
* NET 6654 = abc_11867_new_n345
* NET 6655 = abc_11867_auto_rtlil_cc_2608_muxgate_11710
* NET 6659 = abc_11867_auto_rtlil_cc_2608_muxgate_11702
* NET 6660 = abc_11867_new_n1278
* NET 6661 = abc_11867_new_n1254
* NET 6662 = abc_11867_new_n1256
* NET 6664 = abc_11867_new_n468
* NET 6666 = abc_11867_new_n469
* NET 6668 = abc_11867_new_n696
* NET 6670 = abc_11867_new_n755
* NET 6672 = abc_11867_new_n629
* NET 6673 = abc_11867_new_n695
* NET 6674 = abc_11867_new_n721
* NET 6677 = abc_11867_new_n535
* NET 6681 = subckt_1734_sff1_x4.sff_s
* NET 6682 = subckt_1734_sff1_x4.sff_m
* NET 6684 = subckt_1734_sff1_x4.ckr
* NET 6687 = subckt_1734_sff1_x4.nckr
* NET 6688 = abc_11867_auto_rtlil_cc_2608_muxgate_11816
* NET 6690 = abc_11867_new_n1495
* NET 6691 = mos6502_dihold[6]
* NET 6692 = subckt_1696_sff1_x4.sff_s
* NET 6693 = subckt_1696_sff1_x4.sff_m
* NET 6695 = subckt_1696_sff1_x4.ckr
* NET 6698 = subckt_1696_sff1_x4.nckr
* NET 6699 = abc_11867_new_n1523
* NET 6700 = subckt_89_nmx2_x1.q
* NET 6701 = di[4]
* NET 6708 = mos6502_pc[2]
* NET 6711 = abc_11867_new_n1085
* NET 6713 = abc_11867_new_n1627
* NET 6714 = abc_11867_new_n1626
* NET 6715 = abc_11867_new_n1628
* NET 6716 = abc_11867_new_n428_hfns_2
* NET 6717 = abc_11867_new_n478_hfns_1
* NET 6718 = abc_11867_new_n485_hfns_0
* NET 6719 = abc_11867_new_n1064
* NET 6720 = abc_11867_new_n338
* NET 6721 = abc_11867_new_n1071
* NET 6726 = abc_11867_new_n1564
* NET 6727 = abc_11867_new_n1563
* NET 6728 = abc_11867_new_n1565
* NET 6735 = abc_11867_new_n424
* NET 6739 = mos6502_cond_code[1]
* NET 6744 = subckt_1659_sff1_x4.sff_s
* NET 6746 = subckt_1659_sff1_x4.ckr
* NET 6748 = subckt_1659_sff1_x4.sff_m
* NET 6751 = subckt_1659_sff1_x4.nckr
* NET 6758 = mos6502_compare
* NET 6760 = abc_11867_new_n1261
* NET 6761 = abc_11867_new_n1237
* NET 6765 = abc_11867_new_n1244
* NET 6766 = abc_11867_new_n1276
* NET 6770 = abc_11867_new_n753
* NET 6799 = subckt_1737_sff1_x4.sff_m
* NET 6801 = subckt_1737_sff1_x4.ckr
* NET 6809 = subckt_1695_sff1_x4.sff_m
* NET 6810 = subckt_1695_sff1_x4.ckr
* NET 6814 = subckt_1694_sff1_x4.sff_m
* NET 6815 = subckt_1694_sff1_x4.ckr
* NET 6816 = abc_11867_new_n1079
* NET 6817 = abc_11867_new_n1051
* NET 6818 = abc_11867_new_n1052
* NET 6819 = abc_11867_new_n1056
* NET 6820 = abc_11867_new_n1058
* NET 6821 = abc_11867_new_n1059
* NET 6825 = subckt_1671_sff1_x4.sff_m
* NET 6826 = subckt_1671_sff1_x4.ckr
* NET 6833 = subckt_1737_sff1_x4.sff_s
* NET 6838 = subckt_1737_sff1_x4.nckr
* NET 6841 = abc_11867_new_n1503
* NET 6843 = abc_11867_new_n342
* NET 6844 = abc_11867_new_n1532
* NET 6846 = abc_11867_new_n1508
* NET 6851 = subckt_1695_sff1_x4.sff_s
* NET 6852 = mos6502_dihold[5]
* NET 6855 = subckt_1695_sff1_x4.nckr
* NET 6858 = abc_11867_new_n1515
* NET 6859 = abc_11867_new_n339
* NET 6860 = abc_11867_new_n1473
* NET 6861 = abc_11867_new_n1516
* NET 6863 = subckt_1694_sff1_x4.sff_s
* NET 6864 = mos6502_dihold[4]
* NET 6869 = subckt_1694_sff1_x4.nckr
* NET 6872 = abc_11867_new_n340
* NET 6873 = abc_11867_new_n971
* NET 6874 = abc_11867_new_n1080
* NET 6878 = abc_11867_new_n619_hfns_0
* NET 6879 = abc_11867_new_n1078
* NET 6882 = abc_11867_new_n1612
* NET 6883 = abc_11867_new_n1613
* NET 6887 = abc_11867_new_n1614
* NET 6889 = abc_11867_new_n436
* NET 6893 = abc_11867_new_n1077
* NET 6900 = abc_11867_new_n1049
* NET 6908 = abc_11867_new_n377
* NET 6910 = abc_11867_new_n392
* NET 6911 = subckt_1671_sff1_x4.sff_s
* NET 6918 = subckt_1671_sff1_x4.nckr
* NET 6919 = abc_11867_auto_rtlil_cc_2608_muxgate_11676
* NET 6920 = mos6502_cond_code[2]
* NET 6925 = mos6502_op[3]
* NET 6927 = abc_11867_auto_rtlil_cc_2608_muxgate_11704
* NET 6934 = abc_11867_new_n330
* NET 6936 = abc_11867_new_n1217
* NET 6940 = abc_11867_new_n546
* NET 6946 = abc_11867_new_n1246
* NET 6947 = abc_11867_new_n1250
* NET 6950 = abc_11867_new_n1277
* NET 6954 = abc_11867_new_n1243
* NET 6955 = abc_11867_new_n751
* NET 6957 = abc_11867_new_n745
* NET 6961 = abc_11867_new_n461
* NET 6964 = abc_11867_new_n465
* NET 6966 = abc_11867_new_n685
* NET 6970 = abc_11867_new_n443
* NET 6972 = abc_11867_new_n446
* NET 6975 = do[5]
* NET 7049 = mos6502_pc[3]
* NET 7050 = subckt_1735_sff1_x4.sff_s
* NET 7053 = subckt_1735_sff1_x4.sff_m
* NET 7057 = subckt_1735_sff1_x4.nckr
* NET 7058 = subckt_1735_sff1_x4.ckr
* NET 7059 = abc_11867_new_n1505
* NET 7060 = abc_11867_auto_rtlil_cc_2608_muxgate_11818
* NET 7063 = abc_11867_new_n1511
* NET 7065 = abc_11867_new_n1501
* NET 7066 = abc_11867_new_n1492
* NET 7068 = abc_11867_new_n1524
* NET 7071 = di[3]
* NET 7073 = abc_11867_new_n408
* NET 7075 = subckt_85_nmx2_x1.q
* NET 7076 = abc_11867_new_n1002
* NET 7077 = abc_11867_new_n407
* NET 7081 = abc_11867_new_n406
* NET 7087 = abc_11867_new_n1094
* NET 7088 = abc_11867_new_n1091
* NET 7091 = abc_11867_new_n1095
* NET 7092 = abc_11867_new_n1086
* NET 7093 = abc_11867_new_n1087
* NET 7096 = abc_11867_new_n1093
* NET 7099 = abc_11867_new_n1641
* NET 7102 = abc_11867_new_n1084
* NET 7106 = abc_11867_new_n1637
* NET 7111 = abc_11867_new_n1073
* NET 7112 = abc_11867_new_n1070
* NET 7115 = abc_11867_new_n480
* NET 7116 = abc_11867_new_n1072
* NET 7118 = abc_11867_new_n970
* NET 7120 = abc_11867_new_n1065
* NET 7121 = abc_11867_new_n1066
* NET 7124 = abc_11867_new_n1063
* NET 7126 = abc_11867_new_n963
* NET 7127 = abc_11867_new_n964
* NET 7130 = subckt_1707_sff1_x4.sff_s
* NET 7133 = subckt_1707_sff1_x4.sff_m
* NET 7135 = abc_11867_auto_rtlil_cc_2608_muxgate_11762
* NET 7138 = subckt_1707_sff1_x4.nckr
* NET 7139 = subckt_1707_sff1_x4.ckr
* NET 7140 = mos6502_irhold[7]
* NET 7142 = mos6502_dimux[7]
* NET 7151 = abc_11867_new_n544
* NET 7153 = mos6502_cond_code[0]
* NET 7154 = subckt_1657_sff1_x4.sff_s
* NET 7157 = subckt_1657_sff1_x4.sff_m
* NET 7159 = abc_11867_auto_rtlil_cc_2608_muxgate_11672
* NET 7162 = subckt_1657_sff1_x4.nckr
* NET 7163 = subckt_1657_sff1_x4.ckr
* NET 7164 = abc_11867_new_n1230
* NET 7165 = abc_11867_new_n1251
* NET 7167 = abc_11867_new_n1220
* NET 7169 = abc_11867_new_n464
* NET 7170 = abc_11867_new_n1260
* NET 7171 = abc_11867_new_n1245
* NET 7173 = abc_11867_new_n460
* NET 7175 = abc_11867_new_n673
* NET 7177 = abc_11867_new_n1290
* NET 7178 = abc_11867_new_n1289
* NET 7181 = abc_11867_new_n1306
* NET 7182 = abc_11867_new_n1305
* NET 7184 = abc_11867_new_n540
* NET 7185 = abc_11867_new_n454
* NET 7227 = abc_11867_new_n1238
* NET 7228 = mos6502_pc[4]
* NET 7230 = subckt_1736_sff1_x4.sff_s
* NET 7232 = subckt_1736_sff1_x4.sff_m
* NET 7238 = subckt_1736_sff1_x4.nckr
* NET 7239 = subckt_1736_sff1_x4.ckr
* NET 7240 = abc_11867_new_n1513
* NET 7242 = abc_11867_auto_rtlil_cc_2608_muxgate_11820
* NET 7243 = abc_11867_new_n1510
* NET 7245 = abc_11867_new_n1519
* NET 7246 = abc_11867_new_n1502
* NET 7251 = abc_11867_new_n1517
* NET 7252 = abc_11867_new_n1509
* NET 7257 = mos6502_dihold[3]
* NET 7258 = subckt_1693_sff1_x4.sff_s
* NET 7261 = subckt_1693_sff1_x4.sff_m
* NET 7267 = subckt_1693_sff1_x4.nckr
* NET 7268 = subckt_1693_sff1_x4.ckr
* NET 7273 = abc_11867_new_n968_hfns_1
* NET 7275 = abc_11867_new_n1090
* NET 7277 = abc_11867_new_n367
* NET 7279 = abc_11867_new_n1088
* NET 7280 = abc_11867_new_n1083
* NET 7282 = abc_11867_new_n1625
* NET 7283 = abc_11867_new_n1629
* NET 7285 = abc_11867_new_n1615
* NET 7288 = abc_11867_new_n1603
* NET 7291 = abc_11867_new_n1599
* NET 7294 = abc_11867_new_n1611
* NET 7297 = abc_11867_new_n1578
* NET 7300 = abc_11867_new_n1591
* NET 7304 = abc_11867_new_n1587
* NET 7305 = abc_11867_new_n1574
* NET 7307 = abc_11867_new_n1472
* NET 7308 = abc_11867_new_n576
* NET 7311 = abc_11867_new_n420
* NET 7315 = abc_11867_new_n432_hfns_0
* NET 7320 = abc_11867_new_n412
* NET 7323 = abc_11867_new_n393
* NET 7326 = mos6502_dimux[3]
* NET 7329 = mos6502_op[1]
* NET 7331 = abc_11867_auto_rtlil_cc_2608_muxgate_11700
* NET 7335 = subckt_1665_sff1_x4.sff_s
* NET 7342 = subckt_1665_sff1_x4.sff_m
* NET 7344 = subckt_1665_sff1_x4.ckr
* NET 7345 = mos6502_sed
* NET 7346 = subckt_1665_sff1_x4.nckr
* NET 7347 = abc_11867_new_n1181_hfns_1
* NET 7349 = abc_11867_new_n1223
* NET 7353 = abc_11867_new_n675
* NET 7356 = abc_11867_new_n1218
* NET 7357 = abc_11867_new_n1229
* NET 7358 = abc_11867_new_n1222
* NET 7362 = abc_11867_new_n1226
* NET 7364 = abc_11867_new_n1228
* NET 7367 = abc_11867_new_n538
* NET 7373 = abc_11867_new_n1232
* NET 7381 = abc_11867_new_n1249
* NET 7382 = abc_11867_new_n1282
* NET 7391 = abc_11867_new_n1255
* NET 7394 = abc_11867_new_n437
* NET 7400 = abc_11867_new_n1248
* NET 7404 = abc_11867_new_n1188
* NET 7472 = mos6502_pc[5]
* NET 7475 = abc_11867_auto_rtlil_cc_2608_muxgate_11822
* NET 7476 = abc_11867_new_n1521
* NET 7478 = abc_11867_new_n1528
* NET 7480 = abc_11867_new_n1518
* NET 7481 = abc_11867_new_n1525
* NET 7485 = abc_11867_new_n1542
* NET 7488 = spare_buffer_42.q
* NET 7491 = abc_11867_new_n978
* NET 7492 = abc_11867_new_n394
* NET 7495 = abc_11867_new_n994
* NET 7499 = abc_11867_new_n954_hfns_1
* NET 7506 = subckt_1730_sff1_x4.sff_s
* NET 7509 = subckt_1730_sff1_x4.sff_m
* NET 7512 = subckt_1730_sff1_x4.ckr
* NET 7513 = subckt_1730_sff1_x4.nckr
* NET 7514 = mos6502_abh[6]
* NET 7515 = abc_11867_auto_rtlil_cc_2608_muxgate_11808
* NET 7521 = abc_11867_new_n366
* NET 7522 = abc_11867_new_n1642
* NET 7523 = abc_11867_new_n1636
* NET 7526 = spare_buffer_38.q
* NET 7528 = abc_11867_new_n1462
* NET 7529 = abc_11867_new_n1475
* NET 7532 = abc_11867_new_n1592
* NET 7533 = abc_11867_new_n601
* NET 7534 = abc_11867_new_n986
* NET 7535 = abc_11867_new_n507
* NET 7536 = abc_11867_new_n472
* NET 7540 = abc_11867_new_n1069
* NET 7541 = abc_11867_new_n1074
* NET 7542 = abc_11867_new_n1566
* NET 7543 = abc_11867_new_n1562
* NET 7545 = abc_11867_new_n1060
* NET 7546 = abc_11867_new_n1055
* NET 7547 = abc_11867_new_n378
* NET 7553 = mos6502_irhold[3]
* NET 7555 = subckt_1703_sff1_x4.sff_s
* NET 7558 = subckt_1703_sff1_x4.sff_m
* NET 7560 = abc_11867_auto_rtlil_cc_2608_muxgate_11754
* NET 7561 = subckt_1703_sff1_x4.ckr
* NET 7563 = subckt_1703_sff1_x4.nckr
* NET 7568 = spare_buffer_26.q
* NET 7570 = abc_11867_new_n1202
* NET 7572 = abc_11867_auto_rtlil_cc_2608_muxgate_11688
* NET 7573 = abc_11867_new_n1227
* NET 7574 = abc_11867_new_n1194
* NET 7575 = abc_11867_new_n1235
* NET 7576 = abc_11867_new_n1216
* NET 7578 = abc_11867_new_n1224
* NET 7579 = abc_11867_new_n545
* NET 7582 = abc_11867_new_n1270
* NET 7584 = spare_buffer_22.q
* NET 7588 = abc_11867_new_n1294
* NET 7589 = abc_11867_new_n1295
* NET 7592 = abc_11867_new_n674
* NET 7593 = abc_11867_new_n1198
* NET 7594 = abc_11867_new_n1303
* NET 7595 = abc_11867_new_n1304
* NET 7636 = abc_11867_new_n1543
* NET 7637 = abc_11867_new_n1527
* NET 7639 = abc_11867_new_n1534
* NET 7641 = abc_11867_new_n1533
* NET 7643 = abc_11867_new_n1479
* NET 7645 = spare_buffer_41.q
* NET 7648 = abc_11867_new_n403
* NET 7650 = abc_11867_new_n395
* NET 7655 = abc_11867_new_n402
* NET 7657 = abc_11867_new_n1579
* NET 7658 = abc_11867_new_n361
* NET 7660 = mos6502_abh[7]
* NET 7662 = subckt_1731_sff1_x4.sff_s
* NET 7667 = subckt_1731_sff1_x4.sff_m
* NET 7669 = abc_11867_auto_rtlil_cc_2608_muxgate_11810
* NET 7671 = subckt_1731_sff1_x4.ckr
* NET 7672 = subckt_1731_sff1_x4.nckr
* NET 7675 = abc_11867_new_n1635
* NET 7678 = abc_11867_new_n1624
* NET 7680 = abc_11867_new_n1630
* NET 7682 = spare_buffer_37.q
* NET 7684 = clk_root_br_0
* NET 7686 = abc_11867_new_n1081
* NET 7688 = abc_11867_new_n1076
* NET 7690 = abc_11867_new_n1048
* NET 7691 = abc_11867_new_n1053
* NET 7693 = abc_11867_new_n1067
* NET 7700 = subckt_1706_sff1_x4.sff_s
* NET 7705 = subckt_1706_sff1_x4.sff_m
* NET 7707 = abc_11867_auto_rtlil_cc_2608_muxgate_11760
* NET 7709 = subckt_1706_sff1_x4.ckr
* NET 7710 = subckt_1706_sff1_x4.nckr
* NET 7713 = abc_11867_new_n416
* NET 7716 = mos6502_irhold[6]
* NET 7718 = mos6502_dimux[6]
* NET 7723 = mos6502_dimux[4]
* NET 7727 = spare_buffer_25.q
* NET 7731 = abc_11867_new_n1200
* NET 7732 = abc_11867_new_n1197
* NET 7734 = abc_11867_new_n1225
* NET 7735 = abc_11867_new_n462
* NET 7741 = abc_11867_new_n1234
* NET 7746 = abc_11867_new_n1233
* NET 7749 = abc_11867_new_n467
* NET 7752 = abc_11867_new_n752
* NET 7756 = abc_11867_new_n1242
* NET 7757 = abc_11867_new_n1212
* NET 7759 = abc_11867_new_n1293
* NET 7761 = abc_11867_new_n672
* NET 7763 = spare_buffer_21.q
* NET 7765 = clk_root_bl_0
* NET 7767 = abc_11867_new_n1311
* NET 7770 = abc_11867_new_n1239
* NET 7771 = abc_11867_new_n1318
* NET 7826 = do[4]
* NET 7850 = abc_11867_new_n1549
* NET 7852 = abc_11867_new_n1559
* NET 7855 = abc_11867_new_n1561
* NET 7857 = abc_11867_new_n1571
* NET 7874 = abc_11867_new_n1644
* NET 7875 = abc_11867_new_n1645
* NET 7877 = abc_11867_new_n954_hfns_0
* NET 7879 = abc_11867_new_n362
* NET 7880 = abc_11867_new_n968_hfns_0
* NET 7881 = abc_11867_new_n975
* NET 7884 = abc_11867_new_n399
* NET 7887 = abc_11867_new_n398
* NET 7888 = abc_11867_new_n1062
* NET 7895 = abc_11867_new_n379
* NET 7904 = abc_11867_new_n1189
* NET 7905 = abc_11867_new_n346
* NET 7906 = abc_11867_new_n1199
* NET 7907 = abc_11867_new_n1241
* NET 7908 = abc_11867_new_n541
* NET 7912 = abc_11867_new_n1319
* NET 7913 = abc_11867_new_n1302
* NET 7927 = subckt_81_nmx2_x1.q
* NET 7928 = di[2]
* NET 7929 = abc_11867_new_n1580
* NET 7930 = abc_11867_new_n1568
* NET 7931 = subckt_73_nmx2_x1.q
* NET 7932 = abc_11867_new_n1567
* NET 7933 = abc_11867_new_n360
* NET 7934 = subckt_1692_sff1_x4.sff_s
* NET 7937 = mos6502_dihold[2]
* NET 7940 = subckt_1692_sff1_x4.sff_m
* NET 7942 = subckt_1692_sff1_x4.ckr
* NET 7944 = subckt_1692_sff1_x4.nckr
* NET 7945 = subckt_1747_sff1_x4.sff_s
* NET 7947 = mos6502_pc[15]
* NET 7948 = subckt_1747_sff1_x4.ckr
* NET 7950 = subckt_1747_sff1_x4.sff_m
* NET 7951 = abc_11867_auto_rtlil_cc_2608_muxgate_11842
* NET 7953 = subckt_1747_sff1_x4.nckr
* NET 7957 = abc_11867_new_n1643
* NET 7961 = subckt_77_nmx2_x1.q
* NET 7966 = subckt_1726_sff1_x4.sff_s
* NET 7969 = mos6502_abh[2]
* NET 7971 = subckt_1726_sff1_x4.ckr
* NET 7973 = subckt_1726_sff1_x4.sff_m
* NET 7974 = abc_11867_auto_rtlil_cc_2608_muxgate_11800
* NET 7976 = subckt_1726_sff1_x4.nckr
* NET 7984 = subckt_1704_sff1_x4.sff_s
* NET 7987 = mos6502_irhold[4]
* NET 7988 = subckt_1704_sff1_x4.sff_m
* NET 7991 = abc_11867_auto_rtlil_cc_2608_muxgate_11756
* NET 7993 = subckt_1704_sff1_x4.ckr
* NET 7995 = subckt_1704_sff1_x4.nckr
* NET 7998 = subckt_1664_sff1_x4.sff_s
* NET 8000 = mos6502_cld
* NET 8001 = subckt_1664_sff1_x4.ckr
* NET 8003 = subckt_1664_sff1_x4.sff_m
* NET 8004 = abc_11867_auto_rtlil_cc_2608_muxgate_11686
* NET 8007 = subckt_1664_sff1_x4.nckr
* NET 8010 = abc_11867_new_n435
* NET 8018 = abc_11867_new_n539
* NET 8019 = abc_11867_new_n1180
* NET 8020 = abc_11867_new_n543
* NET 8022 = abc_11867_new_n1326
* NET 8023 = abc_11867_new_n743
* NET 8026 = abc_11867_new_n1308
* NET 8027 = abc_11867_new_n1247
* NET 8029 = abc_11867_new_n1240
* NET 8030 = abc_11867_new_n741
* NET 8049 = abc_11867_new_n1545
* NET 8054 = subckt_1740_sff1_x4.sff_m
* NET 8055 = abc_11867_auto_rtlil_cc_2608_muxgate_11828
* NET 8056 = subckt_1740_sff1_x4.ckr
* NET 8060 = subckt_1741_sff1_x4.sff_m
* NET 8061 = abc_11867_auto_rtlil_cc_2608_muxgate_11830
* NET 8062 = subckt_1741_sff1_x4.ckr
* NET 8063 = abc_11867_new_n1570
* NET 8065 = rdy_hfns_0
* NET 8069 = abc_11867_new_n1582
* NET 8077 = subckt_1690_sff1_x4.sff_m
* NET 8078 = subckt_1690_sff1_x4.ckr
* NET 8082 = subckt_1746_sff1_x4.sff_m
* NET 8083 = subckt_1746_sff1_x4.ckr
* NET 8087 = subckt_1729_sff1_x4.sff_m
* NET 8088 = subckt_1729_sff1_x4.ckr
* NET 8091 = subckt_1725_sff1_x4.sff_m
* NET 8093 = subckt_1725_sff1_x4.ckr
* NET 8097 = abc_11867_new_n542
* NET 8098 = abc_11867_new_n537
* NET 8102 = subckt_1740_sff1_x4.sff_s
* NET 8103 = mos6502_pc[8]
* NET 8106 = subckt_1740_sff1_x4.nckr
* NET 8109 = subckt_1741_sff1_x4.sff_s
* NET 8110 = mos6502_pc[9]
* NET 8113 = subckt_1741_sff1_x4.nckr
* NET 8116 = abc_11867_new_n1584
* NET 8117 = abc_11867_new_n1573
* NET 8120 = subckt_1690_sff1_x4.sff_s
* NET 8121 = mos6502_dihold[0]
* NET 8126 = subckt_1690_sff1_x4.nckr
* NET 8127 = abc_11867_new_n1604
* NET 8128 = abc_11867_new_n364
* NET 8131 = abc_11867_new_n1616
* NET 8132 = abc_11867_new_n1477
* NET 8135 = rdy_hfns_3
* NET 8138 = subckt_1746_sff1_x4.sff_s
* NET 8143 = subckt_1746_sff1_x4.nckr
* NET 8145 = subckt_1729_sff1_x4.sff_s
* NET 8150 = subckt_1729_sff1_x4.nckr
* NET 8154 = subckt_1725_sff1_x4.sff_s
* NET 8159 = subckt_1725_sff1_x4.nckr
* NET 8160 = mos6502_abh[1]
* NET 8161 = abc_11867_auto_rtlil_cc_2608_muxgate_11798
* NET 8168 = mos6502_dimux[5]
* NET 8175 = abc_11867_new_n400
* NET 8185 = abc_11867_new_n396
* NET 8191 = abc_11867_new_n389
* NET 8199 = abc_11867_new_n391
* NET 8202 = abc_11867_new_n404
* NET 8207 = abc_11867_new_n435_hfns_4
* NET 8209 = abc_11867_new_n452
* NET 8215 = abc_11867_new_n435_hfns_3
* NET 8217 = abc_11867_new_n1271
* NET 8220 = abc_11867_new_n742
* NET 8222 = abc_11867_new_n442
* NET 8223 = abc_11867_new_n444
* NET 8226 = abc_11867_new_n448
* NET 8227 = abc_11867_new_n1193
* NET 8231 = abc_11867_new_n1312
* NET 8232 = abc_11867_new_n1320
* NET 8235 = abc_11867_new_n463
* NET 8236 = abc_11867_new_n536
* NET 8237 = abc_11867_new_n435_hfns_2
* NET 8240 = abc_11867_new_n447
* NET 8242 = abc_11867_new_n1310
* NET 8246 = abc_11867_new_n438
* NET 8247 = abc_11867_new_n435_hfns_1
* NET 8248 = abc_11867_new_n1309
* NET 8314 = abc_11867_new_n1539
* NET 8315 = abc_11867_new_n1547
* NET 8321 = abc_11867_new_n1546
* NET 8323 = abc_11867_new_n1535
* NET 8324 = abc_11867_new_n1556
* NET 8325 = abc_11867_new_n1544
* NET 8326 = abc_11867_new_n1526
* NET 8327 = abc_11867_new_n1558
* NET 8329 = mos6502_pc[10]
* NET 8330 = subckt_1742_sff1_x4.sff_s
* NET 8334 = subckt_1742_sff1_x4.sff_m
* NET 8335 = abc_11867_auto_rtlil_cc_2608_muxgate_11832
* NET 8338 = subckt_1742_sff1_x4.nckr
* NET 8339 = subckt_1742_sff1_x4.ckr
* NET 8343 = abc_11867_new_n1583
* NET 8346 = abc_11867_new_n1569
* NET 8347 = abc_11867_new_n1557
* NET 8348 = abc_11867_new_n1593
* NET 8349 = abc_11867_new_n1581
* NET 8350 = rdy_hfns_1
* NET 8355 = abc_11867_new_n1605
* NET 8356 = abc_11867_new_n1617
* NET 8358 = abc_11867_new_n1619
* NET 8359 = abc_11867_new_n365
* NET 8361 = abc_11867_new_n1631
* NET 8362 = abc_11867_new_n1618
* NET 8363 = mos6502_pc[14]
* NET 8366 = abc_11867_new_n1623
* NET 8367 = abc_11867_auto_rtlil_cc_2608_muxgate_11840
* NET 8368 = abc_11867_new_n1633
* NET 8369 = abc_11867_new_n1632
* NET 8372 = mos6502_abh[5]
* NET 8373 = abc_11867_auto_rtlil_cc_2608_muxgate_11806
* NET 8383 = mos6502_dihold[1]
* NET 8385 = subckt_1691_sff1_x4.sff_s
* NET 8389 = subckt_1691_sff1_x4.sff_m
* NET 8391 = subckt_1691_sff1_x4.nckr
* NET 8392 = subckt_1691_sff1_x4.ckr
* NET 8394 = abc_11867_new_n1443
* NET 8399 = mos6502_irhold[5]
* NET 8402 = subckt_1705_sff1_x4.sff_s
* NET 8404 = abc_11867_auto_rtlil_cc_2608_muxgate_11758
* NET 8405 = subckt_1705_sff1_x4.sff_m
* NET 8408 = subckt_1705_sff1_x4.ckr
* NET 8409 = subckt_1705_sff1_x4.nckr
* NET 8410 = abc_11867_new_n390
* NET 8412 = mos6502_dimux[1]
* NET 8417 = mos6502_dimux[2]
* NET 8423 = abc_11867_new_n1341
* NET 8427 = mos6502_dimux[0]
* NET 8430 = mos6502_irhold_valid
* NET 8433 = mos6502_load_reg
* NET 8434 = subckt_1698_sff1_x4.sff_s
* NET 8437 = subckt_1698_sff1_x4.sff_m
* NET 8441 = subckt_1698_sff1_x4.ckr
* NET 8442 = subckt_1698_sff1_x4.nckr
* NET 8443 = abc_11867_new_n1323
* NET 8444 = abc_11867_auto_rtlil_cc_2608_muxgate_11742
* NET 8445 = abc_11867_new_n327
* NET 8446 = abc_11867_new_n1272
* NET 8449 = subckt_950_nmx2_x1.q
* NET 8450 = abc_11867_new_n449
* NET 8451 = abc_11867_new_n1335
* NET 8454 = abc_11867_new_n1284
* NET 8455 = abc_11867_new_n456
* NET 8457 = abc_11867_new_n1328
* NET 8458 = abc_11867_new_n1213
* NET 8459 = abc_11867_new_n1329
* NET 8461 = mos6502_dst_reg[1]
* NET 8463 = subckt_1688_sff1_x4.sff_s
* NET 8466 = subckt_1688_sff1_x4.sff_m
* NET 8467 = abc_11867_auto_rtlil_cc_2608_muxgate_11736
* NET 8470 = subckt_1688_sff1_x4.ckr
* NET 8471 = subckt_1688_sff1_x4.nckr
* NET 8472 = abc_11867_new_n388
* NET 8473 = abc_11867_new_n1317
* NET 8474 = abc_11867_new_n1334
* NET 8475 = abc_11867_new_n1327
* NET 8477 = abc_11867_new_n1330
* NET 8478 = abc_11867_new_n455
* NET 8479 = abc_11867_new_n627
* NET 8480 = abc_11867_new_n440
* NET 8482 = abc_11867_new_n1325
* NET 8483 = abc_11867_new_n445
* NET 8485 = abc_11867_new_n466
* NET 8486 = abc_11867_new_n1301
* NET 8487 = abc_11867_new_n1211
* NET 8488 = abc_11867_new_n534_hfns_1
* NET 8490 = abc_11867_new_n534_hfns_0
* NET 8552 = vdd
* NET 8553 = mos6502_pc[7]
* NET 8555 = subckt_1739_sff1_x4.sff_s
* NET 8560 = subckt_1739_sff1_x4.sff_m
* NET 8561 = abc_11867_auto_rtlil_cc_2608_muxgate_11826
* NET 8564 = subckt_1739_sff1_x4.ckr
* NET 8565 = subckt_1739_sff1_x4.nckr
* NET 8566 = di[1]
* NET 8567 = abc_11867_new_n1530
* NET 8569 = abc_11867_new_n1536
* NET 8570 = abc_11867_new_n1537
* NET 8572 = mos6502_pc[6]
* NET 8573 = subckt_1738_sff1_x4.sff_s
* NET 8577 = abc_11867_auto_rtlil_cc_2608_muxgate_11824
* NET 8580 = subckt_1738_sff1_x4.sff_m
* NET 8582 = subckt_1738_sff1_x4.ckr
* NET 8584 = subckt_1738_sff1_x4.nckr
* NET 8585 = di[0]
* NET 8586 = mos6502_pc[11]
* NET 8588 = subckt_1743_sff1_x4.sff_s
* NET 8593 = subckt_1743_sff1_x4.sff_m
* NET 8596 = clk_root_br_br_0
* NET 8597 = subckt_1743_sff1_x4.ckr
* NET 8598 = subckt_1743_sff1_x4.nckr
* NET 8599 = abc_11867_new_n1586
* NET 8600 = abc_11867_auto_rtlil_cc_2608_muxgate_11834
* NET 8602 = abc_11867_new_n1595
* NET 8603 = abc_11867_new_n1596
* NET 8605 = mos6502_pc[12]
* NET 8607 = subckt_1744_sff1_x4.sff_s
* NET 8609 = subckt_1744_sff1_x4.sff_m
* NET 8615 = subckt_1744_sff1_x4.ckr
* NET 8616 = subckt_1744_sff1_x4.nckr
* NET 8617 = a[15]
* NET 8618 = abc_11867_new_n1598
* NET 8619 = abc_11867_auto_rtlil_cc_2608_muxgate_11836
* NET 8622 = abc_11867_new_n1608
* NET 8623 = abc_11867_new_n1594
* NET 8624 = abc_11867_new_n1607
* NET 8625 = abc_11867_new_n1606
* NET 8627 = rdy_hfns_2
* NET 8630 = abc_11867_new_n1620
* NET 8631 = abc_11867_new_n1610
* NET 8632 = abc_11867_new_n1621
* NET 8634 = mos6502_pc[13]
* NET 8635 = subckt_1745_sff1_x4.sff_s
* NET 8639 = abc_11867_auto_rtlil_cc_2608_muxgate_11838
* NET 8643 = subckt_1745_sff1_x4.sff_m
* NET 8645 = subckt_1745_sff1_x4.ckr
* NET 8646 = a[14]
* NET 8647 = subckt_1745_sff1_x4.nckr
* NET 8648 = mos6502_abh[4]
* NET 8650 = subckt_1728_sff1_x4.sff_s
* NET 8652 = subckt_1728_sff1_x4.sff_m
* NET 8655 = abc_11867_auto_rtlil_cc_2608_muxgate_11804
* NET 8659 = subckt_1728_sff1_x4.ckr
* NET 8660 = subckt_1728_sff1_x4.nckr
* NET 8661 = mos6502_abh[3]
* NET 8663 = subckt_1727_sff1_x4.sff_s
* NET 8665 = a[13]
* NET 8669 = subckt_1727_sff1_x4.sff_m
* NET 8670 = abc_11867_auto_rtlil_cc_2608_muxgate_11802
* NET 8672 = subckt_1727_sff1_x4.ckr
* NET 8674 = clk_root_br_bl_0
* NET 8675 = subckt_1727_sff1_x4.nckr
* NET 8677 = mos6502_irhold[1]
* NET 8678 = subckt_1701_sff1_x4.sff_s
* NET 8683 = subckt_1701_sff1_x4.sff_m
* NET 8684 = abc_11867_auto_rtlil_cc_2608_muxgate_11750
* NET 8687 = subckt_1701_sff1_x4.ckr
* NET 8688 = a[12]
* NET 8689 = subckt_1701_sff1_x4.nckr
* NET 8690 = mos6502_irhold[2]
* NET 8692 = subckt_1702_sff1_x4.sff_s
* NET 8694 = subckt_1702_sff1_x4.sff_m
* NET 8696 = abc_11867_auto_rtlil_cc_2608_muxgate_11752
* NET 8701 = subckt_1702_sff1_x4.ckr
* NET 8702 = subckt_1702_sff1_x4.nckr
* NET 8703 = mos6502_irhold[0]
* NET 8705 = subckt_1700_sff1_x4.sff_s
* NET 8710 = subckt_1700_sff1_x4.sff_m
* NET 8711 = abc_11867_auto_rtlil_cc_2608_muxgate_11748
* NET 8714 = subckt_1700_sff1_x4.ckr
* NET 8715 = subckt_1700_sff1_x4.nckr
* NET 8716 = a[11]
* NET 8717 = mos6502_shift
* NET 8719 = subckt_1678_sff1_x4.sff_s
* NET 8722 = subckt_1678_sff1_x4.sff_m
* NET 8723 = abc_11867_auto_rtlil_cc_2608_muxgate_11716
* NET 8728 = clk_root_bl_br_0
* NET 8729 = subckt_1678_sff1_x4.ckr
* NET 8730 = subckt_1678_sff1_x4.nckr
* NET 8731 = mos6502_store
* NET 8733 = subckt_1683_sff1_x4.sff_s
* NET 8735 = subckt_1683_sff1_x4.sff_m
* NET 8741 = a[10]
* NET 8742 = subckt_1683_sff1_x4.ckr
* NET 8743 = subckt_1683_sff1_x4.nckr
* NET 8744 = abc_11867_new_n1286
* NET 8745 = abc_11867_new_n1287
* NET 8746 = abc_11867_new_n1285
* NET 8747 = abc_11867_auto_rtlil_cc_2608_muxgate_11726
* NET 8750 = subckt_1681_sff1_x4.sff_s
* NET 8752 = subckt_1681_sff1_x4.sff_m
* NET 8758 = clk_root_bl_bl_0
* NET 8759 = subckt_1681_sff1_x4.ckr
* NET 8760 = subckt_1681_sff1_x4.nckr
* NET 8761 = mos6502_load_only
* NET 8763 = abc_11867_auto_rtlil_cc_2608_muxgate_11722
* NET 8764 = abc_11867_new_n1181_hfns_0
* NET 8768 = a[9]
* NET 8769 = abc_11867_new_n1333
* NET 8770 = abc_11867_new_n1331
* NET 8771 = abc_11867_new_n1332
* NET 8775 = abc_11867_new_n451
* NET 8776 = abc_11867_new_n1324
* NET 8778 = abc_11867_new_n1280
* NET 8780 = abc_11867_new_n435_hfns_0
* NET 8781 = abc_11867_new_n453
* NET 8782 = abc_11867_new_n450
* NET 8784 = abc_11867_new_n534_hfns_2
* NET 8785 = abc_11867_new_n534
* NET 8787 = vss
Mtr_16868 8552 7684 7527 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16867 7526 7527 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16866 8552 7527 7526 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16865 8552 7527 7526 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16864 7526 7527 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16863 3788 3811 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16862 4055 3812 3788 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16861 8552 3809 4055 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16860 8246 7565 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16859 7566 7723 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16858 8552 8430 7567 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16857 8552 7987 7564 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16856 7564 7567 7565 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16855 7565 8430 7566 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16854 3494 3490 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16853 3494 4111 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16852 8552 4577 3494 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16851 708 710 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16850 644 4073 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16849 8552 988 713 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16848 8552 926 643 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16847 643 713 710 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16846 710 988 644 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16845 8552 6281 6035 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16844 6035 6032 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16843 8552 6273 6035 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16842 7297 6035 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16841 8552 7684 7683 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16840 7682 7683 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16839 8552 7683 7682 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16838 8552 7683 7682 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16837 7682 7683 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16836 8552 7684 7685 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16835 8674 7685 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16834 8552 7685 8674 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16833 8552 7685 8674 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16832 8674 7685 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16831 8552 7765 5468 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16830 5467 5468 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16829 8552 5468 5467 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16828 8552 5468 5467 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16827 5467 5468 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16826 8552 7765 5674 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16825 5673 5674 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16824 8552 5674 5673 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16823 8552 5674 5673 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16822 5673 5674 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16821 8552 7765 5675 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16820 6512 5675 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16819 8552 5675 6512 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16818 8552 5675 6512 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16817 6512 5675 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16816 8552 7765 5507 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16815 5506 5507 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16814 8552 5507 5506 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16813 8552 5507 5506 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16812 5506 5507 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16811 8552 3956 3425 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16810 3425 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16809 3425 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16808 8552 8553 3425 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16807 3672 3425 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16806 4085 3859 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16805 3796 3860 3859 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16804 3797 7880 3796 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16803 3798 7881 3797 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16802 8552 7499 3798 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16801 7384 7582 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16800 8552 7757 7384 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16799 7382 7384 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16798 8552 3835 3818 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16797 3789 3835 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16796 5371 3814 3789 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16795 3789 3818 5371 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16794 8552 3816 3789 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16793 3816 3814 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16792 5181 5434 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16791 8552 5180 5181 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16790 5179 5181 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16789 8552 7765 5695 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16788 5694 5695 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16787 8552 5695 5694 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16786 8552 5695 5694 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16785 5694 5695 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16784 8552 7765 5696 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16783 6361 5696 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16782 8552 5696 6361 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16781 8552 5696 6361 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16780 6361 5696 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16779 8552 7765 7569 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16778 7568 7569 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16777 8552 7569 7568 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16776 8552 7569 7568 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16775 7568 7569 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16774 8552 7765 7728 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16773 7727 7728 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16772 8552 7728 7727 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16771 8552 7728 7727 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16770 7727 7728 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16769 8552 7765 7729 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16768 8728 7729 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16767 8552 7729 8728 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16766 8552 7729 8728 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16765 8728 7729 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16764 8552 7765 7585 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16763 7584 7585 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16762 8552 7585 7584 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16761 8552 7585 7584 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16760 7584 7585 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16759 8552 7765 7764 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16758 7763 7764 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16757 8552 7764 7763 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16756 8552 7764 7763 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16755 7763 7764 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16754 8552 7765 7766 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16753 8758 7766 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16752 8552 7766 8758 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16751 8552 7766 8758 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16750 8758 7766 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16749 790 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16748 8552 5465 790 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16747 1011 790 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16746 813 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16745 8552 5471 813 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16744 3295 813 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16743 8552 1020 810 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16742 810 1558 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16741 8552 1769 810 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16740 807 810 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16739 8552 2847 2793 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16738 2793 2795 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16737 2793 4230 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16736 8552 2798 2793 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16735 3343 2793 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16734 6379 8246 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16733 8552 8237 6379 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16732 6378 6379 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16731 8552 6029 5838 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16730 5838 6717 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16729 8552 6026 5838 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16728 6007 5838 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16727 2790 5279 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16726 8552 3006 2790 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16725 2789 2790 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16724 5934 7880 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16723 6008 6007 5934 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16722 8552 6027 6008 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16721 243 372 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16720 492 369 243 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16719 8552 1641 492 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16718 8552 6763 2258 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16717 3278 2258 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16716 8552 2258 3278 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16715 8552 2258 3278 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16714 3278 2258 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16713 8552 6763 2342 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16712 3330 2342 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16711 8552 2342 3330 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16710 8552 2342 3330 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16709 3330 2342 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16708 2469 2482 2470 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16707 2470 2471 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16706 8552 2639 2469 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16705 2907 2469 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16704 8552 5465 623 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16703 623 3753 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16702 623 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16701 8552 4139 623 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16700 824 623 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16699 8552 8020 6941 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16698 6941 7735 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16697 8552 8247 6941 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16696 6940 6941 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16695 700 707 642 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16694 641 706 700 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16693 8552 702 641 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16692 702 700 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16691 699 706 702 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16690 8552 1302 706 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16689 707 706 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16688 8552 708 705 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16687 642 705 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16686 640 639 699 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16685 8552 926 640 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16684 926 699 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16683 8552 699 926 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16682 8231 8025 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16681 8025 8490 7911 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16680 8552 8027 7911 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16679 7911 8479 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16678 7910 8242 8025 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16677 7911 8026 7910 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16676 8357 8602 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16675 8358 8355 8357 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16674 8552 8356 8358 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16673 996 994 997 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16672 997 1128 996 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16671 995 1129 997 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16670 997 992 995 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16669 1338 996 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16668 8552 1123 995 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16667 995 993 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16666 5146 4087 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16665 8552 3265 5146 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16664 8082 8083 7958 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16663 7956 8143 8082 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16662 8552 8080 7956 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16661 8080 8082 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16660 8138 8143 8080 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16659 8552 8674 8143 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16658 8083 8143 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16657 8552 8367 8142 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16656 7958 8142 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16655 7954 8039 8138 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16654 8552 8363 7954 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16653 8363 8138 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16652 8552 8138 8363 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16651 2593 2591 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16650 8552 2592 2593 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16649 8741 7545 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16648 8552 7546 8741 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16647 7125 7126 7128 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16646 7128 7127 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16645 8552 7326 7125 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16644 7124 7125 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16643 2701 2703 2603 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16642 2602 2704 2701 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16641 8552 2695 2602 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16640 2695 2701 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16639 2693 2704 2695 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16638 8552 3705 2704 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16637 2703 2704 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16636 8552 2699 2700 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16635 2603 2700 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16634 2601 2613 2693 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16633 8552 5440 2601 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16632 5440 2693 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16631 8552 2693 5440 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16630 2677 2685 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16629 8552 2936 2677 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16628 2675 2677 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16627 8552 1781 1785 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16626 1786 1783 1794 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16625 1784 1988 1786 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16624 1785 2343 1784 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16623 1465 2255 1428 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16622 8552 1956 1428 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16621 1428 2127 1465 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16620 1717 1465 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16619 2111 5150 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16618 8552 2481 2111 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16617 2235 2111 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16616 8226 8780 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16615 8226 8223 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16614 8552 8222 8226 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16613 5461 5211 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16612 5211 5215 5097 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16611 8552 5212 5097 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16610 5097 5209 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16609 5096 5363 5211 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16608 5097 5214 5096 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16607 2773 3317 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16606 2773 2771 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16605 8552 2576 2773 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16604 7364 7367 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16603 7364 7734 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16602 8552 7579 7364 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16601 7164 7167 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16600 7164 7357 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16599 8552 7573 7164 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16598 6553 8030 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16597 6553 8487 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16596 8552 7404 6553 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16595 8552 8240 6553 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16594 8234 8232 8045 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16593 8045 8231 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16592 8552 8473 8234 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16591 8467 8234 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16590 3338 3339 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16589 3340 3551 3339 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16588 3337 3544 3340 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16587 8552 3525 3337 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16586 7578 8780 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16585 7578 8020 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16584 8552 8098 7578 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16583 7183 7770 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16582 8552 8019 7183 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16581 7182 7183 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16580 8552 185 186 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16579 3320 186 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16578 8552 186 3320 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16577 8552 186 3320 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16576 3320 186 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16575 8552 3320 3321 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16574 6026 3321 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16573 8552 3321 6026 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16572 8552 3321 6026 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16571 6026 3321 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16570 8552 3320 1029 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16569 6021 1029 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16568 8552 1029 6021 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16567 8552 1029 6021 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16566 6021 1029 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16565 8552 3320 3161 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16564 6716 3161 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16563 8552 3161 6716 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16562 8552 3161 6716 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16561 6716 3161 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16560 8552 3320 3162 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16559 6284 3162 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16558 8552 3162 6284 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16557 8552 3162 6284 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16556 6284 3162 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16555 8552 3320 819 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16554 4300 819 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16553 8552 819 4300 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16552 8552 819 4300 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16551 4300 819 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16550 8552 7576 6938 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16549 6938 7353 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16548 8552 7592 6938 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16547 6936 6938 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16546 8456 8454 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16545 8552 8455 8456 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16544 8746 8456 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16543 8552 638 635 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16542 1044 635 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16541 8552 635 1044 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16540 8552 635 1044 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16539 1044 635 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16538 8552 1044 1045 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16537 3333 1045 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16536 8552 1045 3333 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16535 8552 1045 3333 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16534 3333 1045 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16533 8552 1044 634 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16532 4139 634 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16531 8552 634 4139 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16530 8552 634 4139 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16529 4139 634 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16528 8552 7228 7240 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16527 8552 8350 6803 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16526 7240 6803 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16525 6335 6336 6334 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16524 6331 6338 6335 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16523 8552 6333 6331 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16522 6333 6335 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16521 6332 6338 6333 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16520 8552 6512 6338 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16519 6336 6338 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16518 8552 6515 6337 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16517 6334 6337 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16516 6330 6329 6332 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16515 8552 6514 6330 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16514 6514 6332 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16513 8552 6332 6514 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16512 8552 2183 2184 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16511 2184 2182 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16510 8552 2789 2184 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16509 2582 2184 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16508 8552 3297 3298 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16507 3298 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16506 6873 6021 3298 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16505 3296 3294 6873 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16504 3298 3295 3296 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16503 6494 6501 6388 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16502 6387 6500 6494 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16501 8552 6493 6387 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16500 6493 6494 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16499 6492 6500 6493 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16498 8552 6512 6500 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16497 6501 6500 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16496 8552 6927 6499 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16495 6388 6499 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16494 6386 6404 6492 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16493 8552 6925 6386 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16492 6925 6492 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16491 8552 6492 6925 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16490 2711 2713 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16489 2713 2942 2616 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16488 8552 5676 2616 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16487 2616 2949 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16486 2615 2947 2713 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16485 2616 2715 2615 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16484 8552 4109 1380 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16483 1380 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16482 1380 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16481 8552 3333 1380 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16480 1591 1380 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16479 8552 6717 2006 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16478 2006 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16477 2006 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16476 8552 3333 2006 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16475 2008 2006 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16474 2944 2949 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16473 8552 5220 2944 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16472 3774 4157 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16471 3773 5915 3774 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16470 8552 3775 3773 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16469 4981 6860 4982 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16468 4982 6279 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16467 8552 4990 4981 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16466 5170 4981 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16465 3827 3648 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16464 8552 3644 3827 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16463 5522 6283 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16462 8552 5843 5522 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16461 5523 5826 5522 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16460 5522 5844 5523 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16459 5523 5621 5625 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16458 5625 8110 5523 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16457 391 2974 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16456 8552 6077 391 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16455 2376 2596 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16454 8552 2374 2376 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16453 3015 3342 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16452 8552 3181 3015 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16451 6772 6972 6675 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16450 6675 8478 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16449 8552 6970 6772 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16448 6674 6772 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16447 5505 7404 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16446 8552 6940 5505 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16445 5275 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16444 8552 5284 5275 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16443 2136 2139 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16442 8552 3275 2136 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16441 2270 2136 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16440 7286 7285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16439 8552 7294 7286 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16438 8131 7286 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16437 6964 8235 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16436 8552 8780 6964 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16435 1772 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16434 1772 6037 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16433 8552 3898 1772 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16432 6636 6720 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16431 7121 6873 6636 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16430 8552 6719 7121 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16429 1103 1318 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16428 8552 1496 1103 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16427 1310 1103 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16426 6883 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16425 6883 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16424 8552 6286 6883 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16423 8552 6022 6883 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16422 1215 2964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16421 8552 2723 1215 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16420 307 310 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16419 216 3680 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16418 8552 988 311 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16417 8552 555 217 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16416 217 311 310 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16415 310 988 216 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16414 986 989 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16413 990 2718 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16412 8552 988 991 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16411 8552 993 987 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16410 987 991 989 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16409 989 988 990 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16408 8552 3657 3021 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16407 3021 3073 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16406 3648 3246 3021 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16405 3020 3655 3648 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16404 3021 3646 3020 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16403 5014 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16402 5014 5013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16401 8552 5562 5014 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16400 8552 6758 5014 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16399 3011 2777 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16398 2632 3000 2777 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16397 2631 2775 2632 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16396 8552 2776 2631 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16395 6671 6770 8552 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16394 6670 7752 6671 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16393 6669 6769 6670 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16392 8552 6955 6669 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16391 4944 5466 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16390 4944 5851 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16389 8552 4943 4944 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16388 8552 5415 4944 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16387 944 947 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16386 945 3849 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16385 8552 1525 948 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16384 8552 1105 946 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16383 946 948 947 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16382 947 1525 945 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16381 1286 1086 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16380 1053 4073 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16379 8552 1525 1089 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16378 8552 1280 1052 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16377 1052 1089 1086 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16376 1086 1525 1053 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16375 975 976 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16374 979 2284 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16373 8552 988 978 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16372 8552 1125 977 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16371 977 978 976 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16370 976 988 979 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16369 7210 7307 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16368 7304 7308 7210 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16367 8552 7326 7304 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16366 1475 1915 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_16365 1472 1716 1405 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16364 1405 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16363 8552 1469 1408 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16362 1408 1477 1406 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16361 1406 1475 1472 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16360 1472 1915 1407 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16359 8552 3414 1469 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_16358 2119 1472 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16357 1407 1732 1408 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16356 2229 2890 8552 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16355 2344 2337 2229 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16354 2228 2338 2344 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16353 8552 6307 2228 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16352 1137 1135 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16351 8552 1138 1137 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16350 3469 1137 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16349 5626 5625 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16348 8552 5645 5626 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16347 5624 5626 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16346 8484 8782 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16345 8485 8483 8484 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16344 8552 8780 8485 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16343 6267 6276 6266 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16342 6266 7320 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16341 8552 6721 6267 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16340 6265 6267 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16339 540 548 541 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16338 541 1128 540 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16337 539 1129 541 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16336 541 542 539 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16335 2504 540 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16334 8552 1123 539 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16333 539 538 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16332 6241 6243 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16331 6243 7535 6244 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16330 8552 6420 6244 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16329 6244 6242 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16328 6240 7536 6243 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16327 6244 7533 6240 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16326 8552 4943 4497 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16325 4496 4943 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16324 4499 5466 4496 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16323 4496 4497 4499 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16322 8552 4495 4496 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16321 4495 5466 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16320 7150 8020 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16319 8552 8247 7150 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16318 7151 7150 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16317 8466 8470 8469 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16316 8464 8471 8466 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16315 8552 8465 8464 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16314 8465 8466 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16313 8463 8471 8465 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16312 8552 8758 8471 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16311 8470 8471 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16310 8552 8467 8468 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16309 8469 8468 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16308 8462 8460 8463 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16307 8552 8461 8462 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16306 8461 8463 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16305 8552 8463 8461 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16304 2261 2273 2198 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16303 2198 2274 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16302 8552 2260 2261 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16301 3262 2261 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16300 8552 1203 246 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16299 246 5470 418 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16298 6235 6237 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16297 6237 7535 6239 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16296 8552 6415 6239 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16295 6239 6238 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16294 6236 7536 6237 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16293 6239 7533 6236 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16292 6400 6433 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16291 7087 6873 6400 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16290 8552 6432 7087 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16289 3913 3915 3801 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16288 3801 3912 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16287 8552 8627 3913 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16286 4217 3913 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16285 8552 4530 1556 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16284 1556 2305 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16283 1556 2159 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16282 8552 1980 1556 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16281 1558 1556 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16280 5955 6107 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16279 6106 6115 5955 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16278 8552 6104 6106 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16277 7940 7942 7868 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16276 7866 7944 7940 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16275 8552 7939 7866 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16274 7939 7940 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16273 7934 7944 7939 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16272 8552 8674 7944 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16271 7942 7944 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16270 8552 8417 7943 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16269 7868 7943 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16268 7865 7936 7934 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16267 8552 7937 7865 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16266 7937 7934 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16265 8552 7934 7937 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16264 8342 8350 8599 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16263 8341 8586 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16262 8552 8341 8342 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16261 7705 7709 7606 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16260 7607 7710 7705 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16259 8552 7701 7607 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16258 7701 7705 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16257 7700 7710 7701 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16256 8552 8728 7710 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16255 7709 7710 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16254 8552 7707 7708 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16253 7606 7708 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16252 7605 7625 7700 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16251 8552 7716 7605 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16250 7716 7700 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16249 8552 7700 7716 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16248 5601 5388 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16247 8552 3840 5601 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16246 7626 7904 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16245 8004 7731 7626 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16244 8552 7732 8004 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16243 8315 8049 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16242 8552 8627 8315 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16241 6474 6476 6382 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16240 6381 6478 6474 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16239 8552 6469 6381 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16238 6469 6474 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16237 6467 6478 6469 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16236 8552 6512 6478 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16235 6476 6478 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16234 8552 6473 6477 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16233 6382 6477 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16232 6380 6402 6467 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16231 8552 6466 6380 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16230 6466 6467 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16229 8552 6467 6466 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16228 3640 3639 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16227 8552 4469 3640 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16226 3812 3640 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16225 3795 6720 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16224 3857 5408 3795 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16223 8552 6268 3857 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16222 1762 2151 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16221 8552 6077 1762 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16220 1959 1762 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16219 4331 4773 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16218 8552 4799 4331 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16217 4330 4331 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16216 6016 6432 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16215 8552 6254 6016 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16214 6439 6016 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16213 8447 8449 8723 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16212 8552 8764 8449 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16211 8448 8446 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16210 8723 8764 8448 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16209 8552 8445 8447 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16208 2937 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16207 2937 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16206 8552 3956 2937 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16205 8552 5826 2937 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16204 8130 8132 8036 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16203 8036 8128 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16202 8552 8127 8130 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16201 8355 8130 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16200 633 1390 632 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16199 631 2566 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16198 8552 631 633 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16197 8552 824 672 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16196 1997 822 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16195 672 823 822 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16194 8779 8778 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16193 8552 8775 8779 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16192 8776 8779 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16191 8552 1725 1461 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16190 1426 1725 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16189 1897 1723 1426 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16188 1426 1461 1897 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16187 8552 1458 1426 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16186 1458 1723 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16185 2219 2248 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16184 5186 2247 2219 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16183 8552 2723 5186 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16182 6077 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16181 6077 5562 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16180 8552 5563 6077 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16179 3005 3004 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16178 2896 2897 3004 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16177 2895 3539 2896 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16176 8552 3535 2895 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16175 7863 7931 8185 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16174 8552 8627 7931 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16173 7862 8121 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16172 8185 8627 7862 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16171 8552 8585 7863 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16170 4704 4961 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16169 8552 4971 4704 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16168 4703 4704 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16167 4095 4094 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16166 4038 4040 4094 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16165 4039 7880 4038 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16164 4037 7881 4039 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16163 8552 7877 4037 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16162 4086 5606 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16161 8552 4085 4086 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16160 4087 4086 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16159 2549 2548 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16158 8552 2572 2549 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16157 2550 2549 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16156 5636 5848 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16155 8552 5641 5636 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16154 5634 5636 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16153 2546 6037 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16152 8552 4109 2546 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16151 3133 2546 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16150 8552 3343 3344 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16149 3344 3552 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16148 8552 4237 3344 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16147 3342 3344 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16146 8552 4536 4315 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16145 4315 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16144 8552 6716 4315 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16143 5644 4315 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16142 8552 4158 4159 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16141 4374 4159 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16140 8552 4159 4374 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16139 8552 4159 4374 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16138 4374 4159 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16137 8552 4374 3908 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16136 8135 3908 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16135 8552 3908 8135 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16134 8552 3908 8135 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16133 8135 3908 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16132 8552 4374 3909 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16131 8627 3909 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16130 8552 3909 8627 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16129 8552 3909 8627 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16128 8627 3909 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16127 8552 4374 4375 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16126 8350 4375 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16125 8552 4375 8350 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16124 8552 4375 8350 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16123 8350 4375 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16122 8552 4374 4136 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16121 8065 4136 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16120 8552 4136 8065 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16119 8552 4136 8065 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16118 8065 4136 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16117 2992 2994 2991 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16116 2990 2995 2992 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16115 8552 2989 2990 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16114 2989 2992 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16113 2988 2995 2989 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16112 8552 3329 2995 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16111 2994 2995 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16110 8552 3055 2993 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16109 2991 2993 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16108 2987 2985 2988 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16107 8552 2986 2987 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16106 2986 2988 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16105 8552 2988 2986 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16104 3349 3389 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16103 3651 3390 3349 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16102 8552 3388 3651 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16101 6269 6276 6270 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16100 6270 7073 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16099 8552 6719 6269 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16098 6268 6269 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16097 199 1203 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16096 8552 5470 199 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16095 198 199 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16094 8552 5124 4942 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16093 4940 5124 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16092 4941 5130 4940 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16091 4940 4942 4941 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16090 8552 4939 4940 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16089 4939 5130 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16088 128 133 131 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16087 129 134 128 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16086 8552 127 129 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16085 127 128 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16084 125 134 127 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16083 8552 1516 134 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16082 133 134 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16081 8552 559 132 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16080 131 132 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16079 126 124 125 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16078 8552 560 126 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16077 560 125 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16076 8552 125 560 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16075 1778 2890 8552 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16074 1777 3717 1778 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16073 1776 1775 1777 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16072 8552 2159 1776 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_16071 8552 1201 1074 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16070 1074 1202 1599 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16069 8552 3898 1042 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16068 1042 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16067 1042 5013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16066 8552 4300 1042 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16065 1201 1042 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16064 2130 2707 2131 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16063 2131 2517 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16062 8552 2129 2130 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16061 2128 2130 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16060 8552 3753 1377 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16059 1377 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16058 1377 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16057 8552 4139 1377 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16056 1790 1377 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16055 8091 8093 7970 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16054 7967 8159 8091 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16053 8552 8090 7967 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16052 8090 8091 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16051 8154 8159 8090 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16050 8552 8674 8159 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16049 8093 8159 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16048 8552 8161 8158 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16047 7970 8158 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16046 7965 8041 8154 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16045 8552 8160 7965 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16044 8160 8154 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16043 8552 8154 8160 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16042 4230 6537 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16041 8552 5280 4230 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16040 3375 3750 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16039 8552 3750 3506 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16038 3503 5790 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16037 8552 3503 3375 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16036 3375 3506 3505 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16035 3505 5790 3375 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16034 3502 3505 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16033 8552 3505 3502 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16032 7570 7347 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16031 8552 7345 7570 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16030 5668 6307 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16029 8552 6077 5668 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16028 4503 4501 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16027 4503 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16026 8552 7315 4503 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16025 8552 3657 2225 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16024 2225 2270 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16023 2272 2267 2225 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16022 2224 3655 2272 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16021 2225 2268 2224 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16020 1756 1757 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16019 1951 1758 1756 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16018 8552 2260 1951 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16017 1892 2255 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16016 8552 2127 1892 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16015 1890 1892 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16014 3715 3716 3714 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16013 8552 3860 3714 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16012 3714 3717 3715 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16011 3875 3715 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16010 3680 3682 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16009 3683 4281 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16008 8552 4075 3684 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16007 8552 8417 3681 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16006 3681 3684 3682 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16005 3682 4075 3683 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16004 7643 4988 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16003 7643 5438 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16002 8552 5557 7643 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16001 8365 8627 8366 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16000 8364 8363 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15999 8552 8364 8365 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15998 7185 8781 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15997 8552 8780 7185 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15996 2337 3753 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15995 2337 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15994 8552 6717 2337 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15993 4988 6026 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15992 4988 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15991 8552 6029 4988 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15990 4984 6026 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15989 4984 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15988 8552 6717 4984 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15987 1141 1144 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15986 1057 2718 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15985 8552 1525 1146 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15984 8552 1140 1056 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15983 1056 1146 1144 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15982 1144 1525 1057 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15981 5087 5171 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15980 5427 5166 5087 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15979 8552 8065 5427 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15978 2492 2498 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_15977 2497 2500 2491 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15976 2491 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15975 8552 2493 2495 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15974 2495 2670 2494 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15973 2494 2492 2497 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15972 2497 2498 2496 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15971 8552 3414 2493 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_15970 2671 2497 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15969 2496 2930 2495 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15968 8552 2008 1854 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15967 2343 2004 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15966 1854 2005 2004 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15965 4532 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15964 4532 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15963 8552 3956 4532 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15962 937 734 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15961 652 4073 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15960 8552 779 735 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15959 8552 931 651 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15958 651 735 734 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15957 734 779 652 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15956 1513 1343 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15955 1344 2284 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15954 8552 1525 1345 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15953 8552 1505 1342 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15952 1342 1345 1343 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15951 1343 1525 1344 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15950 960 963 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15949 962 3680 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15948 8552 1525 964 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15947 8552 959 961 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15946 961 964 963 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15945 963 1525 962 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15944 5919 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15943 5919 7353 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15942 8552 7184 5919 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15941 8552 8490 5919 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15940 5915 6940 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15939 5915 6673 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15938 8552 7592 5915 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15937 8552 8490 5915 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15936 2160 3956 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15935 2160 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15934 8552 3767 2160 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15933 550 551 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15932 553 3849 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15931 8552 779 552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15930 8552 548 549 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15929 549 552 551 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15928 551 779 553 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15927 8552 6307 4760 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15926 4760 4999 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15925 8552 6077 4760 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15924 5212 4760 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15923 8552 3657 1740 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15922 1740 1741 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15921 1738 1926 1740 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15920 1739 3655 1738 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15919 1740 1923 1739 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15918 7540 7109 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15917 7110 8128 7109 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15916 7107 7880 7110 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15915 7108 7881 7107 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15914 8552 7877 7108 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15913 2735 2746 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15912 8552 8135 2735 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15911 2734 2735 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15910 5913 6368 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15909 8552 8019 5913 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15908 5912 5913 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15907 8552 3460 3461 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15906 3861 3461 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15905 8552 3461 3861 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15904 8552 3461 3861 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15903 3861 3461 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15902 8552 3861 3862 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15901 7499 3862 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15900 8552 3862 7499 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15899 8552 3862 7499 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15898 7499 3862 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15897 8552 3861 3708 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15896 7877 3708 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15895 8552 3708 7877 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15894 8552 3708 7877 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15893 7877 3708 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15892 6097 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15891 8552 6095 6097 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15890 6761 6097 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15889 6849 7228 6777 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15888 8552 6861 6777 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15887 6777 7643 6849 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15886 7251 6849 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15885 3486 3956 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15884 8552 5465 3486 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15883 3744 3486 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15882 322 327 222 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15881 221 326 322 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15880 8552 319 221 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15879 319 322 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15878 318 326 319 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15877 8552 1516 326 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15876 327 326 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15875 8552 328 325 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15874 222 325 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15873 220 240 318 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15872 8552 765 220 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15871 765 318 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15870 8552 318 765 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15869 8552 3657 1726 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15868 1726 1907 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15867 1725 1902 1726 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15866 1724 3655 1725 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15865 1726 1723 1724 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15864 8621 8622 8510 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15863 8552 8618 8510 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15862 8510 8624 8621 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15861 8619 8621 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15860 8552 805 180 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15859 180 2974 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15858 8552 5033 180 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15857 179 180 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15856 8552 4792 1770 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15855 1770 2572 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15854 8552 2334 1770 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15853 1769 1770 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15852 7642 8572 7597 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15851 8552 7641 7597 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15850 7597 7643 7642 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15849 8323 7642 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15848 285 288 209 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15847 210 290 285 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15846 8552 282 210 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15845 282 285 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15844 281 290 282 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15843 8552 1302 290 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15842 288 290 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15841 8552 291 289 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15840 209 289 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15839 208 238 281 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15838 8552 538 208 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15837 538 281 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15836 8552 281 538 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15835 2908 2911 2909 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15834 2909 2907 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15833 8552 2906 2908 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15832 3826 2908 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15831 8552 5471 3332 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15830 3332 5562 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15829 3332 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15828 8552 4139 3332 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15827 5280 3332 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15826 8552 5046 5047 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15825 5047 5043 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15824 5044 5280 5047 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15823 5045 6957 5044 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15822 5047 8023 5045 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15821 8609 8615 8509 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15820 8508 8616 8609 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15819 8552 8608 8508 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15818 8608 8609 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15817 8607 8616 8608 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15816 8552 8674 8616 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15815 8615 8616 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15814 8552 8619 8614 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15813 8509 8614 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15812 8507 8506 8607 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15811 8552 8605 8507 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15810 8605 8607 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15809 8552 8607 8605 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15808 2260 1763 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15807 2260 1537 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15806 8552 1771 2260 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15805 8552 2986 7536 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15804 8552 1567 368 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15803 7536 368 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15802 8569 8323 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15801 8552 8326 8569 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15800 4206 4061 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15799 8552 4646 4206 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15798 2127 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15797 2127 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15796 8552 3490 2127 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15795 8552 7049 2127 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15794 2914 3085 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15793 8552 2936 2914 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15792 3246 2914 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15791 8552 1567 372 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15790 8552 2986 373 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15789 372 373 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15788 4083 4690 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15787 8552 4079 4083 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15786 7974 7697 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15785 7604 8741 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15784 8552 8394 7698 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15783 8552 7969 7603 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15782 7603 7698 7697 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15781 7697 8394 7604 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15780 8655 8379 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15779 8380 8688 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15778 8552 8394 8381 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15777 8552 8648 8378 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15776 8378 8381 8379 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15775 8379 8394 8380 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15774 7515 7517 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15773 7518 8646 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15772 8552 8394 7519 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15771 8552 7514 7516 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15770 7516 7519 7517 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15769 7517 8394 7518 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15768 6452 6719 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15767 8552 6878 6452 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15766 6453 6452 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15765 8552 4577 4561 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15764 4561 6717 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15763 4561 5562 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15762 8552 8717 4561 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15761 4787 4561 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15760 245 1203 415 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15759 414 5470 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15758 8552 414 245 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15757 5407 5408 5409 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15756 5409 6872 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15755 8552 6262 5407 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15754 5406 5407 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15753 3518 4139 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15752 8552 5036 3518 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15751 3516 3518 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15750 5290 5294 5076 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15749 5077 5295 5290 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15748 8552 5286 5077 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15747 5286 5290 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15746 5285 5295 5286 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15745 8552 6361 5295 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15744 5294 5295 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15743 8552 5292 5293 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15742 5076 5293 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15741 5075 5110 5285 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15740 8552 5284 5075 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15739 5284 5285 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15738 8552 5285 5284 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15737 8552 2567 2349 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15736 2349 2346 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15735 8552 3317 2349 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15734 2587 2349 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15733 7117 7115 7119 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15732 7119 7118 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15731 8552 8648 7117 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15730 7116 7117 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15729 7854 8135 7855 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15728 7921 8110 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15727 8552 7921 7854 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15726 5965 5968 5925 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15725 5926 5970 5965 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15724 8552 5961 5926 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15723 5961 5965 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15722 5960 5970 5961 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15721 8552 6232 5970 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15720 5968 5970 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15719 8552 5966 5969 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15718 5925 5969 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15717 5924 5923 5960 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15716 8552 5958 5924 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15715 5958 5960 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15714 8552 5960 5958 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15713 6825 6826 6742 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15712 6743 6918 6825 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15711 8552 6823 6743 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15710 6823 6825 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15709 6911 6918 6823 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15708 8552 8728 6918 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15707 6826 6918 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15706 8552 7331 6917 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15705 6742 6917 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15704 6741 6794 6911 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15703 8552 7329 6741 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15702 7329 6911 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15701 8552 6911 7329 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15700 1496 3254 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15699 8552 3673 1496 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15698 7677 7875 7602 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15697 8552 7675 7602 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15696 7602 7874 7677 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15695 7951 7677 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15694 3341 3553 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15693 8552 3776 3341 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15692 8423 4217 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15691 8552 4553 8423 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15690 5776 4529 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15689 8552 4530 5776 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15688 8775 8782 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15687 8552 8780 8775 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15686 6307 3753 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15685 6307 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15684 8552 6029 6307 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15683 333 336 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15682 226 3709 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15681 8552 983 337 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15680 8552 764 225 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15679 225 337 336 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15678 336 983 226 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15677 5265 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15676 8552 5263 5265 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15675 5684 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15674 8552 5565 5684 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15673 6446 6026 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15672 6446 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15671 8552 6029 6446 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15670 8552 6027 6446 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15669 1955 5183 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15668 8552 1951 1955 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15667 1952 1955 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15666 1908 2508 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15665 8552 3269 1908 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15664 1907 1908 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15663 3539 4153 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15662 8552 4148 3539 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15661 8552 7937 7655 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15660 8552 8135 7656 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15659 7655 7656 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15658 4951 4698 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15657 4698 7535 4615 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15656 8552 4723 4615 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15655 4615 4697 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15654 4614 7536 4698 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15653 4615 7533 4614 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15652 980 982 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15651 985 2284 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15650 8552 983 984 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15649 8552 1124 981 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15648 981 984 982 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15647 982 983 985 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15646 7271 8132 7197 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15645 7197 7658 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15644 8552 7657 7271 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15643 7929 7271 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15642 8602 8346 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15641 8602 8348 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15640 8552 8349 8602 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15639 8552 8347 8602 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15638 8552 3677 2932 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15637 2932 3678 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15636 8552 7723 2932 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15635 2931 2932 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15634 6438 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15633 6438 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15632 8552 6286 6438 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15631 8552 6271 6438 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15630 1754 1758 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15629 1753 1757 1754 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15628 8552 2723 1753 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15627 3000 2998 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15626 3000 2999 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15625 8552 3326 3000 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15624 5088 7880 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15623 5180 6007 5088 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15622 8552 6283 5180 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15621 2745 2572 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15620 2745 4792 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15619 8552 4530 2745 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15618 8552 2159 2745 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15617 680 565 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15616 568 2284 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15615 8552 779 567 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15614 8552 1127 566 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15613 566 567 565 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15612 565 779 568 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15611 559 563 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15610 562 3680 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15609 8552 779 564 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15608 8552 560 561 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15607 561 564 563 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15606 563 779 562 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15605 8552 7257 7081 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15604 8552 8065 7082 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15603 7081 7082 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15602 715 718 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15601 646 4073 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15600 8552 983 719 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15599 8552 925 645 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15598 645 719 718 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15597 718 983 646 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15596 8552 4520 4521 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15595 4521 4714 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15594 8552 4518 4521 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15593 4519 4521 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15592 4093 5824 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15591 8552 4095 4093 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15590 4092 4093 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15589 5119 5466 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15588 5119 6290 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15587 8552 5790 5119 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15586 8552 5415 5119 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15585 8044 8226 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15584 8457 8220 8044 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15583 8552 8454 8457 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15582 1520 5214 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15581 8552 1522 1520 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15580 1757 1520 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15579 7741 7743 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15578 7743 8220 7628 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15577 8552 8247 7628 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15576 7628 8235 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15575 7627 8455 7743 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15574 7628 7746 7627 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15573 2561 2890 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15572 2560 4792 2562 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15571 2569 2562 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15570 2562 6878 2561 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15569 8552 3048 2560 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15568 3270 4502 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15567 3271 5408 3270 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15566 8552 4096 3271 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15565 8552 4536 3889 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15564 3889 6040 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15563 8552 3964 3889 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15562 4075 3889 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15561 364 7536 242 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15560 242 1016 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15559 8552 6077 364 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15558 363 364 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15557 4229 4362 4197 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15556 4196 4364 4229 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15555 8552 4227 4196 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15554 4227 4229 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15553 4357 4364 4227 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15552 8552 6361 4364 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15551 4362 4364 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15550 8552 4823 4363 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15549 4197 4363 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15548 4195 4194 4357 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15547 8552 4358 4195 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15546 4358 4357 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15545 8552 4357 4358 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15544 725 726 648 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15543 648 1128 725 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15542 647 1129 648 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15541 648 720 647 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15540 2252 725 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15539 8552 1123 647 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15538 647 721 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15537 8552 7761 6960 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15536 6960 8490 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15535 8552 8240 6960 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15534 6957 6960 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15533 8552 6940 5509 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15532 5509 6673 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15531 5509 7184 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15530 8552 8490 5509 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15529 5508 5509 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15528 7326 7073 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15527 8417 8202 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15526 8552 3490 402 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15525 402 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15524 402 5192 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15523 8552 5465 402 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15522 499 402 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15521 6249 6246 6248 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15520 6248 6247 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15519 8552 7076 6249 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15518 6245 6249 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15517 3366 3469 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15516 3866 3462 3366 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15515 8552 4092 3866 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15514 6891 7126 6783 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15513 6783 7127 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15512 8552 7142 6891 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15511 7088 6891 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15510 8077 8078 7941 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15509 7938 8126 8077 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15508 8552 8075 7938 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15507 8075 8077 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15506 8120 8126 8075 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15505 8552 8674 8126 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15504 8078 8126 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15503 8552 8427 8124 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15502 7941 8124 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15501 7935 8035 8120 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15500 8552 8121 7935 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15499 8121 8120 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15498 8552 8120 8121 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15497 1747 1498 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15496 8552 1496 1747 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15495 4098 6276 4097 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15494 4097 8185 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15493 8552 4099 4098 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15492 4096 4098 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15491 3367 3472 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15490 7826 3469 3367 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15489 8552 3718 7826 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15488 7533 3898 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15487 8552 6717 7533 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15486 2148 4979 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15485 8552 1954 2148 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15484 7988 7993 7899 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15483 7897 7995 7988 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15482 8552 7989 7897 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15481 7989 7988 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15480 7984 7995 7989 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15479 8552 8728 7995 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15478 7993 7995 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15477 8552 7991 7992 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15476 7899 7992 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15475 7896 7986 7984 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15474 8552 7987 7896 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15473 7987 7984 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15472 8552 7984 7987 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15471 1966 2566 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15470 1966 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15469 8552 4577 1966 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15468 6887 8372 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15467 6887 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15466 8552 7315 6887 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15465 3336 5510 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15464 3335 3334 3336 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15463 8552 3333 3335 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15462 2685 3082 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15461 2685 2933 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15460 8552 2927 2685 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15459 8552 3083 2685 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15458 3401 3400 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15457 8552 3429 3401 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15456 3658 3401 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15455 4487 5415 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15454 4487 4943 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15453 8552 5466 4487 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15452 5600 5604 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15451 5517 5601 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15450 8552 8394 5605 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15449 8552 6000 5516 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15448 5516 5605 5604 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15447 5604 8394 5517 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15446 5402 5147 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15445 5063 5146 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15444 8552 8394 5149 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15443 8552 6251 5062 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15442 5062 5149 5147 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15441 5147 8394 5063 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15440 4215 4082 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15439 4080 4083 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15438 8552 8394 4084 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15437 8552 5998 4081 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15436 4081 4084 4082 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15435 4082 8394 4080 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15434 8552 2277 1934 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15433 1934 2937 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15432 8552 3657 1934 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15431 1931 1934 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15430 8552 2508 1730 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15429 1730 3269 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15428 8552 3657 1730 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15427 1729 1730 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15426 1768 3136 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15425 1768 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15424 8552 6718 1768 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15423 1546 1369 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15422 1546 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15421 8552 3753 1546 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15420 2209 3048 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15419 2208 2334 2336 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15418 3318 2336 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15417 2336 2337 2209 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15416 8552 2890 2208 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15415 3007 5279 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15414 8552 3006 3007 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15413 5080 7880 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15412 5142 6007 5080 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15411 8552 6271 5142 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15410 2293 2147 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15409 2149 2148 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15408 8552 8394 2150 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15407 8552 5188 2146 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15406 2146 2150 2147 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15405 2147 8394 2149 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15404 3269 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15403 3269 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15402 8552 3956 3269 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15401 8552 6708 3269 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15400 3049 2971 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15399 2891 2890 2971 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15398 2889 3314 2891 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15397 8552 3315 2889 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15396 1298 5214 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15395 8552 1297 1298 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15394 2251 1298 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15393 2738 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15392 8552 3956 2738 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15391 3297 2738 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15390 2767 2784 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15389 8552 4577 2767 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15388 3164 2767 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15387 6973 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15386 8552 8780 6973 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15385 6972 6973 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15384 5994 6246 5933 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15383 5933 5996 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15382 8552 6241 5994 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15381 5993 5994 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15380 3722 7118 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15379 3723 7115 3722 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15378 8552 4522 3723 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15377 1210 1212 1062 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15376 1061 1214 1210 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15375 8552 1206 1061 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15374 1206 1210 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15373 1204 1214 1206 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15372 8552 2028 1214 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15371 1212 1214 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15370 8552 2191 1213 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15369 1062 1213 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15368 1060 1059 1204 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15367 8552 1203 1060 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15366 1203 1204 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15365 8552 1204 1203 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15364 8552 5915 5918 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15363 5918 5919 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15362 5918 5916 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15361 8552 5917 5918 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15360 6123 5918 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15359 8552 1996 1852 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15358 1852 1995 2171 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15357 5672 5668 5534 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15356 5534 5669 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15355 8552 5666 5672 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15354 5856 5672 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15353 752 759 660 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15352 659 761 752 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15351 8552 753 659 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15350 753 752 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15349 751 761 753 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15348 8552 1516 761 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15347 759 761 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15346 8552 680 760 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15345 660 760 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15344 658 657 751 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15343 8552 1127 658 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15342 1127 751 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15341 8552 751 1127 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15340 2265 2263 2199 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15339 2199 2511 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15338 8552 2936 2265 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15337 2267 2265 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15336 8552 6286 3322 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15335 3322 3749 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15334 3322 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15333 8552 6716 3322 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15332 3334 3322 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15331 8552 1790 1792 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15330 1792 1791 2170 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15329 8552 5470 1177 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15328 1177 1203 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15327 1177 1390 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15326 8552 2566 1177 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15325 2784 1177 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15324 5547 5598 5394 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15323 5393 5599 5547 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15322 8552 5545 5393 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15321 5545 5547 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15320 5593 5599 5545 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15319 8552 6232 5599 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15318 5598 5599 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15317 8552 5600 5597 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15316 5394 5597 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15315 5391 5515 5593 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15314 8552 6000 5391 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15313 6000 5593 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15312 8552 5593 6000 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15311 2537 2151 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15310 8552 6077 2537 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15309 5580 4693 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15308 8552 3838 5580 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15307 2191 2372 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15306 8552 2374 2191 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15305 599 609 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15304 599 363 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15303 8552 360 599 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15302 4213 4275 4177 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15301 4176 4276 4213 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15300 8552 4212 4176 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15299 4212 4213 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15298 4268 4276 4212 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15297 8552 6232 4276 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15296 4275 4276 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15295 8552 4215 4274 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15294 4177 4274 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15293 4175 4174 4268 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15292 8552 5998 4175 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15291 5998 4268 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15290 8552 4268 5998 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15289 2123 3857 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15288 2122 2121 2123 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15287 8552 3261 2122 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15286 3538 3765 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15285 8552 5044 3538 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15284 6104 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15283 8552 6316 6104 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15282 5089 5174 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15281 5171 5169 5089 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15280 8552 5170 5171 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15279 7617 7658 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15278 8349 8132 7617 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15277 8552 7657 8349 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15276 2277 8412 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15275 2277 3677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15274 8552 3678 2277 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15273 4104 4529 4042 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15272 8552 8359 4042 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15271 4042 4530 4104 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15270 4105 4104 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15269 6298 6300 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15268 6301 6299 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15267 8552 6739 6302 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15266 8552 6296 6297 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15265 6297 6302 6300 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15264 6300 6739 6301 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15263 8480 8246 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15262 8552 8215 8480 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15261 2559 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15260 2559 6717 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15259 8552 5562 2559 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15258 6722 6721 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15257 8552 6878 6722 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15256 6637 6722 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15255 8369 8625 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15254 8369 8361 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15253 8552 8362 8369 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15252 8552 8623 8369 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15251 2548 5470 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15250 2548 3753 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15249 8552 5563 2548 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15248 6296 6063 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15247 5940 6062 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15246 8552 6920 6065 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15245 8552 6060 5939 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15244 5939 6065 6063 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15243 6063 6920 5940 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15242 5916 7184 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15241 5916 6673 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15240 8552 6940 5916 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15239 8552 8490 5916 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15238 7172 8222 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15237 7173 8246 7172 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15236 8552 8247 7173 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15235 2161 5562 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15234 2161 6717 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15233 8552 3964 2161 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15232 8552 1702 1445 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15231 1425 1702 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15230 1879 1447 1425 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15229 1425 1445 1879 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15228 8552 1443 1425 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15227 1443 1447 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15226 8552 4027 3301 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15225 3301 4533 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15224 8552 3300 3301 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15223 4327 3301 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15222 3498 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15221 3498 3749 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15220 8552 6286 3498 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15219 8552 6716 3498 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15218 6711 6026 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15217 6711 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15216 8552 6717 6711 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15215 8552 7514 6711 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15214 4068 4070 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15213 4069 4941 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15212 8552 4075 4072 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15211 8552 7718 4071 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15210 4071 4072 4070 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15209 4070 4075 4069 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15208 4184 4306 6735 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15207 8552 8350 4306 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15206 4185 4727 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15205 6735 8350 4185 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15204 8552 4305 4184 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15203 8552 6027 3809 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15202 8552 8627 3810 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15201 3809 3810 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15200 8552 3648 3385 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15199 3346 3648 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15198 3825 3644 3346 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15197 3346 3385 3825 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15196 8552 3382 3346 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15195 3382 3644 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15194 7295 7528 7209 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15193 7209 7529 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15192 8552 7947 7295 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15191 7523 7295 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15190 5649 6072 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15189 8552 6466 5649 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15188 5647 5649 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15187 1802 2764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15186 8552 4577 1802 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15185 2015 1802 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15184 7583 8030 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15183 8552 8240 7583 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15182 8023 7583 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15181 8552 8483 6771 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15180 6771 8222 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15179 8552 8237 6771 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15178 6673 6771 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15177 7192 7251 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15176 7245 7243 7192 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15175 8552 8350 7245 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15174 7477 7478 7479 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15173 8552 7476 7479 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15172 7479 7637 7477 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15171 7475 7477 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15170 1288 1290 1287 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15169 1284 1291 1288 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15168 8552 1283 1284 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15167 1283 1288 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15166 1281 1291 1283 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15165 8552 1302 1291 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15164 1290 1291 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15163 8552 1286 1289 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15162 1287 1289 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15161 1282 1279 1281 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15160 8552 1280 1282 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15159 1280 1281 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15158 8552 1281 1280 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15157 8552 1552 1549 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15156 1549 1553 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15155 1549 1772 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15154 8552 2559 1549 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15153 2974 1549 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15152 3163 3168 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15151 3168 5046 3041 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15150 8552 5280 3041 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15149 3041 6111 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15148 3040 3164 3168 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15147 3041 3165 3040 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15146 8552 6282 3760 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15145 3760 3767 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15144 8552 5562 3760 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15143 7115 3760 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15142 1885 1882 1814 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15141 1814 2105 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15140 8552 1883 1885 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15139 2108 1885 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15138 6724 7115 6639 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15137 6639 7118 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15136 8552 8160 6724 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15135 6817 6724 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15134 8580 8582 8500 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15133 8499 8584 8580 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15132 8552 8575 8499 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15131 8575 8580 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15130 8573 8584 8575 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15129 8552 8596 8584 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15128 8582 8584 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15127 8552 8577 8583 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15126 8500 8583 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15125 8498 8497 8573 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15124 8552 8572 8498 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15123 8572 8573 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15122 8552 8573 8572 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15121 59 61 58 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15120 60 63 59 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15119 8552 57 60 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15118 57 59 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15117 55 63 57 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15116 8552 1302 63 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15115 61 63 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15114 8552 259 62 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15113 58 62 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15112 54 53 55 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15111 8552 274 54 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15110 274 55 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15109 8552 55 274 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15108 2263 2139 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15107 8552 3275 2263 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15106 4714 7643 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15105 8552 4715 4714 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15104 2138 3445 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15103 8552 2137 2138 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15102 3154 3502 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15101 8552 4139 3154 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15100 5237 5239 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15099 5071 5440 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15098 8552 6312 5240 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15097 8552 5365 5070 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15096 5070 5240 5239 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15095 5239 6312 5071 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15094 8334 8339 8337 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15093 8332 8338 8334 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15092 8552 8333 8332 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15091 8333 8334 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15090 8330 8338 8333 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15089 8552 8596 8338 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15088 8339 8338 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15087 8552 8335 8336 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15086 8337 8336 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15085 8331 8328 8330 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15084 8552 8329 8331 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15083 8329 8330 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15082 8552 8330 8329 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15081 6406 6770 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15080 6407 6955 6544 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15079 6543 6544 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15078 6544 7752 6406 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15077 8552 6668 6407 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15076 4498 6283 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15075 4498 4499 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15074 8552 5415 4498 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15073 4584 4587 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15072 4585 6125 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15071 8552 8764 4588 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15070 8552 4583 4586 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15069 4586 4588 4587 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15068 4587 8764 4585 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15067 1361 4027 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15066 8552 2159 1361 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15065 1539 1361 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15064 1318 1320 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15063 1321 3254 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15062 8552 1862 1322 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15061 8552 3673 1319 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15060 1319 1322 1320 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15059 1320 1862 1321 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15058 2927 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15057 2927 6043 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15056 8552 3956 2927 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15055 8552 7228 2927 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15054 7100 7099 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15053 8552 7106 7100 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15052 7522 7100 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15051 5528 5643 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15050 5641 5644 5528 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15049 8552 6062 5641 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15048 3936 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15047 3936 4135 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15046 8552 6718 3936 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15045 8552 5471 3936 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15044 6136 8490 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15043 8552 8240 6136 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15042 7917 8321 7853 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15041 7853 8324 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15040 8552 8627 7917 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15039 7852 7917 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15038 6463 6462 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15037 8552 6878 6463 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15036 6727 6463 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15035 5108 6115 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15034 5274 5505 5108 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15033 8552 5272 5274 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15032 6427 6426 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15031 8552 6878 6427 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15030 6699 6427 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15029 1019 4529 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15028 1019 4750 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15027 8552 1553 1019 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15026 8552 1552 1019 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15025 1065 1114 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15024 1323 1113 1065 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15023 8552 2260 1323 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15022 927 931 929 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15021 929 1128 927 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15020 928 1129 929 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15019 929 925 928 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15018 2248 927 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15017 8552 1123 928 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15016 928 926 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15015 4701 5160 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15014 8552 4744 4701 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15013 4700 4701 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15012 4157 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15011 4157 5562 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15010 8552 5471 4157 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15009 8552 4139 4157 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15008 8552 7049 7059 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15007 8552 8065 6805 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15006 7059 6805 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15005 8552 5013 3511 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15004 3511 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15003 3511 6026 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15002 8552 4139 3511 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15001 3512 3511 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15000 8552 6040 1371 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14999 1371 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14998 1371 4577 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14997 8552 5465 1371 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14996 1566 1371 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14995 7342 7344 7224 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14994 7223 7346 7342 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14993 8552 7337 7223 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14992 7337 7342 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14991 7335 7346 7337 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14990 8552 8728 7346 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14989 7344 7346 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14988 8552 7572 7343 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14987 7224 7343 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14986 7222 7221 7335 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14985 8552 7345 7222 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14984 7345 7335 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14983 8552 7335 7345 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14982 8552 2176 2175 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14981 2175 2571 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14980 2175 2350 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14979 8552 2174 2175 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14978 2173 2175 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14977 2232 3009 2372 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14976 2373 2592 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14975 8552 2373 2232 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14974 2970 3049 2979 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14973 2969 2968 2970 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14972 8552 3307 2969 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14971 8552 4143 2583 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14970 2583 2582 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14969 2583 2587 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14968 8552 2783 2583 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14967 2591 2583 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14966 6897 7126 6787 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14965 6787 7127 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14964 8552 7723 6897 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14963 7112 6897 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14962 5542 5577 5368 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14961 5369 5578 5542 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14960 8552 5540 5369 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14959 5540 5542 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14958 5572 5578 5540 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14957 8552 6232 5578 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14956 5577 5578 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14955 8552 5543 5576 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14954 5368 5576 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14953 5367 5512 5572 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14952 8552 6271 5367 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14951 6271 5572 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14950 8552 5572 6271 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14949 6278 6276 6277 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14948 6277 8175 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14947 8552 6462 6278 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14946 6275 6278 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14945 2617 3297 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14944 8552 3531 2617 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14943 2618 3133 2617 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14942 2617 3767 2618 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14941 2618 2741 2743 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14940 2743 6284 2618 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14939 4505 6860 4504 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14938 4504 4502 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14937 8552 4503 4505 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14936 4520 4505 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14935 2255 7326 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14934 2255 3677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14933 8552 3678 2255 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14932 3300 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14931 3300 3490 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14930 8552 5465 3300 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14929 8552 3171 2894 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14928 2997 2996 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14927 2894 2893 2996 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14926 2998 4577 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14925 2998 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14924 8552 2784 2998 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14923 6541 8237 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14922 6541 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14921 8552 6644 6541 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14920 4294 4292 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14919 8552 4320 4294 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14918 4518 4294 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14917 1733 2508 1693 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14916 8552 1956 1693 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14915 1693 3269 1733 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14914 1916 1733 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14913 6966 6964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14912 6966 7592 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14911 8552 8488 6966 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14910 8552 8240 6966 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14909 4697 4305 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14908 8552 8350 4697 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14907 6879 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14906 6879 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14905 8552 6717 6879 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14904 8552 8372 6879 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14903 75 77 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14902 78 3843 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14901 8552 983 79 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14900 8552 276 76 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14899 76 79 77 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14898 77 983 78 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14897 338 340 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14896 228 2718 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14895 8552 983 342 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14894 8552 992 227 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14893 227 342 340 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14892 340 983 228 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14891 8552 817 818 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14890 1180 818 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14889 8552 818 1180 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14888 8552 818 1180 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14887 1180 818 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14886 8552 1180 1181 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14885 6037 1181 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14884 8552 1181 6037 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14883 8552 1181 6037 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14882 6037 1181 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14881 8552 1180 1025 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14880 6285 1025 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14879 8552 1025 6285 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14878 8552 1025 6285 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14877 6285 1025 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14876 2180 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14875 2180 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14874 8552 3898 2180 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14873 8552 6021 2180 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14872 8552 8785 8786 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14871 8784 8786 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14870 8552 8786 8784 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14869 8552 8786 8784 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14868 8784 8786 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14867 8552 8784 8489 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14866 8488 8489 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14865 8552 8489 8488 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14864 8552 8489 8488 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14863 8488 8489 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14862 8552 8784 8491 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14861 8490 8491 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14860 8552 8491 8490 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14859 8552 8491 8490 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14858 8490 8491 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14857 5191 5841 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14856 8552 5196 5191 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14855 5189 5191 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14854 3183 3541 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14853 8552 3180 3183 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14852 3181 3183 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14851 7754 8220 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14850 8552 8455 7754 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14849 7752 7754 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14848 3970 3969 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14847 8552 4826 3970 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14846 3968 3970 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14845 6367 6370 6366 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14844 6366 6664 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14843 8552 7315 6367 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14842 6365 6367 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14841 8552 1021 1022 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14840 1022 4750 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14839 8552 2161 1022 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14838 1020 1022 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14837 8552 8098 8230 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14836 8230 8097 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14835 8230 8235 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14834 8552 8780 8230 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14833 8778 8230 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14832 8199 8690 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14831 4235 4371 4201 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14830 4200 4373 4235 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14829 8552 4233 4200 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14828 4233 4235 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14827 4367 4373 4233 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14826 8552 6361 4373 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14825 4371 4373 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14824 8552 4584 4372 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14823 4201 4372 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14822 4199 4198 4367 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14821 8552 4583 4199 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14820 4583 4367 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14819 8552 4367 4583 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14818 4468 4472 4471 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14817 8552 6934 4472 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14816 4470 4469 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14815 4471 6934 4470 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14814 8552 4473 4468 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14813 1929 1928 1824 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14812 1824 2511 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14811 8552 2936 1929 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14810 1926 1929 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14809 1915 3110 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14808 8552 1323 1915 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14807 3669 3676 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14806 3670 3672 3669 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14805 8552 3673 3670 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14804 8552 2344 1853 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14803 1853 1997 1998 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14802 5033 4350 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14801 4580 4358 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14800 8191 8703 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14799 5537 6115 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14798 5685 5683 5537 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14797 8552 5684 5685 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14796 8511 8632 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14795 8639 8630 8511 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14794 8552 8631 8639 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14793 1009 2986 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14792 7912 8778 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14791 8552 8030 7912 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14790 6447 8648 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14789 6447 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14788 8552 6272 6447 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14787 7097 7115 7098 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14786 7098 7118 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14785 8552 7660 7097 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14784 7096 7097 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14783 6548 6549 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14782 8552 7767 6548 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14781 8473 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14780 8552 8472 8473 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14779 5651 5655 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14778 5531 5660 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14777 8552 5656 5659 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14776 8552 6060 5530 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14775 5530 5659 5655 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14774 5655 5656 5531 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14773 601 599 600 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14772 600 608 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14771 8552 793 601 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14770 783 601 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14769 5557 8237 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14768 8552 7315 5557 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14767 1358 4532 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14766 8552 1552 1358 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14765 8694 8701 8531 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14764 8530 8702 8694 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14763 8552 8693 8530 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14762 8693 8694 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14761 8692 8702 8693 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14760 8552 8728 8702 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14759 8701 8702 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14758 8552 8696 8699 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14757 8531 8699 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14756 8529 8528 8692 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14755 8552 8690 8529 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14754 8690 8692 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14753 8552 8692 8690 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14752 6635 7660 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14751 6635 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14750 8552 7315 6635 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14749 6881 6879 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14748 8552 6878 6881 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14747 6882 6881 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14746 2782 2579 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14745 8552 2578 2782 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14744 7118 4027 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14743 8552 4533 7118 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14742 5864 5867 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14741 5868 8412 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14740 8552 6307 5869 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14739 8552 5865 5866 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14738 5866 5869 5867 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14737 5867 6307 5868 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14736 7301 7300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14735 8552 7304 7301 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14734 7532 7301 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14733 6347 6100 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14732 5954 6660 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14731 8552 8764 6101 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14730 8552 6339 5953 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14729 5953 6101 6100 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14728 6100 8764 5954 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14727 8763 8766 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14726 8550 8778 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14725 8552 8764 8767 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14724 8552 8761 8549 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14723 8549 8767 8766 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14722 8766 8764 8550 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14721 6424 6422 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14720 8552 6878 6424 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14719 6844 6424 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14718 8098 7979 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14717 7893 8168 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14716 8552 8430 7980 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14715 8552 8399 7894 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14714 7894 7980 7979 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14713 7979 8430 7893 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14712 5819 7273 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14711 5818 6007 5819 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14710 8552 6290 5818 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14709 5587 5415 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14708 5587 5790 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14707 8552 5466 5587 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14706 5890 7349 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14705 5890 6320 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14704 8552 5891 5890 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14703 8552 8478 5890 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14702 5032 5043 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14701 5031 5243 5032 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14700 8552 5041 5031 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14699 1069 4577 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14698 8552 2784 1069 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14697 1070 3531 1069 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14696 1069 1154 1070 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14695 1070 1157 3903 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14694 3903 6021 1070 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14693 5469 5470 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14692 5469 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14691 8552 6284 5469 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14690 8552 8350 5469 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14689 8552 5974 5975 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14688 5927 5974 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14687 6293 6433 5927 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14686 5927 5975 6293 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14685 8552 5971 5927 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14684 5971 6433 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14683 2350 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14682 2350 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14681 8552 5562 2350 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14680 8552 3333 2350 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14679 7688 7689 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14678 7622 8359 7689 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14677 7623 7880 7622 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14676 7624 7881 7623 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14675 8552 7877 7624 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14674 7615 7637 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14673 8049 7639 7615 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14672 8552 7636 8049 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14671 2112 2251 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14670 2481 2252 2112 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14669 8552 2260 2481 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14668 1018 3898 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14667 8552 6282 1018 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14666 1154 1018 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14665 8552 4279 4277 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14664 4178 4279 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14663 4281 4498 4178 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14662 4178 4277 4281 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14661 8552 4280 4178 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14660 4280 4498 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14659 8046 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14658 8248 8246 8046 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14657 8552 8247 8248 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14656 3002 6530 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14655 8552 5280 3002 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14654 3001 3002 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14653 8552 5137 4948 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14652 4946 5137 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14651 4947 6872 4946 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14650 4946 4948 4947 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14649 8552 4945 4946 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14648 4945 6872 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14647 7212 7307 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14646 7543 7308 7212 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14645 8552 8412 7543 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14644 4118 4115 4119 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14643 4117 4122 4118 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14642 8552 4116 4117 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14641 4116 4118 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14640 4114 4122 4116 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14639 8552 4121 4122 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14638 4115 4122 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14637 8552 4123 4120 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14636 4119 4120 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14635 4113 4112 4114 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14634 8552 8430 4113 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14633 8430 4114 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14632 8552 4114 8430 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14631 8552 3657 2217 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14630 2217 2648 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14629 2644 2482 2217 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14628 2216 3655 2644 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14627 2217 2639 2216 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14626 8552 6037 3949 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14625 3949 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14624 8552 6284 3949 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14623 3946 3949 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14622 8552 8235 6953 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14621 6953 8020 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14620 6953 7394 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14619 8552 8247 6953 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14618 6954 6953 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14617 8552 6284 5472 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14616 5472 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14615 5472 5470 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14614 8552 8350 5472 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14613 5891 5472 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14612 1394 1399 1397 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14611 1395 1400 1394 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14610 8552 1393 1395 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14609 1393 1394 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14608 1391 1400 1393 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14607 8552 2028 1400 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14606 1399 1400 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14605 8552 2593 1398 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14604 1397 1398 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14603 1392 1389 1391 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14602 8552 1390 1392 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14601 1390 1391 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14600 8552 1391 1390 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14599 1430 1476 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14598 1917 3273 1430 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14597 8552 1477 1917 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14596 8632 8358 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14595 8552 8627 8632 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14594 1845 2890 8552 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_14593 1996 4529 1845 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_14592 1844 1983 1996 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_14591 8552 3716 1844 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_14590 8552 5562 4998 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14589 4998 5563 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14588 8552 6716 4998 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14587 5446 4998 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14586 8552 6644 6529 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14585 6529 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14584 6529 7394 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14583 8552 8237 6529 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14582 6530 6529 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14581 8552 6037 1186 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14580 1186 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14579 1186 3898 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14578 8552 3531 1186 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14577 1372 1186 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14576 8552 6027 5525 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14575 5526 6290 5637 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14574 5527 6271 5526 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14573 5525 6022 5527 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14572 2297 2299 2207 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14571 2206 2300 2297 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14570 8552 2291 2206 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14569 2291 2297 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14568 2290 2300 2291 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14567 8552 3705 2300 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14566 2299 2300 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14565 8552 2293 2298 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14564 2207 2298 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14563 2205 2204 2290 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14562 8552 5188 2205 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14561 5188 2290 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14560 8552 2290 5188 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14559 4627 5263 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14558 5843 4750 4627 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14557 8552 4999 5843 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14556 4954 6246 4953 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14555 4953 5143 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14554 8552 4951 4954 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14553 4952 4954 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14552 4562 5870 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14551 4562 4339 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14550 8552 4338 4562 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14549 5400 5398 5403 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14548 5401 5405 5400 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14547 8552 5399 5401 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14546 5399 5400 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14545 5396 5405 5399 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14544 8552 6232 5405 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14543 5398 5405 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14542 8552 5402 5404 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14541 5403 5404 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14540 5397 5395 5396 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14539 8552 6251 5397 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14538 6251 5396 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14537 8552 5396 6251 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14536 2748 1546 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14535 8552 4027 2748 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14534 6125 6377 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14533 6125 7177 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14532 8552 6128 6125 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14531 1742 2277 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14530 8552 2937 1742 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14529 1741 1742 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14528 2151 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14527 2151 3898 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14526 8552 5013 2151 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14525 2571 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14524 2571 2983 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14523 8552 3295 2571 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14522 1976 1772 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14521 1976 1768 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14520 8552 4792 1976 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14519 2325 2760 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14518 2325 2328 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14517 8552 6307 2325 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14516 5178 5176 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14515 8552 5432 5178 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14514 5426 5178 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14513 6274 6287 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14512 8552 6878 6274 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14511 6273 6274 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14510 2508 8417 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14509 2508 3677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14508 8552 3678 2508 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14507 4154 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14506 4154 4111 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14505 8552 3960 4154 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14504 8552 3767 4154 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14503 6721 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14502 6721 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14501 8552 6717 6721 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14500 8552 8648 6721 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14499 6726 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14498 6726 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14497 8552 6286 6726 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14496 8552 6283 6726 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14495 3345 3639 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14494 3811 4469 3345 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14493 8552 8627 3811 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14492 1849 2890 8552 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_14491 1988 4530 1849 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_14490 1848 1987 1988 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_14489 8552 3717 1848 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_14488 8552 8349 8119 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14487 8119 8348 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14486 8119 8346 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14485 8552 8347 8119 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14484 8623 8119 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14483 8552 168 158 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14482 1760 158 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14481 8552 158 1760 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14480 8552 158 1760 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14479 1760 158 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14478 8552 1760 1761 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14477 6043 1761 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14476 8552 1761 6043 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14475 8552 1761 6043 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14474 6043 1761 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14473 8552 1760 1357 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14472 6286 1357 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14471 8552 1357 6286 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14470 8552 1357 6286 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14469 6286 1357 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14468 8552 1760 1528 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14467 6029 1528 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14466 8552 1528 6029 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14465 8552 1528 6029 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14464 6029 1528 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14463 8552 1760 157 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14462 6718 157 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14461 8552 157 6718 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14460 8552 157 6718 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14459 6718 157 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14458 3480 4327 3368 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14457 3368 6095 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14456 8552 3478 3480 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14455 3479 3480 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14454 6848 7049 6776 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14453 8552 6846 6776 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14452 6776 7643 6848 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14451 7252 6848 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14450 6260 6276 6261 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14449 6261 7311 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14448 8552 6711 6260 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14447 6259 6260 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14446 1801 2764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14445 8552 4300 1801 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14444 2016 1801 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14443 8552 3721 3719 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14442 3719 4103 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14441 8552 3884 3719 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14440 3718 3719 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14439 8552 6285 2547 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14438 2547 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14437 8552 3136 2547 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14436 2749 2547 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14435 737 746 656 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14434 655 745 737 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14433 8552 740 655 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14432 740 737 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14431 736 745 740 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14430 8552 1302 745 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14429 746 745 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14428 8552 944 744 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14427 656 744 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14426 654 653 736 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14425 8552 1105 654 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14424 1105 736 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14423 8552 736 1105 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14422 8552 8209 8015 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14421 8015 8782 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14420 8552 8780 8015 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14419 8478 8015 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14418 7547 7716 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14417 1369 1390 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14416 3136 1567 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14415 8552 5192 820 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14414 820 4111 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14413 820 5563 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14412 8552 4139 820 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14411 1030 820 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14410 5988 6250 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14409 5363 8433 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14408 6902 7126 6791 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14407 6791 7127 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14406 8552 8412 6902 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14405 6900 6902 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14404 7232 7239 7190 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14403 7189 7238 7232 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14402 8552 7231 7189 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14401 7231 7232 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14400 7230 7238 7231 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14399 8552 8596 7238 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14398 7239 7238 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14397 8552 7242 7237 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14396 7190 7237 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14395 7188 7187 7230 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14394 8552 7228 7188 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14393 7228 7230 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14392 8552 7230 7228 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14391 7873 8359 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14390 8362 8132 7873 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14389 8552 8131 8362 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14388 1138 5214 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14387 8552 1140 1138 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14386 8552 3150 2552 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14385 2551 2554 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14384 2552 2553 2554 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14383 943 5412 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14382 8552 1100 943 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14381 2760 2784 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14380 8552 6716 2760 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14379 5459 5462 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14378 5463 5460 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14377 8552 5461 5464 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14376 8552 5872 5458 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14375 5458 5464 5462 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14374 5462 5461 5463 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14373 8054 8056 7918 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14372 7919 8106 8054 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14371 8552 8052 7919 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14370 8052 8054 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14369 8102 8106 8052 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14368 8552 8596 8106 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14367 8056 8106 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14366 8552 8055 8108 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14365 7918 8108 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14364 7916 8032 8102 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14363 8552 8103 7916 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14362 8103 8102 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14361 8552 8102 8103 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14360 6473 6068 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14359 5941 6466 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14358 8552 6075 6069 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14357 8552 6303 5942 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14356 5942 6069 6068 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14355 6068 6075 5941 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14354 7317 8215 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14353 8552 7315 7317 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14352 7528 7317 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14351 6840 7065 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14350 8552 7066 6840 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14349 7246 6840 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14348 8552 6763 6706 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14347 7684 6706 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14346 8552 6706 7684 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14345 8552 6706 7684 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14344 7684 6706 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14343 8552 6763 6762 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14342 7765 6762 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14341 8552 6762 7765 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14340 8552 6762 7765 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14339 7765 6762 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14338 8552 4311 4312 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14337 6763 4312 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14336 8552 4312 6763 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14335 8552 4312 6763 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14334 6763 4312 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14333 5130 5415 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14332 5130 5139 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14331 8552 6022 5130 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14330 8552 3668 2919 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14329 2919 3106 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14328 8552 3657 2919 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14327 3247 2919 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14326 4346 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14325 4346 5465 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14324 8552 5471 4346 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14323 8552 8461 4346 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14322 2803 2783 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14321 2803 3180 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14320 8552 2587 2803 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14319 4628 4754 4755 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14318 4753 4751 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14317 8552 4753 4628 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14316 5607 5993 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14315 8552 5609 5607 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14314 5606 5607 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14313 5956 6115 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14312 6358 6364 5956 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14311 8552 6109 6358 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14310 3111 5408 3025 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14309 3025 6288 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14308 8552 5631 3111 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14307 3110 3111 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14306 619 1390 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14305 8552 2566 619 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14304 817 619 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14303 6748 6746 6653 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14302 6651 6751 6748 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14301 8552 6747 6651 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14300 6747 6748 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14299 6744 6751 6747 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14298 8552 8728 6751 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14297 6746 6751 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14296 8552 6919 6749 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14295 6653 6749 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14294 6650 6745 6744 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14293 8552 6920 6650 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14292 6920 6744 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14291 8552 6744 6920 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14290 8552 3121 3124 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14289 3124 3125 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14288 8552 3120 3124 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14287 3280 3124 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14286 3264 3262 3263 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14285 3263 3271 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14284 8552 3261 3264 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14283 3392 3264 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14282 2513 2940 2512 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14281 8552 2942 2512 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14280 2512 3479 2513 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14279 2511 2513 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14278 8024 8246 7909 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14277 7909 8098 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14276 8552 8247 8024 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14275 7908 8024 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14274 8552 8483 6114 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14273 6114 6644 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14272 8552 8237 6114 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14271 6111 6114 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14270 4555 4759 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14269 4554 7315 4555 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14268 8552 4553 4554 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14267 5569 5693 5504 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14266 5501 5692 5569 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14265 8552 5568 5501 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14264 5568 5569 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14263 5687 5692 5568 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14262 8552 6361 5692 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14261 5693 5692 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14260 8552 5910 5691 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14259 5504 5691 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14258 5497 5538 5687 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14257 8552 5907 5497 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14256 5907 5687 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14255 8552 5687 5907 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14254 5922 6674 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14253 8552 6378 5922 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14252 8552 5046 1580 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14251 1580 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14250 1580 3753 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14249 8552 3490 1580 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14248 1791 1580 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14247 7090 7096 7091 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14246 7089 7087 7090 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14245 8552 7088 7089 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14244 3414 2949 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14243 8552 5676 3414 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14242 2226 2273 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14241 2938 2274 2226 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14240 8552 2723 2938 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14239 4462 4466 4461 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14238 4463 4467 4462 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14237 8552 4460 4463 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14236 4460 4462 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14235 4459 4467 4460 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14234 8552 6232 4467 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14233 4466 4467 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14232 8552 4464 4465 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14231 4461 4465 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14230 4457 4458 4459 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14229 8552 6022 4457 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14228 6022 4459 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14227 8552 4459 6022 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14226 7874 7957 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14225 8552 8369 7874 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14224 3526 3519 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14223 8552 3318 3526 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14222 983 2734 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14221 8552 1129 983 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14220 2928 2933 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14219 8552 2927 2928 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14218 2926 2928 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14217 3417 5580 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_14216 3420 3482 3354 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14215 3354 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14214 8552 3412 3356 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14213 3356 3415 3355 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14212 3355 3417 3420 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14211 3420 5580 3357 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14210 8552 3414 3412 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_14209 3411 3420 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14208 3357 3671 3356 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14207 2655 3066 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_14206 2657 3660 2597 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14205 2597 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14204 8552 2652 2599 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14203 2599 2659 2598 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14202 2598 2655 2657 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14201 2657 3066 2600 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14200 8552 3414 2652 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_14199 3646 2657 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14198 2600 3665 2599 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14197 8552 3677 3679 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14196 3679 3678 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14195 8552 7142 3679 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14194 3676 3679 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14193 1064 1113 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14192 1116 1114 1064 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14191 8552 2723 1116 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14190 3978 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14189 3978 4111 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14188 8552 5046 3978 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14187 8552 3964 3978 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14186 8552 8383 7887 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14185 8552 8627 7964 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14184 7887 7964 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14183 6766 8240 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14182 6766 6954 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14181 8552 8490 6766 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14180 2761 2760 2627 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14179 2627 2890 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14178 8552 2763 2761 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14177 2847 2761 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14176 8552 632 630 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14175 831 630 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14174 8552 630 831 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14173 8552 630 831 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14172 831 630 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14171 8552 831 830 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14170 6040 830 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14169 8552 830 6040 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14168 8552 830 6040 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14167 6040 830 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14166 8552 831 627 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14165 6717 627 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14164 8552 627 6717 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14163 8552 627 6717 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14162 6717 627 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14161 8552 831 832 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14160 6282 832 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14159 8552 832 6282 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14158 8552 832 6282 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14157 6282 832 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14156 3325 3311 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14155 3308 3307 3311 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14154 3309 3759 3308 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14153 8552 3310 3309 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14152 8552 2160 2162 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14151 2162 2161 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14150 8552 6077 2162 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14149 4127 2162 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14148 7690 7502 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14147 7503 7933 7502 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14146 7500 7880 7503 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14145 7501 7881 7500 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14144 8552 7499 7501 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14143 8552 836 837 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14142 835 837 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14141 8552 837 835 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14140 8552 837 835 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14139 835 837 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14138 8552 835 833 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14137 3960 833 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14136 8552 833 3960 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14135 8552 833 3960 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14134 3960 833 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14133 8552 835 834 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14132 5046 834 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14131 8552 834 5046 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14130 8552 834 5046 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14129 5046 834 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14128 2177 2571 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14127 8552 2176 2177 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14126 2354 2177 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14125 2577 2579 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14124 8552 2578 2577 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14123 2999 2577 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14122 8552 8236 7406 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14121 7406 8246 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14120 8552 8237 7406 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14119 7404 7406 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14118 8552 8634 8631 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14117 8552 8627 8629 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14116 8631 8629 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14115 8552 2764 1198 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14114 1198 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14113 8552 4139 1198 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14112 1381 1198 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14111 8722 8729 8539 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14110 8538 8730 8722 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14109 8552 8720 8538 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14108 8720 8722 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14107 8719 8730 8720 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14106 8552 8728 8730 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14105 8729 8730 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14104 8552 8723 8727 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14103 8539 8727 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14102 8537 8536 8719 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14101 8552 8717 8537 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14100 8717 8719 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14099 8552 8719 8717 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14098 6247 6000 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14097 5613 6246 5519 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14096 5519 5612 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14095 8552 7495 5613 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14094 5611 5613 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14093 5102 6072 5246 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14092 5101 6758 5102 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14091 8552 8717 5101 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14090 4805 4810 4639 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14089 4638 4809 4805 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14088 8552 4802 4638 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14087 4802 4805 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14086 4801 4809 4802 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14085 8552 6361 4809 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14084 4810 4809 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14083 8552 5035 4808 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14082 4639 4808 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14081 4637 4636 4801 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14080 8552 5036 4637 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14079 5036 4801 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14078 8552 4801 5036 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14077 8552 4577 1605 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14076 1605 3898 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14075 1605 5013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14074 8552 4139 1605 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14073 1602 1605 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14072 8359 8634 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14071 7277 7947 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14070 5436 5188 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14069 792 4027 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14068 8552 2159 792 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14067 3799 3897 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14066 3880 7115 3799 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14065 8552 6022 3880 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14064 4557 4751 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14063 4778 4789 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14062 8552 4562 4778 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14061 3824 3831 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14060 3831 3827 3792 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14059 8552 3832 3792 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14058 3792 3828 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14057 3791 3825 3831 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14056 3792 3826 3791 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14055 1118 4700 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14054 8552 1116 1118 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14053 3326 6530 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14052 8552 5280 3326 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14051 8710 8714 8534 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14050 8535 8715 8710 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14049 8552 8706 8535 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14048 8706 8710 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14047 8705 8715 8706 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14046 8552 8728 8715 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14045 8714 8715 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14044 8552 8711 8713 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14043 8534 8713 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14042 8533 8532 8705 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14041 8552 8703 8533 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14040 8703 8705 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14039 8552 8705 8703 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14038 3478 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14037 3478 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14036 8552 6282 3478 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14035 8552 3750 3478 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14034 3288 4750 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14033 8552 4529 3288 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14032 5341 5189 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14031 8552 5186 5341 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14030 6515 6517 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14029 6392 6936 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14028 8552 8764 6519 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14027 8552 6514 6393 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14026 6393 6519 6517 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14025 6517 8764 6392 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14024 8552 3479 2941 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14023 2941 3083 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14022 8552 2940 2941 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14021 3657 2941 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14020 6663 7749 6664 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14019 6767 7173 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14018 8552 6767 6663 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14017 5677 5680 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14016 5536 5895 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14015 8552 7347 5681 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14014 8552 5676 5535 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14013 5535 5681 5680 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14012 5680 7347 5536 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14011 7544 7542 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14010 8552 7543 7544 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14009 7932 7544 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14008 2967 2965 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14007 2964 2966 2967 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14006 8552 8731 2964 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14005 4750 4577 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14004 4750 3898 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14003 8552 6282 4750 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14002 1841 1977 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14001 3315 1978 1841 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14000 8552 7535 3315 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13999 8552 1373 1375 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13998 1783 1376 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13997 1375 1374 1376 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13996 8552 1030 1033 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13995 1995 1032 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13994 1033 1031 1032 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13993 6927 6929 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13992 6754 7573 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13991 8552 8764 6930 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13990 8552 6925 6753 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13989 6753 6930 6929 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13988 6929 8764 6754 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13987 8552 2272 2135 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13986 2134 2272 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13985 2517 2133 2134 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13984 2134 2135 2517 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13983 8552 2132 2134 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13982 2132 2133 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13981 8552 7251 7250 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13980 7250 7481 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13979 7250 7252 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13978 8552 7246 7250 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13977 8326 7250 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13976 1993 3318 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13975 8552 1992 1993 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13974 2000 1993 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13973 3130 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13972 8552 6718 3130 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13971 3294 3130 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13970 119 121 118 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13969 120 123 119 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13968 8552 117 120 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13967 117 119 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13966 115 123 117 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13965 8552 1516 123 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13964 121 123 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13963 8552 313 122 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13962 118 122 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13961 114 113 115 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13960 8552 554 114 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13959 554 115 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13958 8552 115 554 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13957 8552 4751 4187 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13956 4187 4747 4318 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13955 8552 2981 2186 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13954 2186 3335 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13953 8552 2185 2186 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13952 2374 2186 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13951 8552 8781 8016 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13950 8016 8450 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13949 8552 8237 8016 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13948 8030 8016 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13947 5821 6246 5820 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13946 5820 6006 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13945 8552 6428 5821 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13944 5822 5821 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13943 795 604 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13942 604 602 605 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13941 8552 3295 605 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13940 605 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13939 603 1009 604 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13938 605 5192 603 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13937 4731 4735 4622 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13936 4621 4737 4731 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13935 8552 4729 4621 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13934 4729 4731 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13933 4728 4737 4729 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13932 8552 5835 4737 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13931 4735 4737 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13930 8552 7142 4736 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13929 4622 4736 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13928 4620 4619 4728 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13927 8552 4727 4620 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13926 4727 4728 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13925 8552 4728 4727 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13924 8552 8223 8017 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13923 8017 8222 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13922 8552 8780 8017 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13921 8240 8017 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13920 7225 7400 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13919 8552 7579 7225 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13918 7226 7593 7225 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13917 7225 7756 7226 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13916 7226 7379 7381 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13915 7381 8023 7226 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13914 269 271 206 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13913 207 273 269 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13912 8552 265 207 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13911 265 269 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13910 264 273 265 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13909 8552 1302 273 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13908 271 273 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13907 8552 517 272 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13906 206 272 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13905 205 235 264 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13904 8552 720 205 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13903 720 264 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13902 8552 264 720 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13901 7094 7092 7279 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13900 7095 7093 7094 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13899 8552 7102 7095 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13898 3733 3736 3732 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13897 3734 3738 3733 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13896 8552 3731 3734 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13895 3731 3733 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13894 3730 3738 3731 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13893 8552 4121 3738 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13892 3736 3738 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13891 8552 3735 3737 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13890 3732 3737 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13889 3729 3728 3730 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13888 8552 3750 3729 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13887 3750 3730 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13886 8552 3730 3750 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13885 7180 8098 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13884 7184 8246 7180 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13883 8552 8247 7184 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13882 8617 7091 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13881 8552 7275 8617 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13880 5216 6077 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13879 5216 6307 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13878 8552 4999 5216 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13877 2156 2328 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13876 8552 4533 2156 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13875 2155 2156 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13874 388 4350 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13873 388 805 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13872 8552 2974 388 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13871 2960 2961 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13870 2960 3956 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13869 8552 3964 2960 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13868 2507 2949 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13867 8552 5676 2507 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13866 3261 2507 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13865 616 5033 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13864 616 805 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13863 8552 2974 616 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13862 613 807 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13861 613 2976 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13860 8552 391 613 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13859 4772 5011 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13858 8552 5231 4772 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13857 5215 4772 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13856 4302 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13855 4302 6037 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13854 8552 6029 4302 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13853 8552 5440 4302 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13852 8552 4750 1970 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13851 1970 4027 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13850 1970 4529 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13849 8552 2159 1970 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13848 2153 1970 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13847 161 7536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13846 160 1016 162 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13845 360 162 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13844 162 369 161 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13843 8552 1015 160 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13842 5823 5822 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13841 8552 6008 5823 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13840 5824 5823 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13839 7207 7307 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13838 7291 7308 7207 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13837 8552 7723 7291 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13836 8552 2644 2643 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13835 2606 2644 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13834 2904 2639 2606 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13833 2606 2643 2904 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13832 8552 2640 2606 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13831 2640 2639 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13830 935 941 939 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13829 936 940 935 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13828 8552 934 936 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13827 934 935 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13826 933 940 934 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13825 8552 1302 940 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13824 941 940 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13823 8552 937 938 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13822 939 938 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13821 932 930 933 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13820 8552 931 932 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13819 931 933 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13818 8552 933 931 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13817 8552 6718 4578 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13816 4578 4577 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13815 8552 5563 4578 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13814 5043 4578 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13813 8552 3490 407 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13812 407 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13811 407 5465 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13810 8552 4300 407 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13809 498 407 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13808 7069 7472 7070 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13807 8552 7068 7070 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13806 7070 7643 7069 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13805 7481 7069 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13804 914 918 917 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13803 915 919 914 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13802 8552 913 915 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13801 913 914 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13800 911 919 913 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13799 8552 1302 919 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13798 918 919 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13797 8552 920 916 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13796 917 916 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13795 912 910 911 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13794 8552 1092 912 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13793 1092 911 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13792 8552 911 1092 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13791 4102 4529 4041 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13790 8552 8128 4041 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13789 4041 4530 4102 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13788 4103 4102 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13787 7879 8586 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13786 7933 8110 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13785 6095 5220 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13784 4133 5790 4132 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13783 4131 8731 4133 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13782 8552 5036 4131 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13781 4339 4564 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13780 8552 4342 4339 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13779 3650 3396 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13778 3650 3392 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13777 8552 3824 3650 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13776 2506 2504 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13775 3872 2505 2506 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13774 8552 2723 3872 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13773 4616 5440 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13772 8552 5843 4616 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13771 4617 4715 4616 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13770 4616 5844 4617 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13769 4617 4710 4712 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13768 4712 8103 4617 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13767 2145 6324 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13766 5817 8572 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13765 5518 7880 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13764 5609 6007 5518 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13763 8552 6022 5609 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13762 8552 5166 4618 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13761 4718 4719 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13760 4618 4717 4719 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13759 6682 6684 6622 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13758 6623 6687 6682 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13757 8552 6685 6623 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13756 6685 6682 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13755 6681 6687 6685 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13754 8552 8596 6687 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13753 6684 6687 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13752 8552 6688 6686 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13751 6622 6686 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13750 6620 6683 6681 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13749 8552 6708 6620 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13748 6708 6681 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13747 8552 6681 6708 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13746 1477 1318 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13745 8552 1496 1477 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13744 1876 5624 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13743 8552 1753 1876 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13742 5909 6115 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13741 5910 5911 5909 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13740 8552 5908 5910 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13739 7177 7178 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13738 8552 7582 7177 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13737 6138 5634 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13736 8552 5551 6138 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13735 6728 8160 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13734 6728 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13733 8552 7315 6728 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13732 1748 2138 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13731 1752 1755 1745 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13730 1745 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13729 8552 1746 1751 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13728 1751 1747 1749 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13727 1749 1748 1752 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13726 1752 2138 1750 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13725 8552 3414 1746 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13724 2133 1752 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13723 1750 1945 1751 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13722 3085 3082 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13721 3085 3668 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13720 8552 3106 3085 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13719 8552 3083 3085 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13718 3022 3832 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13717 3395 3655 3022 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13716 8552 3654 3395 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13715 5209 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13714 5209 5013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13713 8552 5465 5209 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13712 8552 6514 5209 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13711 5439 5438 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13710 8552 5557 5439 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13709 8132 5439 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13708 3653 4662 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13707 3652 4258 3653 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13706 8552 4064 3652 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13705 8552 3490 3436 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13704 3436 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13703 3436 6026 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13702 8552 8572 3436 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13701 3685 3436 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13700 5930 5984 7311 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13699 8552 8065 5984 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13698 5931 6691 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13697 7311 8065 5931 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13696 8552 6234 5930 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13695 7770 7184 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13694 7770 7593 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13693 8552 8030 7770 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13692 8552 8240 7770 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13691 7392 7391 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13690 8552 8487 7392 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13689 8026 7392 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13688 8552 4320 4183 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13687 4183 4292 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13686 5166 4520 4183 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13685 4182 4289 5166 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13684 4183 5169 4182 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13683 2973 2972 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13682 8552 3509 2973 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13681 2978 2973 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13680 8552 4747 4539 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13679 8552 4758 4540 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13678 4539 4540 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13677 7157 7163 7160 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13676 7158 7162 7157 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13675 8552 7156 7158 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13674 7156 7157 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13673 7154 7162 7156 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13672 8552 8728 7162 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13671 7163 7162 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13670 8552 7159 7161 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13669 7160 7161 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13668 7155 7152 7154 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13667 8552 7153 7155 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13666 7153 7154 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13665 8552 7154 7153 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13664 1487 2277 1431 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13663 1431 2937 1487 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13662 8552 1956 1431 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13661 8552 6286 3169 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13660 3169 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13659 3169 3767 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13658 8552 3333 3169 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13657 3171 3169 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13656 8552 8235 7396 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13655 7396 8236 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13654 7396 7394 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13653 8552 8237 7396 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13652 8027 7396 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13651 7486 8553 7487 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13650 8552 7485 7487 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13649 7487 7643 7486 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13648 8325 7486 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13647 6785 6816 7686 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13646 6784 6874 6785 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13645 8552 6893 6784 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13644 4205 4243 4163 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13643 4162 4244 4205 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13642 8552 4203 4162 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13641 4203 4205 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13640 4238 4244 4203 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13639 8552 6232 4244 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13638 4243 4244 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13637 8552 4206 4242 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13636 4163 4242 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13635 4161 4160 4238 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13634 8552 5790 4161 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13633 5790 4238 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13632 8552 4238 5790 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13631 4816 4820 4643 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13630 4642 4821 4816 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13629 8552 4813 4642 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13628 4813 4816 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13627 4811 4821 4813 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13626 8552 6361 4821 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13625 4820 4821 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13624 8552 5267 4819 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13623 4643 4819 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13622 4641 4640 4811 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13621 8552 5263 4641 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13620 5263 4811 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13619 8552 4811 5263 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13618 4629 5010 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13617 4773 5893 4629 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13616 8552 5014 4773 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13615 8552 3551 3010 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13614 3013 3341 3012 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13613 3014 3011 3013 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13612 3010 3544 3014 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13611 2222 2505 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13610 2501 2504 2222 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13609 8552 2260 2501 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13608 2936 2940 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13607 2936 3479 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13606 8552 3083 2936 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13605 7680 7283 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13604 8552 7282 7680 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13603 6668 6673 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13602 8552 8490 6668 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13601 8646 7279 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13600 8552 7280 8646 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13599 8116 8069 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13598 8552 8350 8116 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13597 5798 5801 5797 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13596 5799 5802 5798 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13595 8552 5796 5799 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13594 5796 5798 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13593 5795 5802 5796 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13592 8552 6232 5802 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13591 5801 5802 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13590 8552 5976 5800 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13589 5797 5800 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13588 5793 5794 5795 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13587 8552 6311 5793 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13586 6311 5795 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13585 8552 5795 6311 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13584 2516 2515 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13583 2699 2518 2516 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13582 8552 2706 2699 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13581 2664 3254 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13580 2664 3092 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13579 8552 3102 2664 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13578 2965 2955 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13577 2955 6021 2956 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13576 8552 3531 2956 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13575 2956 3297 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13574 2954 3295 2955 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13573 2956 3137 2954 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13572 3544 3968 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13571 8552 3973 3544 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13570 7356 7592 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13569 7356 7576 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13568 8552 7353 7356 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13567 5966 5584 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13566 5514 5580 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13565 8552 6934 5585 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13564 8552 5958 5513 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13563 5513 5585 5584 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13562 5584 6934 5514 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13561 5543 5372 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13560 5373 5371 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13559 8552 6934 5374 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13558 8552 6271 5370 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13557 5370 5374 5372 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13556 5372 6934 5373 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13555 3092 8168 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13554 3092 3677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13553 8552 3678 3092 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13552 2921 3668 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13551 8552 3106 2921 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13550 3073 2921 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13549 8552 3478 2946 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13548 2946 3471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13547 8552 3885 2946 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13546 2945 2946 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13545 3520 3762 3376 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13544 3376 6092 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13543 8552 3761 3520 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13542 3519 3520 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13541 7170 8478 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13540 7170 7373 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13539 8552 7169 7170 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13538 7298 7297 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13537 8552 7305 7298 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13536 7657 7298 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13535 4464 4246 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13534 4165 4247 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13533 8552 6934 4248 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13532 8552 6022 4164 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13531 4164 4248 4246 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13530 4246 6934 4165 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13529 612 4358 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13528 612 805 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13527 8552 2974 612 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13526 6662 6964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13525 6662 7391 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13524 8552 8030 6662 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13523 6238 6234 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13522 8552 8065 6238 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13521 4099 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13520 4099 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13519 8552 6282 4099 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13518 8552 4522 4099 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13517 6242 6410 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13516 8552 8065 6242 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13515 5811 7880 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13514 5989 6007 5811 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13513 8552 6311 5989 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13512 7280 7278 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13511 7206 7521 7278 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13510 7204 7880 7206 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13509 7205 7881 7204 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13508 8552 7877 7205 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13507 2144 4529 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13506 8552 4530 2144 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13505 2532 2144 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13504 5812 5814 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13503 5815 5817 5814 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13502 5816 7273 5815 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13501 5813 7881 5816 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13500 8552 7877 5813 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13499 4691 4949 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13498 8552 4955 4691 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13497 4690 4691 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13496 8552 4928 4930 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13495 4930 4929 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13494 8552 5415 4930 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13493 4927 4930 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13492 8552 8098 7372 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13491 7372 7394 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13490 8552 8247 7372 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13489 7592 7372 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13488 6507 6511 6390 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13487 6391 6513 6507 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13486 8552 6504 6391 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13485 6504 6507 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13484 6502 6513 6504 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13483 8552 6512 6513 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13482 6511 6513 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13481 8552 6655 6510 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13480 6390 6510 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13479 6389 6405 6502 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13478 8552 6758 6389 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13477 6758 6502 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13476 8552 6502 6758 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13475 942 1462 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13474 1308 1463 942 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13473 8552 2260 1308 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13472 5810 7049 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13471 8552 6285 1036 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13470 1036 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13469 1036 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13468 8552 6021 1036 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13467 1189 1036 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13466 6345 6349 6344 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13465 6346 6350 6345 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13464 8552 6343 6346 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13463 6343 6345 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13462 6342 6350 6343 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13461 8552 6361 6350 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13460 6349 6350 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13459 8552 6347 6348 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13458 6344 6348 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13457 6341 6340 6342 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13456 8552 6339 6341 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13455 6339 6342 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13454 8552 6342 6339 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13453 5174 5826 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13452 4799 5498 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13451 6654 7153 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13450 6426 6251 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13449 6426 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13448 8552 7315 6426 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13447 2939 4286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13446 8552 2938 2939 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13445 6433 6271 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13444 6257 6005 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13443 6257 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13442 8552 7315 6257 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13441 2943 2949 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13440 8552 6925 2943 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13439 2942 2943 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13438 8018 8098 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13437 8552 8247 8018 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13436 5889 5888 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13435 8552 5892 5889 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13434 793 791 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13433 669 802 791 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13432 670 794 669 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13431 671 795 670 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13430 8552 792 671 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13429 684 4027 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13428 8552 1363 684 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13427 7560 7325 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13426 7218 7326 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13425 8552 8423 7328 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13424 8552 7553 7217 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13423 7217 7328 7325 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13422 7325 8423 7218 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13421 8404 8171 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13420 7981 8168 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13419 8552 8423 8172 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13418 8552 8399 7982 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13417 7982 8172 8171 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13416 8171 8423 7981 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13415 7135 6905 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13414 6731 7142 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13413 8552 8423 6906 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13412 8552 7140 6732 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13411 6732 6906 6905 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13410 6905 8423 6731 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13409 3106 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13408 3106 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13407 8552 3490 3106 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13406 8552 8572 3106 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13405 7101 7307 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13404 7282 7308 7101 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13403 8552 7718 7282 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13402 5109 6115 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13401 5292 5914 5109 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13400 8552 5275 5292 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13399 8684 8413 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13398 8414 8412 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13397 8552 8423 8415 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13396 8552 8677 8411 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13395 8411 8415 8413 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13394 8413 8423 8414 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13393 8781 8181 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13392 7994 8412 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13391 8552 8430 8183 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13390 8552 8677 7990 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13389 7990 8183 8181 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13388 8181 8430 7994 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13387 8552 6878 4989 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13386 4989 4988 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13385 8552 6077 4989 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13384 4987 4989 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13383 2772 1999 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13382 2772 2172 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13381 8552 1998 2772 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13380 8552 2000 2772 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13379 8552 4527 4528 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13378 4525 4527 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13377 4526 6279 4525 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13376 4525 4528 4526 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13375 8552 4524 4525 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13374 4524 6279 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13373 3272 6288 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13372 3273 5408 3272 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13371 8552 5631 3273 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13370 7142 6735 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13369 8552 2569 2568 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13368 2568 2570 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13367 8552 2756 2568 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13366 2567 2568 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13365 575 576 574 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13364 573 578 575 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13363 8552 572 573 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13362 572 575 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13361 571 578 572 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13360 8552 1516 578 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13359 576 578 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13358 8552 980 577 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13357 574 577 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13356 570 569 571 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13355 8552 1124 570 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13354 1124 571 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13353 8552 571 1124 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13352 5099 6514 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13351 5656 5218 5099 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13350 8552 5216 5656 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13349 6809 6810 6703 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13348 6704 6855 6809 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13347 8552 6807 6704 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13346 6807 6809 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13345 6851 6855 6807 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13344 8552 8596 6855 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13343 6810 6855 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13342 8552 8168 6857 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13341 6703 6857 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13340 6702 6778 6851 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13339 8552 6852 6702 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13338 6852 6851 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13337 8552 6851 6852 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13336 8552 1558 804 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13335 804 1020 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13334 804 1769 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13333 8552 6077 804 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13332 805 804 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13331 4572 4575 4571 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13330 4570 4576 4572 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13329 8552 4569 4570 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13328 4569 4572 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13327 4567 4576 4569 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13326 8552 6361 4576 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13325 4575 4576 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13324 8552 4573 4574 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13323 4571 4574 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13322 4568 4566 4567 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13321 8552 4754 4568 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13320 4754 4567 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13319 8552 4567 4754 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13318 152 154 151 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13317 153 156 152 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13316 8552 150 153 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13315 150 152 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13314 148 156 150 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13313 8552 1516 156 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13312 154 156 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13311 8552 338 155 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13310 151 155 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13309 147 146 148 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13308 8552 992 147 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13307 992 148 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13306 8552 148 992 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13305 4188 4799 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13304 4328 4327 4188 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13303 8552 4334 4328 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13302 6289 6288 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13301 6821 6873 6289 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13300 8552 6287 6821 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13299 5987 6246 5932 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13298 5932 5988 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13297 8552 6235 5987 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13296 5985 5987 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13295 8665 7686 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13294 8552 7688 8665 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13293 4781 4785 4632 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13292 4633 4786 4781 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13291 8552 4777 4633 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13290 4777 4781 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13289 4776 4786 4777 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13288 8552 6512 4786 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13287 4785 4786 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13286 8552 4778 4784 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13285 4632 4784 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13284 4631 4630 4776 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13283 8552 5870 4631 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13282 5870 4776 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13281 8552 4776 5870 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13280 3551 4153 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13279 8552 3979 3551 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13278 5976 5980 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13277 5929 5978 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13276 8552 6934 5981 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13275 8552 6311 5928 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13274 5928 5981 5980 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13273 5980 6934 5929 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13272 2113 2247 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13271 3838 2248 2113 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13270 8552 2260 3838 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13269 8353 8623 8354 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13268 8354 8625 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13267 8552 8627 8353 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13266 8622 8353 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13265 4673 4260 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13264 4171 4258 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13263 8552 6934 4261 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13262 8552 6283 4170 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13261 4170 4261 4260 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13260 4260 6934 4171 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13259 8552 3285 3284 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13258 3460 3283 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13257 3284 3282 3283 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13256 1021 1009 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13255 1021 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13254 8552 5471 1021 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13253 7171 7173 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13252 7171 7593 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13251 8552 8490 7171 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13250 3828 2916 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13249 2916 3654 2917 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13248 8552 3657 2917 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13247 2917 3658 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13246 2915 3832 2916 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13245 2917 3655 2915 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13244 167 5470 168 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13243 166 1203 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13242 8552 166 167 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13241 8453 8474 8452 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13240 8552 8764 8452 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13239 8452 8459 8453 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13238 8451 8453 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13237 8552 6316 5865 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13236 8552 6283 5855 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13235 5865 5855 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13234 8552 6307 2158 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13233 2158 2337 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13232 2158 2760 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13231 8552 2161 2158 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13230 2157 2158 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13229 1722 2255 1721 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13228 1721 2127 1722 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13227 8552 1956 1721 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13226 6634 6843 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13225 7093 6873 6634 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13224 8552 6711 7093 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13223 1106 5214 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13222 8552 1105 1106 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13221 2505 1106 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13220 8601 8603 8505 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13219 8552 8599 8505 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13218 8505 8602 8601 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13217 8600 8601 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13216 301 304 214 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13215 215 306 301 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13214 8552 298 215 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13213 298 301 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13212 297 306 298 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13211 8552 1516 306 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13210 304 306 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13209 8552 550 305 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13208 214 305 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13207 213 239 297 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13206 8552 548 213 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13205 548 297 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13204 8552 297 548 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13203 8552 6373 6375 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13202 6375 6374 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13201 6375 6666 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13200 8552 6376 6375 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13199 6372 6375 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13198 8552 3753 825 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13197 825 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13196 825 3490 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13195 8552 5465 825 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13194 827 825 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13193 8552 6717 3917 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13192 3917 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13191 8552 5562 3917 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13190 3915 3917 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13189 6318 8000 6319 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13188 6317 7345 6318 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13187 8552 6316 6317 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13186 8318 8350 8567 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13185 8317 8572 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13184 8552 8317 8318 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13183 1350 1355 1353 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13182 1351 1356 1350 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13181 8552 1349 1351 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13180 1349 1350 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13179 1347 1356 1349 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13178 8552 1367 1356 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13177 1355 1356 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13176 8552 1521 1354 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13175 1353 1354 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13174 1348 1346 1347 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13173 8552 1522 1348 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13172 1522 1347 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13171 8552 1347 1522 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13170 1913 2128 1819 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13169 1819 1924 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13168 8552 1910 1913 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13167 1911 1913 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13166 8552 3433 2126 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13165 2498 2125 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13164 2126 2124 2125 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13163 6720 6311 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13162 6872 6022 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13161 6843 6290 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13160 8652 8659 8519 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13159 8518 8660 8652 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13158 8552 8651 8518 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13157 8651 8652 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13156 8650 8660 8651 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13155 8552 8674 8660 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13154 8659 8660 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13153 8552 8655 8658 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13152 8519 8658 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13151 8517 8516 8650 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13150 8552 8648 8517 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13149 8648 8650 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13148 8552 8650 8648 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13147 8552 1995 1787 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13146 1788 1790 2182 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13145 1789 1996 1788 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13144 1787 1791 1789 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13143 6279 6283 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13142 4473 4943 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13141 8552 1372 1071 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13140 1072 1193 2346 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13139 1073 1189 1072 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13138 1071 1373 1073 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13137 4511 4514 4510 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13136 4512 4515 4511 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13135 8552 4509 4512 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13134 4509 4511 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13133 4508 4515 4509 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13132 8552 5835 4515 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13131 4514 4515 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13130 8552 4516 4513 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13129 4510 4513 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13128 4507 4506 4508 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13127 8552 4715 4507 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13126 4715 4508 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13125 8552 4508 4715 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13124 7126 3140 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13123 3140 3745 3034 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13122 8552 3137 3034 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13121 3034 3136 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13120 3033 3531 3140 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13119 3034 3753 3033 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13118 1977 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13117 8552 3956 1977 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13116 4792 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13115 4792 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13114 8552 6285 4792 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13113 4541 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13112 4541 4111 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13111 8552 6282 4541 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13110 2220 2252 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13109 5551 2251 2220 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13108 8552 2723 5551 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13107 2305 3767 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13106 2305 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13105 8552 6282 2305 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13104 8711 8422 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13103 8424 8427 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13102 8552 8423 8425 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13101 8552 8703 8421 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13100 8421 8425 8422 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13099 8422 8423 8424 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13098 4100 4099 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13097 8552 6878 4100 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13096 4295 4100 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13095 8552 3657 2611 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13094 2611 2926 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13093 2672 2675 2611 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13092 2610 3655 2672 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13091 2611 2671 2610 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13090 8209 8174 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13089 7985 8175 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13088 8552 8430 8177 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13087 8552 8410 7983 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13086 7983 8177 8174 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13085 8174 8430 7985 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13084 8782 8429 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13083 8428 8427 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13082 8552 8430 8431 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13081 8552 8703 8426 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13080 8426 8431 8429 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13079 8429 8430 8428 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13078 636 3158 638 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13077 637 8350 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13076 8552 637 636 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13075 4579 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13074 4579 5465 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13073 8552 5563 4579 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13072 8552 8065 4579 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13071 1486 1755 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13070 1484 1915 1409 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13069 1409 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13068 8552 1480 1412 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13067 1412 1479 1410 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13066 1410 1486 1484 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13065 1484 1755 1411 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13064 8552 3414 1480 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13063 1737 1484 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13062 1411 1487 1412 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13061 8223 8203 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13060 8012 8202 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13059 8552 8430 8204 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13058 8552 8199 8011 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13057 8011 8204 8203 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13056 8203 8430 8012 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13055 3287 3285 3462 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13054 3286 3463 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13053 8552 3286 3287 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13052 8316 8315 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13051 8561 8321 8316 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13050 8552 8314 8561 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13049 8552 2904 2902 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13048 2905 2904 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13047 4247 2911 2905 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13046 2905 2902 4247 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13045 8552 2903 2905 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13044 2903 2911 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13043 1914 1919 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13042 1919 1917 1821 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13041 8552 2949 1821 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13040 1821 5676 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13039 1820 1915 1919 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13038 1821 1916 1820 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13037 7955 8369 7876 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13036 7876 7957 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13035 8552 8065 7955 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13034 7875 7955 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13033 5521 6311 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13032 8552 5843 5521 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13031 5520 7049 5521 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13030 5521 5844 5520 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13029 5520 5617 5619 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13028 5619 8586 5520 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13027 7546 7274 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13026 7200 7658 7274 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13025 7198 7273 7200 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13024 7199 7881 7198 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13023 8552 7877 7199 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13022 6489 8000 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13021 6934 8065 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13020 4563 5036 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13019 1008 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13018 8552 6717 1008 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13017 2542 1008 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13016 5392 5803 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13015 8552 5812 5392 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13014 5390 5392 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13013 8552 6708 6690 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13012 8552 8065 6689 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13011 6690 6689 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13010 5840 6271 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13009 8552 5843 5840 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13008 5842 8553 5840 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13007 5840 5844 5842 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13006 5842 5839 5841 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13005 5841 7947 5842 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13004 6312 6316 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13003 4558 4747 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13002 8568 8570 8496 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13001 8552 8567 8496 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13000 8496 8569 8568 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12999 8577 8568 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12998 3925 3929 3786 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12997 3787 3930 3925 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12996 8552 3921 3787 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12995 3921 3925 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12994 3920 3930 3921 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12993 8552 4121 3930 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12992 3929 3930 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12991 8552 3927 3928 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12990 3786 3928 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12989 3785 3802 3920 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12988 8552 4747 3785 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12987 4747 3920 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12986 8552 3920 4747 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12985 4059 3650 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12984 8552 3651 4059 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12983 8552 6285 1797 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12982 1797 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12981 1797 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12980 8552 3964 1797 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12979 1870 1797 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12978 7127 3134 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12977 3134 5192 3032 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12976 8552 6021 3032 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12975 3032 3133 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12974 3031 3294 3134 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12973 3032 3295 3031 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12972 7614 8627 7850 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12971 7635 8103 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12970 8552 7635 7614 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12969 2982 2979 2981 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12968 2980 2978 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12967 8552 2980 2982 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12966 7950 7948 7872 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12965 7870 7953 7950 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12964 8552 7949 7870 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12963 7949 7950 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12962 7945 7953 7949 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12961 8552 8674 7953 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12960 7948 7953 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12959 8552 7951 7952 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12958 7872 7952 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12957 7869 7946 7945 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12956 8552 7947 7869 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12955 7947 7945 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12954 8552 7945 7947 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12953 8371 8368 8370 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12952 8552 8366 8370 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12951 8370 8369 8371 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12950 8367 8371 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12949 4517 4718 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12948 4516 4519 4517 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12947 8552 4706 4516 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12946 8063 8346 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12945 8552 8347 8063 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12944 2573 3767 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12943 2573 2764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12942 8552 3960 2573 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12941 6107 7353 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12940 8552 7592 6107 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12939 6789 6817 7691 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12938 6788 6818 6789 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12937 8552 6900 6788 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12936 4670 4676 4607 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12935 4608 4677 4670 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12934 8552 4668 4608 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12933 4668 4670 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12932 4667 4677 4668 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12931 8552 6232 4677 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12930 4676 4677 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12929 8552 4673 4675 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12928 4607 4675 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12927 4606 4605 4667 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12926 8552 6283 4606 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12925 6283 4667 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12924 8552 4667 6283 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12923 2920 3254 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12922 2920 3668 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12921 8552 3106 2920 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12920 2798 2586 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12919 2798 2764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12918 8552 3960 2798 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12917 7574 8237 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12916 7574 8098 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12915 8552 8246 7574 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12914 4344 4564 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12913 8552 4342 4344 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12912 4788 4344 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12911 3275 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12910 3275 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12909 8552 5013 3275 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12908 8552 4715 3275 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12907 3668 7718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12906 3668 3677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12905 8552 3678 3668 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12904 3472 4999 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12903 3472 3471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12902 8552 3885 3472 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12901 8455 8780 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12900 8455 8209 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12899 8552 8782 8455 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12898 7653 8132 7598 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12897 7598 7933 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12896 8552 7932 7653 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12895 7930 7653 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12894 8552 8121 7492 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12893 8552 8627 7270 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12892 7492 7270 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12891 4623 5643 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12890 4744 5644 4623 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12889 8552 4754 4744 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12888 7884 8566 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12887 8552 8135 7884 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12886 6672 6964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12885 6672 7184 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12884 8552 8490 6672 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12883 8552 8240 6672 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12882 3306 3493 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12881 8552 4792 3306 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12880 3305 3306 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12879 7650 8585 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12878 8552 8627 7650 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12877 5410 7880 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12876 5411 6007 5410 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12875 8552 5851 5411 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12874 8552 5446 5447 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12873 5853 5447 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12872 8552 5447 5853 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12871 8552 5447 5853 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12870 5853 5447 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12869 8552 5853 5852 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12868 6272 5852 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12867 8552 5852 6272 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12866 8552 5852 6272 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12865 6272 5852 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12864 8552 5853 5854 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12863 7315 5854 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12862 8552 5854 7315 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12861 8552 5854 7315 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12860 7315 5854 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12859 8552 195 194 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12858 193 194 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12857 8552 194 193 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12856 8552 194 193 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12855 193 194 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12854 8552 193 191 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12853 5563 191 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12852 8552 191 5563 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12851 8552 191 5563 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12850 5563 191 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12849 8552 193 192 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12848 5471 192 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12847 8552 192 5471 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12846 8552 192 5471 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12845 5471 192 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12844 610 2159 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12843 8552 1980 610 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12842 609 610 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12841 8552 2847 2800 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12840 2800 4230 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12839 8552 2798 2800 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12838 3058 2800 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12837 8552 6132 5706 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12836 5706 5702 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12835 8552 5703 5706 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12834 5957 5706 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12833 8552 1564 1434 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12832 1434 1566 1992 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12831 5435 6246 5437 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12830 5437 5436 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12829 8552 7534 5435 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12828 5434 5435 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12827 5255 5258 5073 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12826 5074 5259 5255 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12825 8552 5251 5074 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12824 5251 5255 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12823 5250 5259 5251 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12822 8552 6361 5259 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12821 5258 5259 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12820 8552 5496 5257 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12819 5073 5257 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12818 5072 5105 5250 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12817 8552 5498 5072 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12816 5498 5250 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12815 8552 5250 5498 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12814 8552 3898 1039 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12813 1039 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12812 1039 5013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12811 8552 3531 1039 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12810 1382 1039 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12809 6723 7115 6638 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12808 6638 7118 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12807 8552 8372 6723 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12806 6816 6723 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12805 4573 4791 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12804 8552 4565 4573 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12803 3254 2538 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12802 2539 2537 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12801 8552 2949 2540 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12800 8552 4319 2536 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12799 2536 2540 2538 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12798 2538 2949 2539 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12797 3673 2141 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12796 2142 2537 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12795 8552 2949 2143 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12794 8552 2145 2140 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12793 2140 2143 2141 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12792 2141 2949 2142 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12791 175 2976 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12790 8552 807 175 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12789 181 4346 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12788 8552 2974 181 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12787 4978 4977 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12786 4978 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12785 8552 7315 4978 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12784 1452 1716 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12783 1454 2498 1401 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12782 1401 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12781 8552 1449 1403 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12780 1403 1455 1402 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12779 1402 1452 1454 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12778 1454 1716 1404 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12777 8552 3414 1449 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12776 1447 1454 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12775 1404 1722 1403 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12774 2661 2936 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12773 8552 3078 2661 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12772 3654 2661 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12771 3661 4693 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12770 8552 3838 3661 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12769 3660 3661 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12768 1552 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12767 1552 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12766 8552 6040 1552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12765 6526 6662 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12764 8552 6661 6526 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12763 6252 5998 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12762 6252 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12761 8552 6272 6252 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12760 2659 2920 2607 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12759 2607 3665 2659 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12758 8552 3257 2607 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12757 4529 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12756 4529 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12755 8552 5471 4529 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12754 6644 6736 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12753 6646 7073 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12752 8552 8430 6737 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12751 8552 6910 6645 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12750 6645 6737 6736 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12749 6736 8430 6646 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12748 7159 6933 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12747 6756 7367 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12746 8552 6934 6935 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12745 8552 7153 6755 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12744 6755 6935 6933 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12743 6933 6934 6756 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12742 6919 6922 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12741 6752 7169 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12740 8552 6934 6923 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12739 8552 6920 6750 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12738 6750 6923 6922 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12737 6922 6934 6752 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12736 8552 3398 3250 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12735 3250 3395 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12734 8552 3411 3250 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12733 3389 3250 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12732 2564 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12731 2564 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12730 8552 5465 2564 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12729 8552 4300 2564 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12728 7394 7319 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12727 7216 7320 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12726 8552 8430 7322 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12725 8552 7323 7215 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12724 7215 7322 7319 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12723 7319 8430 7216 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12722 502 504 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12721 505 4068 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12720 8552 988 506 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12719 8552 721 503 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12718 503 506 504 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12717 504 988 505 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12716 8229 8487 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12715 8552 8227 8229 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12714 8458 8229 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12713 6321 6889 6322 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12712 6322 7735 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12711 8552 6466 6321 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12710 6320 6321 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12709 3267 5408 3268 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12708 3268 6859 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12707 8552 6265 3267 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12706 3266 3267 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12705 7923 7857 7856 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12704 8552 7855 7856 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12703 7856 8063 7923 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12702 8061 7923 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12701 4548 4550 4547 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12700 4549 4552 4548 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12699 8552 4546 4549 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12698 4546 4548 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12697 4545 4552 4546 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12696 8552 6512 4552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12695 4550 4552 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12694 8552 4554 4551 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12693 4547 4551 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12692 4544 4543 4545 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12691 8552 4758 4544 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12690 4758 4545 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12689 8552 4545 4758 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12688 8552 3898 2752 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12687 2752 3956 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12686 8552 2986 2752 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12685 2754 2752 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12684 8552 7358 7166 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12683 7166 7362 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12682 7166 7356 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12681 8552 8019 7166 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12680 7165 7166 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12679 4125 4126 4124 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12678 4124 4217 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12677 8552 4553 4125 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12676 4123 4125 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12675 8552 6718 3764 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12674 3764 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12673 3764 6717 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12672 8552 5192 3764 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12671 3763 3764 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12670 1782 2890 8552 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_12669 1781 2161 1782 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_12668 1780 1779 1781 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_12667 8552 2572 1780 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_12666 8552 6285 5195 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12665 5195 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12664 8552 5192 5195 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12663 7308 5195 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12662 7261 7268 7196 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12661 7195 7267 7261 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12660 8552 7260 7195 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12659 7260 7261 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12658 7258 7267 7260 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12657 8552 8596 7267 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12656 7268 7267 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12655 8552 7326 7265 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12654 7196 7265 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12653 7194 7193 7258 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12652 8552 7257 7194 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12651 7257 7258 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12650 8552 7258 7257 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12649 8552 1037 1038 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12648 1038 1997 2584 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12647 2190 2189 3755 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12646 2188 2187 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12645 8552 2188 2190 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12644 7133 7139 7136 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12643 7134 7138 7133 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12642 8552 7132 7134 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12641 7132 7133 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12640 7130 7138 7132 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12639 8552 8728 7138 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12638 7139 7138 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12637 8552 7135 7137 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12636 7136 7137 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12635 7131 7129 7130 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12634 8552 7140 7131 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12633 7140 7130 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12632 8552 7130 7140 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12631 3400 7142 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12630 3400 3677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12629 8552 3678 3400 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12628 4537 5643 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12627 4538 5644 4537 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12626 8552 5870 4538 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12625 1843 2890 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12624 1842 1980 1982 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12623 2769 1982 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12622 1982 2315 1843 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12621 8552 3048 1842 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12620 5205 5207 5066 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12619 5065 5208 5205 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12618 8552 5200 5065 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12617 5200 5205 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12616 5198 5208 5200 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12615 8552 6512 5208 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12614 5207 5208 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12613 8552 5459 5204 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12612 5066 5204 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12611 5064 5095 5198 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12610 8552 5872 5064 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12609 5872 5198 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12608 8552 5198 5872 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12607 8552 1798 1438 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12606 1439 1602 1999 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12605 1437 1596 1439 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12604 1438 1590 1437 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12603 1363 2764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12602 8552 4300 1363 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12601 7904 8237 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12600 7904 8236 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12599 8552 8246 7904 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12598 8232 7770 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12597 8232 7912 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12596 8552 7771 8232 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12595 8552 8019 8232 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12594 1743 2277 1694 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12593 8552 1956 1694 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12592 1694 2937 1743 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12591 1744 1743 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12590 3396 3411 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12589 3396 3398 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12588 8552 3395 3396 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12587 8552 3479 2510 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12586 2510 2942 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12585 8552 2940 2510 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12584 2509 2510 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12583 8768 7691 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12582 8552 7690 8768 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12581 6115 8240 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12580 6115 8019 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12579 8552 8490 6115 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12578 7771 8488 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12577 7771 7593 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12576 8552 7592 7771 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12575 8552 8240 7771 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12574 4322 5557 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12573 8552 4321 4322 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12572 4320 4322 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12571 7482 7480 7483 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12570 7483 7481 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12569 8552 8350 7482 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12568 7478 7482 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12567 8552 2803 2638 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12566 2805 2804 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12565 2638 2802 2804 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12564 8552 4476 4478 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12563 4477 4476 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12562 4483 6720 4477 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12561 4477 4478 4483 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12560 8552 4475 4477 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12559 4475 6720 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12558 8552 2117 2118 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12557 2116 2117 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12556 4258 2128 2116 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12555 2116 2118 4258 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12554 8552 2115 2116 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12553 2115 2128 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12552 7531 7528 7530 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12551 7530 7529 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12550 8552 8363 7531 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12549 7678 7531 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12548 3543 3765 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12547 8552 5044 3543 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12546 3541 3543 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12545 8552 3944 3319 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12544 3319 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12543 3317 3516 3319 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12542 3316 3314 3317 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12541 3319 3315 3316 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12540 8552 2976 178 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12539 178 391 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12538 8552 807 178 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12537 177 178 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12536 3856 5408 3794 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12535 3794 6720 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12534 8552 6268 3856 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12533 3854 3856 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12532 8552 6282 3292 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12531 3292 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12530 3292 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12529 8552 4522 3292 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12528 3291 3292 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12527 86 89 85 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12526 87 90 86 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12525 8552 84 87 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12524 84 86 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12523 82 90 84 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12522 8552 1302 90 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12521 89 90 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12520 8552 534 88 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12519 85 88 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12518 81 80 82 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12517 8552 532 81 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12516 532 82 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12515 8552 82 532 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12514 3082 2945 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12513 8552 2944 3082 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12512 8552 4927 4926 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12511 4925 4927 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12510 4937 6433 4925 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12509 4925 4926 4937 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12508 8552 4924 4925 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12507 4924 6433 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12506 5107 5269 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12505 5267 6115 5107 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12504 8552 5265 5267 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12503 1925 1926 1823 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12502 1823 1931 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12501 8552 1923 1925 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12500 1924 1925 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12499 2499 5406 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12498 8552 2501 2499 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12497 2192 2588 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12496 8552 2376 2192 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12495 4156 5702 4155 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12494 4155 4157 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12493 8552 4154 4156 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12492 4153 4156 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12491 6109 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12490 8552 6352 6109 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12489 6291 6290 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12488 8552 6316 6291 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12487 7973 7971 7892 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12486 7890 7976 7973 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12485 8552 7972 7890 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12484 7972 7973 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12483 7966 7976 7972 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12482 8552 8674 7976 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12481 7971 7976 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12480 8552 7974 7975 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12479 7892 7975 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12478 7889 7968 7966 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12477 8552 7969 7889 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12476 7969 7966 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12475 8552 7966 7969 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12474 5272 7347 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12473 8552 5270 5272 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12472 5914 8227 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12471 8552 6940 5914 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12470 7509 7512 7508 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12469 7510 7513 7509 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12468 8552 7507 7510 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12467 7507 7509 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12466 7506 7513 7507 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12465 8552 8674 7513 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12464 7512 7513 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12463 8552 7515 7511 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12462 7508 7511 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12461 7505 7504 7506 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12460 8552 7514 7505 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12459 7514 7506 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12458 8552 7506 7514 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12457 3974 6966 3805 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12456 3805 4157 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12455 8552 3972 3974 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12454 3973 3974 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12453 608 607 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12452 494 1019 607 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12451 493 492 494 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12450 8552 684 493 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12449 6422 6250 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12448 6422 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12447 8552 7315 6422 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12446 4533 3753 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12445 4533 6037 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12444 8552 4109 4533 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12443 328 330 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12442 224 3709 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12441 8552 988 332 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12440 8552 765 223 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12439 223 332 330 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12438 330 988 224 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12437 259 261 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12436 204 3843 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12435 8552 988 262 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12434 8552 274 203 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12433 203 262 261 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12432 261 988 204 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12431 291 293 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12430 212 3849 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12429 8552 988 295 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12428 8552 538 211 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12427 211 295 293 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12426 293 988 212 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12425 5018 5246 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12424 5020 8427 5017 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12423 5017 6307 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12422 8552 5016 5022 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12421 5022 5237 5019 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12420 5019 5018 5020 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12419 5020 5246 5021 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12418 8552 6307 5016 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12417 5015 5020 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12416 5021 5790 5022 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12415 8552 3677 3421 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12414 3421 3678 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12413 8552 7718 3421 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12412 3666 3421 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12411 3493 5192 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12410 3493 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12409 8552 5013 3493 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12408 1292 1293 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12407 1295 4068 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12406 8552 1525 1296 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12405 8552 1297 1294 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12404 1294 1296 1293 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12403 1293 1525 1295 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12402 8552 5438 4983 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12401 4983 5557 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12400 8552 4988 4983 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12399 5169 4983 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12398 8552 3467 3468 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12397 4299 3468 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12396 8552 3468 4299 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12395 8552 3468 4299 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12394 4299 3468 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12393 8552 4299 4283 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12392 7273 4283 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12391 8552 4283 7273 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12390 8552 4283 7273 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12389 7273 4283 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12388 1313 1915 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12387 1315 1309 1312 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12386 1312 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12385 8552 1311 1317 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12384 1317 1310 1314 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12383 1314 1313 1315 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12382 1315 1915 1316 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12381 8552 3414 1311 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12380 1723 1315 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12379 1316 1916 1317 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12378 2898 2788 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12377 2636 3000 2788 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12376 2637 2787 2636 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12375 8552 3007 2637 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12374 6630 6700 7320 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12373 8552 8135 6700 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12372 6631 6864 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12371 7320 8135 6631 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12370 8552 6701 6630 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12369 8552 4299 4101 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12368 7880 4101 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12367 8552 4101 7880 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12366 8552 4101 7880 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12365 7880 4101 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12364 2975 2974 2977 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12363 2977 4046 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12362 8552 4138 2975 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12361 2976 2975 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12360 6395 6413 7713 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12359 8552 8065 6413 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12358 6396 6852 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12357 7713 8065 6396 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12356 8552 6410 6395 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12355 8552 5465 4764 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12354 4764 5013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12353 4764 6026 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12352 8552 6514 4764 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12351 5669 4764 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12350 8552 4541 4542 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12349 5849 4542 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12348 8552 4542 5849 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12347 8552 4542 5849 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12346 5849 4542 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12345 8552 5849 5850 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12344 6254 5850 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12343 8552 5850 6254 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12342 8552 5850 6254 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12341 6254 5850 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12340 8552 5849 4991 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12339 6878 4991 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12338 8552 4991 6878 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12337 8552 4991 6878 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12336 6878 4991 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12335 8552 5785 3837 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12334 3793 5785 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12333 3835 3832 3793 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12332 3793 3837 3835 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12331 8552 3833 3793 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12330 3833 3832 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12329 1905 3657 1818 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12328 1818 1907 1905 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12327 1817 1914 1818 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12326 1818 2122 1817 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12325 1901 1905 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12324 8552 1902 1817 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12323 1817 2120 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12322 1707 1709 1708 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12321 1708 2511 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12320 8552 2936 1707 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12319 1706 1707 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12318 3664 3685 3663 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12317 3663 3666 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12316 8552 3673 3664 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12315 3662 3664 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12314 8552 7364 7359 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12313 7359 7358 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12312 8552 7356 7359 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12311 7357 7359 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12310 106 111 109 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12309 107 112 106 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12308 8552 105 107 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12307 105 106 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12306 103 112 105 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12305 8552 1516 112 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12304 111 112 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12303 8552 307 110 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12302 109 110 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12301 104 102 103 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12300 8552 555 104 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12299 555 103 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12298 8552 103 555 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12297 2913 4469 2912 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12296 2912 3639 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12295 8552 2910 2913 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12294 2911 2913 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12293 1704 1706 1705 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12292 1705 1886 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12291 8552 1710 1704 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12290 1882 1704 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12289 1543 1978 1433 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12288 1433 1977 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12287 8552 1641 1543 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12286 1765 1543 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12285 253 256 201 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12284 202 257 253 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12283 8552 250 202 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12282 250 253 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12281 248 257 250 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12280 8552 1302 257 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12279 256 257 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12278 8552 502 255 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12277 201 255 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12276 200 234 248 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12275 8552 721 200 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12274 721 248 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12273 8552 248 721 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12272 8552 3058 3174 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12271 3174 3061 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12270 3174 3546 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12269 8552 3973 3174 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12268 3175 3174 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12267 8552 2586 1799 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12266 1799 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12265 1799 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12264 8552 5013 1799 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12263 1798 1799 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12262 4556 4754 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12261 6889 4557 4556 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12260 8552 4558 6889 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12259 3249 3246 3248 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12258 3248 3247 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12257 8552 3646 3249 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12256 3641 3249 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12255 8552 4324 3374 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12254 3372 3485 3637 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12253 3373 3484 3372 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12252 3374 4330 3373 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12251 3030 3285 3126 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12250 3029 3291 3030 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12249 8552 3288 3029 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12248 6729 7115 6640 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12247 6640 7118 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12246 8552 7969 6729 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12245 6820 6729 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12244 8643 8645 8515 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12243 8514 8647 8643 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12242 8552 8637 8514 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12241 8637 8643 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12240 8635 8647 8637 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12239 8552 8674 8647 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12238 8645 8647 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12237 8552 8639 8642 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12236 8515 8642 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12235 8513 8512 8635 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12234 8552 8634 8513 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12233 8634 8635 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12232 8552 8635 8634 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12231 1641 2764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12230 8552 3531 1641 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12229 1553 2764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12228 8552 2586 1553 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12227 8477 8237 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12226 8477 8236 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12225 8552 8235 8477 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12224 8771 8485 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12223 8771 8486 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12222 8552 8487 8771 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12221 1489 1491 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12220 1413 3254 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12219 8552 1928 1493 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12218 8552 3673 1414 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12217 1414 1493 1491 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12216 1491 1928 1413 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12215 7525 7523 7957 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12214 7524 7522 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12213 8552 7524 7525 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12212 8552 8362 8360 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12211 8360 8625 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12210 8552 8623 8360 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12209 8630 8360 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12208 3281 3280 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12207 8552 4285 3281 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12206 4832 4835 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12205 4645 6548 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12204 8552 8764 4837 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12203 8552 4833 4644 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12202 4644 4837 4835 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12201 4835 8764 4645 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12200 2887 2727 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12199 2887 2550 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12198 8552 2732 2887 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12197 8552 3885 2887 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12196 8552 3763 3380 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12195 3771 3530 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12194 3380 3529 3530 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12193 1066 1114 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12192 1119 1113 1066 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12191 8552 7877 1119 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12190 8034 8116 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12189 8335 8343 8034 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12188 8552 8117 8335 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12187 8552 4532 2310 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12186 2310 3716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12185 2310 2315 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12184 8552 3717 2310 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12183 2307 2310 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12182 8552 1772 1773 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12181 1773 2160 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12180 1773 2559 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12179 8552 2161 1773 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12178 1771 1773 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12177 8552 7749 6667 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12176 6666 6768 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12175 6667 6665 6768 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12174 8552 8027 7634 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12173 7634 8479 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12172 7767 8490 7634 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12171 7633 8242 7767 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12170 7634 8026 7633 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12169 8552 2986 164 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12168 1015 165 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12167 164 163 165 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12166 7061 7063 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12165 7060 7243 7061 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12164 8552 7059 7060 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12163 3883 4105 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12162 8552 4108 3883 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12161 3881 3883 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12160 3299 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12159 8552 5013 3299 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12158 3745 3299 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12157 6356 6362 6359 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12156 6357 6363 6356 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12155 8552 6355 6357 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12154 6355 6356 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12153 6353 6363 6355 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12152 8552 6361 6363 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12151 6362 6363 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12150 8552 6358 6360 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12149 6359 6360 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12148 6354 6351 6353 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12147 8552 6352 6354 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12146 6352 6353 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12145 8552 6353 6352 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12144 8552 6717 3941 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12143 3941 5562 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12142 8552 6716 3941 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12141 3942 3941 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12140 3083 2949 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12139 8552 6925 3083 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12138 6795 7175 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12137 6955 7169 6795 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12136 8552 8480 6955 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12135 5228 5229 5069 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12134 5068 5232 5228 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12133 8552 5223 5068 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12132 5223 5228 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12131 5221 5232 5223 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12130 8552 6512 5232 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12129 5229 5232 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12128 8552 6659 5230 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12127 5069 5230 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12126 5067 5100 5221 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12125 8552 5220 5067 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12124 5220 5221 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12123 8552 5221 5220 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12122 6894 7126 6786 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12121 6786 7127 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12120 8552 8168 6894 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12119 6893 6894 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12118 7732 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12117 8552 8000 7732 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12116 2139 8427 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12115 2139 3677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12114 8552 3678 2139 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12113 2918 2920 2883 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12112 8552 3257 2883 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12111 2883 3665 2918 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12110 3065 2918 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12109 8552 4139 3804 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12108 3804 3944 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12107 3969 3960 3804 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12106 3803 7115 3969 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12105 3804 3942 3803 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12104 6377 8478 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12103 8552 8240 6377 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12102 313 315 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12101 219 3680 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12100 8552 983 316 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12099 8552 554 218 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12098 218 316 315 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12097 315 983 219 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12096 5911 8227 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12095 8552 7353 5911 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12094 2519 2517 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12093 8552 2707 2519 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12092 2518 2519 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12091 2502 5406 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12090 8552 2501 2502 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12089 2500 2502 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12088 4795 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12087 4795 5013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12086 8552 5562 4795 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12085 8552 7905 4795 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12084 5844 3716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12083 8552 3717 5844 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12082 5059 8478 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12081 5059 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12080 8552 5280 5059 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12079 8552 6378 5059 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12078 3547 6717 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12077 3547 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12076 8552 4109 3547 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12075 8552 3531 3547 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12074 920 922 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12073 923 3843 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12072 8552 1525 924 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12071 8552 1092 921 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12070 921 924 922 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12069 922 1525 923 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12068 7575 7741 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12067 8552 7573 7575 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12066 8446 8213 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12065 8213 8217 8043 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12064 8552 8235 8043 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12063 8043 8215 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12062 8042 8226 8213 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12061 8043 8220 8042 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12060 6394 6433 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12059 7485 6860 6394 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12058 8552 6408 7485 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12057 2486 2498 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12056 2488 2499 2485 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12055 2485 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12054 8552 2484 2490 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12053 2490 2666 2487 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12052 2487 2486 2488 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12051 2488 2498 2489 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12050 8552 3414 2484 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12049 2662 2488 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12048 2489 2678 2490 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12047 728 730 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12046 650 4068 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12045 8552 779 731 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12044 8552 726 649 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12043 649 731 730 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12042 730 779 650 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12041 1521 1524 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12040 1421 3709 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12039 8552 1525 1527 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12038 8552 1522 1420 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12037 1420 1527 1524 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12036 1524 1525 1421 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12035 8552 8349 8340 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12034 8340 8346 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12033 8552 8347 8340 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12032 8343 8340 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12031 8552 6447 6449 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12030 6449 6446 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12029 8552 6637 6449 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12028 7288 6449 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12027 6770 7394 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12026 6770 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12025 8552 8222 6770 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12024 8552 8237 6770 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12023 777 782 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12022 666 2718 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12021 8552 779 780 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12020 8552 994 665 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12019 665 780 782 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12018 782 779 666 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12017 4824 7181 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12016 8552 4822 4824 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12015 4823 4824 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12014 8552 4985 4739 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12013 4739 4987 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12012 4739 4984 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12011 8552 4986 4739 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12010 7529 4739 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12009 8552 415 413 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12008 628 413 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12007 8552 413 628 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12006 8552 413 628 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12005 628 413 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12004 8552 628 629 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12003 4111 629 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12002 8552 629 4111 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12001 8552 629 4111 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12000 4111 629 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11999 8552 628 412 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11998 4536 412 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11997 8552 412 4536 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11996 8552 412 4536 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11995 4536 412 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11994 1341 1338 1340 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11993 1340 1339 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11992 8552 2260 1341 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11991 2101 1341 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11990 4593 4598 4595 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11989 4594 4597 4593 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11988 8552 4592 4594 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11987 4592 4593 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11986 4590 4597 4592 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11985 8552 6361 4597 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11984 4598 4597 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11983 8552 4832 4596 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11982 4595 4596 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11981 4591 4589 4590 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11980 8552 4833 4591 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11979 4833 4590 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11978 8552 4590 4833 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11977 8552 3960 3003 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11976 3003 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11975 3003 3767 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11974 8552 5563 3003 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11973 3170 3003 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11972 6945 8235 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11971 8552 8780 6945 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11970 7169 6945 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11969 7718 7311 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11968 8168 7713 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11967 3289 2952 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11966 2952 6021 2953 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11965 8552 3297 2953 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11964 2953 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11963 2951 3294 2952 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11962 2953 3295 2951 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11961 4128 6934 4129 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11960 4129 4127 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11959 8552 8430 4128 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11958 4126 4128 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11957 7723 7320 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11956 8552 6717 828 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11955 828 3898 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11954 828 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11953 8552 4139 828 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11952 1373 828 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11951 8552 4483 4484 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11950 4482 4483 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11949 4481 4479 4482 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11948 4482 4484 4481 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11947 8552 4480 4482 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11946 4480 4479 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11945 8389 8392 8388 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11944 8386 8391 8389 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11943 8552 8387 8386 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11942 8387 8389 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11941 8385 8391 8387 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11940 8552 8674 8391 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11939 8392 8391 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11938 8552 8412 8390 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11937 8388 8390 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11936 8384 8382 8385 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11935 8552 8383 8384 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11934 8383 8385 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11933 8552 8385 8383 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11932 3446 5408 3361 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11931 3361 4502 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11930 8552 4096 3446 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11929 3445 3446 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11928 8405 8408 8406 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11927 8401 8409 8405 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11926 8552 8403 8401 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11925 8403 8405 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11924 8402 8409 8403 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11923 8552 8728 8409 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11922 8408 8409 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11921 8552 8404 8407 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11920 8406 8407 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11919 8400 8398 8402 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11918 8552 8399 8400 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11917 8399 8402 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11916 8552 8402 8399 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11915 2281 4968 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11914 8552 1119 2281 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11913 1456 1305 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11912 1306 3254 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11911 8552 1709 1307 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11910 8552 3673 1304 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11909 1304 1307 1305 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11908 1305 1709 1306 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11907 3290 3289 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11906 8552 5440 3290 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11905 3484 1967 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11904 3484 2157 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11903 8552 1966 3484 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11902 2628 2997 2771 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11901 2770 2769 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11900 8552 2770 2628 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11899 8552 4727 4723 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11898 8552 8065 4724 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11897 4723 4724 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11896 8670 8395 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11895 8396 8716 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11894 8552 8394 8397 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11893 8552 8661 8393 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11892 8393 8397 8395 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11891 8395 8394 8396 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11890 8373 8375 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11889 8376 8665 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11888 8552 8394 8377 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11887 8552 8372 8374 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11886 8374 8377 8375 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11885 8375 8394 8376 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11884 7669 7084 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11883 7085 8617 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11882 8552 8394 7086 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11881 8552 7660 7083 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11880 7083 7086 7084 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11879 7084 8394 7085 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11878 6368 8030 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11877 6368 8487 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11876 8552 8227 6368 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11875 8552 8240 6368 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11874 8161 8164 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11873 7978 8768 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11872 8552 8394 8167 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11871 8552 8160 7977 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11870 7977 8167 8164 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11869 8164 8394 7978 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11868 8552 7252 7064 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11867 7064 7065 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11866 8552 7066 7064 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11865 7243 7064 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11864 1822 2101 1922 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11863 1921 3266 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11862 8552 1921 1822 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11861 8552 1553 1162 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11860 1162 4750 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11859 1162 4529 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11858 8552 1552 1162 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11857 1538 1162 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11856 4486 4487 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11855 8552 6288 4486 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11854 4485 4486 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11853 6397 6720 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11852 6846 6860 6397 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11851 8552 6417 6846 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11850 8552 8325 7920 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11849 7920 8324 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11848 7920 8323 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11847 8552 8326 7920 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11846 8347 7920 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11845 8552 2105 1878 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11844 1813 2105 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11843 2107 1879 1813 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11842 1813 1878 2107 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11841 8552 1877 1813 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11840 1877 1879 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11839 749 5214 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11838 8552 959 749 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11837 1114 749 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11836 1504 5214 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11835 8552 1505 1504 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11834 2274 1504 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11833 8552 8236 7775 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11832 7775 8222 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11831 8552 8247 7775 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11830 8486 7775 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11829 2619 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11828 2963 3767 2619 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11827 8552 3744 2963 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11826 4950 4952 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11825 8552 5142 4950 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11824 4949 4950 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11823 1809 1812 1807 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11822 1808 1811 1809 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11821 8552 1806 1808 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11820 1806 1809 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11819 1805 1811 1806 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11818 8552 2028 1811 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11817 1812 1811 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11816 8552 2192 1810 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11815 1807 1810 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11814 1804 1803 1805 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11813 8552 5470 1804 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11812 5470 1805 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11811 8552 1805 5470 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11810 8552 3178 3179 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11809 3179 4839 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11808 8552 3546 3179 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11807 3180 3179 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11806 8552 8097 7176 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11805 7176 8098 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11804 8552 8247 7176 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11803 7175 7176 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11802 8552 5127 5126 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11801 5078 5127 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11800 5124 6843 5078 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11799 5078 5126 5124 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11798 8552 5122 5078 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11797 5122 6843 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11796 8552 2711 2614 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11795 2707 2710 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11794 2614 2709 2710 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11793 8552 613 615 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11792 615 616 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11791 615 614 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11790 8552 612 615 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11789 5214 615 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11788 8552 8478 6371 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11787 6371 8240 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11786 8552 8480 6371 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11785 6370 6371 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11784 8552 6040 1191 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11783 1191 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11782 1191 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11781 8552 3333 1191 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11780 1193 1191 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11779 5261 7589 5106 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11778 5106 5912 5261 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11777 8552 5260 5106 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11776 354 358 232 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11775 233 359 354 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11774 8552 350 233 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11773 350 354 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11772 349 359 350 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11771 8552 1367 359 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11770 358 359 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11769 8552 356 357 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11768 232 357 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11767 231 241 349 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11766 8552 767 231 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11765 767 349 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11764 8552 349 767 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11763 8552 5562 626 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11762 626 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11761 626 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11760 8552 4139 626 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11759 625 626 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11758 8552 6339 5893 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11757 8552 8717 5894 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11756 5893 5894 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11755 5683 7404 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11754 8552 7353 5683 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11753 5908 7347 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11752 8552 5907 5908 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11751 3455 3458 3365 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11750 3364 3459 3455 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11749 8552 3450 3364 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11748 3450 3455 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11747 3448 3459 3450 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11746 8552 3705 3459 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11745 3458 3459 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11744 8552 3452 3457 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11743 3365 3457 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11742 3363 3362 3448 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11741 8552 4522 3363 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11740 4522 3448 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11739 8552 3448 4522 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11738 3066 5150 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11737 8552 2481 3066 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11736 1379 1586 1795 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11735 1378 1777 1379 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11734 8552 1995 1378 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11733 4237 6670 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11732 8552 5280 4237 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11731 8444 8451 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11730 8552 8443 8444 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11729 1159 1009 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11728 1159 3490 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11727 8552 5562 1159 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11726 1494 1498 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11725 8552 1496 1494 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11724 1937 1494 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11723 3142 3141 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11722 8552 5790 3142 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11721 3485 3142 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11720 3535 5044 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11719 8552 4143 3535 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11718 3761 6717 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11717 3761 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11716 8552 6286 3761 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11715 8552 6026 3761 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11714 3762 6026 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11713 3762 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11712 8552 5013 3762 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11711 8552 4139 3762 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11710 4986 5192 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11709 4986 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11708 8552 6718 4986 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11707 3709 3711 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11706 3712 4526 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11705 8552 4075 3713 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11704 8552 8412 3710 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11703 3710 3713 3711 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11702 3711 4075 3712 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11701 2284 2286 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11700 2203 8427 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11699 8552 4530 2288 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11698 8552 5440 2202 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11697 2202 2288 2286 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11696 2286 4530 2203 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11695 356 346 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11694 230 3709 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11693 8552 779 347 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11692 8552 767 229 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11691 229 347 346 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11690 346 779 230 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11689 534 536 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11688 535 3843 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11687 8552 779 537 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11686 8552 532 533 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11685 533 537 536 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11684 536 779 535 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11683 7362 7734 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11682 8552 7578 7362 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11681 8552 5465 3893 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11680 3893 3956 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11679 3893 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11678 8552 5466 3893 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11677 4064 3893 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11676 4073 4076 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11675 4078 4935 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11674 8552 4075 4077 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11673 8552 7142 4074 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11672 4074 4077 4076 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11671 4076 4075 4078 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11670 8552 4985 4531 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11669 4531 4984 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11668 8552 4986 4531 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11667 6860 4531 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11666 1948 2139 1831 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11665 8552 1956 1831 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11664 1831 3275 1948 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11663 1946 1948 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11662 1091 5214 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11661 8552 1280 1091 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11660 2247 1091 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11659 3525 3528 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11658 3379 4152 3528 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11657 3377 3763 3379 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11656 3378 3526 3377 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11655 8552 3527 3378 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11654 3313 3314 3312 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11653 3312 3315 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11652 8552 4563 3313 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11651 3310 3313 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11650 5588 5587 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11649 8552 6843 5588 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11648 5586 5588 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11647 8552 5826 5548 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11646 8552 8065 5550 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11645 5548 5550 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11644 2223 2274 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11643 3274 2273 2223 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11642 8552 7877 3274 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11641 3293 3716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11640 8552 3717 3293 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11639 3885 3293 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11638 8552 6298 6093 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11637 5952 6298 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11636 6092 6654 5952 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11635 5952 6093 6092 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11634 8552 6090 5952 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11633 6090 6654 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11632 8552 8450 7577 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11631 7577 8209 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11630 7577 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11629 8552 8780 7577 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11628 7576 7577 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11627 5103 5245 5243 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11626 8552 7315 5245 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11625 5104 6307 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11624 5243 7315 5104 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11623 8552 6312 5103 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11622 2245 2664 2218 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11621 2218 3090 2245 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11620 8552 3257 2218 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11619 7491 7493 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11618 7493 7535 7494 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11617 8552 7492 7494 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11616 7494 7650 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11615 7490 7536 7493 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11614 7494 7533 7490 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11613 3028 7127 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11612 3121 7126 3028 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11611 8552 8427 3121 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11610 971 972 969 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11609 970 974 971 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11608 8552 968 970 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11607 968 971 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11606 967 974 968 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11605 8552 1516 974 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11604 972 974 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11603 8552 975 973 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11602 969 973 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11601 966 965 967 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11600 8552 1125 966 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11599 1125 967 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11598 8552 967 1125 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11597 2110 3652 2109 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11596 2109 2107 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11595 8552 2108 2110 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11594 4469 2110 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11593 8552 2732 2541 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11592 2541 2550 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11591 2541 2727 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11590 8552 3885 2541 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11589 3120 2541 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11588 584 587 586 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11587 583 588 584 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11586 8552 582 583 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11585 582 584 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11584 581 588 582 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11583 8552 1516 588 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11582 587 588 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11581 8552 986 585 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11580 586 585 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11579 580 579 581 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11578 8552 993 580 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11577 993 581 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11576 8552 581 993 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11575 2129 2272 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11574 8552 2133 2129 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11573 8560 8564 8495 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11572 8494 8565 8560 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11571 8552 8556 8494 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11570 8556 8560 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11569 8555 8565 8556 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11568 8552 8596 8565 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11567 8564 8565 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11566 8552 8561 8563 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11565 8495 8563 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11564 8493 8492 8555 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11563 8552 8553 8493 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11562 8553 8555 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11561 8552 8555 8553 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11560 6730 7126 6641 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11559 6641 7127 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11558 8552 8417 6730 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11557 6819 6730 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11556 8593 8597 8504 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11555 8503 8598 8593 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11554 8552 8589 8503 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11553 8589 8593 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11552 8588 8598 8589 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11551 8552 8596 8598 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11550 8597 8598 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11549 8552 8600 8595 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11548 8504 8595 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11547 8502 8501 8588 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11546 8552 8586 8502 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11545 8586 8588 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11544 8552 8588 8586 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11543 1131 1127 1068 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11542 1068 1128 1131 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11541 1067 1129 1068 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11540 1068 1124 1067 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11539 2273 1131 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11538 8552 1123 1067 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11537 1067 1125 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11536 6676 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11535 6677 8222 6676 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11534 8552 8247 6677 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11533 7629 7907 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11532 7756 8220 7629 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11531 8552 8455 7756 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11530 3735 3725 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11529 3726 3750 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11528 8552 8627 3727 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11527 8552 4305 3724 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11526 3724 3727 3725 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11525 3725 8627 3726 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11524 2514 2517 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11523 2515 2707 2514 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11522 8552 8627 2515 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11521 2716 2949 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11520 8552 5220 2716 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11519 2715 2716 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11518 3255 3254 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11517 8552 3673 3255 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11516 3257 3255 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11515 369 4111 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11514 8552 5563 369 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11513 4490 5390 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11512 8552 3846 4490 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11511 3863 3865 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11510 3784 3866 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11509 8552 8394 3868 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11508 8552 6005 3783 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11507 3783 3868 3865 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11506 3865 8394 3784 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11505 4683 4493 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11504 4492 4490 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11503 8552 8394 4494 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11502 8552 6250 4491 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11501 4491 4494 4493 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11500 4493 8394 4492 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11499 3452 3116 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11498 3027 3281 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11497 8552 8394 3118 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11496 8552 4522 3026 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11495 3026 3118 3116 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11494 3116 8394 3027 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11493 8552 6887 6886 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11492 6886 6883 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11491 8552 6882 6886 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11490 7285 6886 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11489 4027 5563 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11488 4027 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11487 8552 3753 4027 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11486 1759 1757 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11485 1954 1758 1759 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11484 8552 7877 1954 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11483 4338 5562 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11482 4338 6040 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11481 8552 4577 4338 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11480 8552 8717 4338 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11479 3693 3442 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11478 3360 3441 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11477 8552 8394 3444 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11476 8552 4501 3359 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11475 3359 3444 3442 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11474 3442 8394 3360 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11473 2527 2280 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11472 2201 2281 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11471 8552 8394 2283 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11470 8552 4977 2200 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11469 2200 2283 2280 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11468 2280 8394 2201 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11467 3777 5915 3778 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11466 3778 4157 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11465 8552 3775 3777 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11464 3776 3777 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11463 8552 1592 1436 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11462 1586 1585 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11461 1436 1584 1585 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11460 6373 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11459 6373 6940 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11458 8552 7184 6373 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11457 8552 8490 6373 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11456 2176 3956 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11455 2176 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11454 8552 6286 2176 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11453 8552 3964 2176 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11452 1851 2890 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11451 1850 2572 1990 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11450 2578 1990 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11449 1990 2161 1851 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11448 8552 3048 1850 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11447 6401 6859 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11446 7111 6873 6401 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11445 8552 6721 7111 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11444 2320 2318 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11443 2320 2743 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11442 8552 2321 2320 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11441 8552 2963 2320 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11440 1975 1769 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11439 1975 1535 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11438 8552 1766 1975 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11437 8552 1768 1975 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11436 5444 5643 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11435 5445 5644 5444 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11434 8552 6466 5445 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11433 7632 7908 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11432 8022 7906 7632 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11431 8552 7761 8022 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11430 6624 6841 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11429 6688 7246 6624 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11428 8552 6690 6688 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11427 5389 5990 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11426 8552 5805 5389 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11425 5388 5389 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11424 4955 4960 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11423 4958 4957 4960 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11422 4959 7880 4958 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11421 4956 7881 4959 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11420 8552 7877 4956 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11419 8552 8097 8021 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11418 8021 8235 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11417 8552 8215 8021 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11416 8487 8021 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11415 6264 6276 6263 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11414 6263 7713 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11413 8552 6879 6264 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11412 6262 6264 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11411 1767 1772 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11410 8552 2760 1767 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11409 1766 1767 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11408 8552 3657 1703 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11407 1703 1890 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11406 1702 1706 1703 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11405 1701 3655 1702 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11404 1703 1710 1701 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11403 8552 805 380 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11402 380 2974 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11401 8552 4350 380 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11400 378 380 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11399 4962 6246 4964 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11398 4964 4963 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11397 8552 7491 4962 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11396 4961 4962 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11395 5053 5057 5055 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11394 5054 5058 5053 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11393 8552 5052 5054 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11392 5052 5053 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11391 5050 5058 5052 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11390 8552 6361 5058 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11389 5057 5058 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11388 8552 5274 5056 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11387 5055 5056 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11386 5051 5049 5050 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11385 8552 5270 5051 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11384 5270 5050 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11383 8552 5050 5270 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11382 7208 7307 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11381 7294 7308 7208 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11380 8552 8168 7294 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11379 4066 4247 4067 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11378 4067 5112 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11377 8552 4064 4066 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11376 4065 4066 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11375 8552 3898 1594 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11374 1594 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11373 1594 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11372 8552 4577 1594 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11371 1596 1594 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11370 4150 4157 4149 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11369 4149 6373 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11368 8552 4147 4150 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11367 4148 4150 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11366 4210 4255 4169 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11365 4168 4256 4210 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11364 8552 4208 4168 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11363 4208 4210 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11362 4250 4256 4208 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11361 8552 6232 4256 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11360 4255 4256 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11359 8552 4471 4254 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11358 4169 4254 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11357 4167 4166 4250 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11356 8552 4943 4167 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11355 4943 4250 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11354 8552 4250 4943 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11353 6082 6088 5951 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11352 5950 6089 6082 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11351 8552 6081 5950 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11350 6081 6082 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11349 6080 6089 6081 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11348 8552 6512 6089 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11347 6088 6089 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11346 8552 6323 6087 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11345 5951 6087 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11344 5949 5948 6080 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11343 8552 6324 5949 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11342 6324 6080 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11341 8552 6080 6324 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11340 5185 5408 5093 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11339 5093 6279 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11338 8552 6275 5185 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11337 5183 5185 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11336 3720 3897 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11335 3721 7115 3720 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11334 8552 6027 3721 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11333 786 1147 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11332 786 1013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11331 8552 3678 786 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11330 1149 1147 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11329 1149 1151 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11328 8552 3678 1149 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11327 8475 8022 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11326 8552 8023 8475 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11325 8459 8457 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11324 8552 8458 8459 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11323 8770 8477 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11322 8552 8478 8770 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11321 1299 1456 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11320 8552 1496 1299 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11319 1712 1299 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11318 2483 2922 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11317 8552 2936 2483 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11316 2482 2483 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11315 4106 5643 4108 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11314 4107 6878 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11313 8552 4107 4106 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11312 3055 3175 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11311 8552 3772 3055 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11310 6299 5873 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11309 5874 5872 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11308 8552 6920 5875 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11307 8552 5870 5871 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11306 5871 5875 5873 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11305 5873 6920 5874 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11304 7181 7589 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11303 7181 7182 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11302 8552 7595 7181 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11301 8443 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11300 8552 8433 8443 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11299 6455 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11298 6455 6037 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11297 8552 6718 6455 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11296 8552 6311 6455 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11295 2732 2566 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11294 2732 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11293 8552 3753 2732 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11292 2574 2572 2575 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11291 2575 2890 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11290 8552 2573 2574 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11289 2576 2574 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11288 3765 3946 3766 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11287 3766 4140 3765 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11286 8552 3950 3766 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11285 2114 2247 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11284 4079 2248 2114 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11283 8552 7877 4079 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11282 6432 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11281 6432 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11280 8552 6717 6432 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11279 8552 7660 6432 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11278 517 519 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11277 520 4068 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11276 8552 983 521 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11275 8552 720 518 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11274 518 521 519 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11273 519 983 520 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11272 2239 2499 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11271 2242 2235 2193 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11270 2193 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11269 8552 2237 2195 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11268 2195 2245 2194 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11267 2194 2239 2242 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11266 2242 2499 2196 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11265 8552 3414 2237 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11264 2639 2242 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11263 2196 3090 2195 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11262 6713 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11261 6713 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11260 8552 6286 6713 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11259 8552 6290 6713 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11258 543 545 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11257 546 3849 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11256 8552 983 547 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11255 8552 542 544 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11254 544 547 545 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11253 545 983 546 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11252 4695 5408 4613 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11251 4613 6433 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11250 8552 4965 4695 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11249 4693 4695 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11248 5413 5619 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11247 8552 5445 5413 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11246 5412 5413 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11245 4500 4499 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11244 8552 5415 4500 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11243 4527 4500 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11242 2169 2170 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11241 8552 2570 2169 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11240 2172 2169 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11239 5804 5985 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11238 8552 5818 5804 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11237 5803 5804 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11236 8552 3753 3147 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11235 3147 5563 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11234 8552 5470 3147 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11233 3144 3147 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11232 7368 8098 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11231 8552 8247 7368 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11230 7367 7368 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11229 8552 5790 5131 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11228 5131 5466 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11227 8552 5415 5131 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11226 5127 5131 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11225 8552 8553 8314 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11224 8552 8627 8048 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11223 8314 8048 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11222 8552 3171 3042 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11221 3042 3170 3553 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11220 8427 8185 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11219 8412 8175 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11218 6659 7165 6658 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11217 6658 6947 6659 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11216 8552 6761 6658 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11215 5533 5662 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11214 5532 5864 5664 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11213 5660 5664 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11212 5664 5877 5533 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11211 8552 7115 5532 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11210 1360 1364 4292 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11209 1359 1362 1360 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11208 8552 1358 1359 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11207 4225 4355 4193 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11206 4192 4356 4225 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11205 8552 4223 4192 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11204 4223 4225 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11203 4349 4356 4223 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11202 8552 6361 4356 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11201 4355 4356 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11200 8552 5261 4354 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11199 4193 4354 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11198 4191 4190 4349 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11197 8552 4350 4191 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11196 4350 4349 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11195 8552 4349 4350 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11194 170 179 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11193 169 181 171 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11192 1123 171 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11191 171 177 170 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11190 8552 374 169 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11189 7323 7987 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11188 7558 7561 7557 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11187 7559 7563 7558 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11186 8552 7556 7559 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11185 7556 7558 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11184 7555 7563 7556 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11183 8552 8728 7563 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11182 7561 7563 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11181 8552 7560 7562 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11180 7557 7562 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11179 7554 7552 7555 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11178 8552 7553 7554 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11177 7553 7555 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11176 8552 7555 7553 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11175 3441 4088 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11174 8552 3274 3441 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11173 4310 4532 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11172 8552 4533 4310 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11171 6276 4310 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11170 2949 3300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11169 2949 4027 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11168 8552 4533 2949 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11167 4313 5644 4186 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11166 4186 4318 4313 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11165 8552 5643 4186 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11164 6128 6378 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11163 6128 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11162 8552 8478 6128 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11161 2168 2890 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11160 2166 6878 2167 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11159 2178 2167 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11158 2167 3716 2168 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11157 8552 3048 2166 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11156 244 1567 396 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11155 395 2986 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11154 8552 395 244 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11153 3931 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11152 3931 4132 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11151 8552 6037 3931 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11150 8552 6284 3931 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11149 618 2986 815 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11148 617 1567 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11147 8552 617 618 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11146 5035 5038 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11145 5039 7382 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11144 8552 8764 5040 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11143 8552 5036 5037 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11142 5037 5040 5038 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11141 5038 8764 5039 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11140 3150 3493 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11139 3150 3716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11138 8552 3494 3150 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11137 8552 4532 3150 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11136 8552 2727 2729 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11135 2729 2732 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11134 2729 3885 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11133 8552 2760 2729 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11132 5408 2729 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11131 3886 3885 3800 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11130 3800 4040 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11129 8552 4313 3886 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11128 3884 3886 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11127 8020 7720 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11126 7611 7718 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11125 8552 8430 7721 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11124 8552 7716 7610 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11123 7610 7721 7720 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11122 7720 8430 7611 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11121 3746 3744 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11120 3742 3753 3743 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11119 7307 3743 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11118 3743 3745 3746 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11117 8552 5192 3742 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11116 8552 1738 1735 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11115 1736 1738 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11114 2117 1923 1736 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11113 1736 1735 2117 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11112 8552 1734 1736 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11111 1734 1923 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11110 3674 3672 3675 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11109 3675 3676 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11108 8552 3673 3674 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11107 3671 3674 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11106 3548 5059 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11105 8552 3547 3548 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11104 3546 3548 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11103 8552 4473 4474 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11102 4474 4929 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11101 8552 5415 4474 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11100 4476 4474 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11099 5141 5139 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11098 8552 5415 5141 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11097 5137 5141 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11096 2364 2370 2215 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11095 2214 2371 2364 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11094 8552 2363 2214 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11093 2363 2364 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11092 2362 2371 2363 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11091 8552 3329 2371 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11090 2370 2371 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11089 8552 2805 2368 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11088 2215 2368 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11087 2213 2212 2362 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11086 8552 2566 2213 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11085 2566 2362 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11084 8552 2362 2566 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11083 8552 3898 3900 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11082 3900 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11081 8552 4577 3900 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11080 3897 3900 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11079 2623 2749 2968 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11078 2622 2958 2623 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11077 8552 2748 2622 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11076 8352 8350 8618 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11075 8351 8605 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11074 8552 8351 8352 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11073 2524 2530 2528 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11072 2525 2531 2524 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11071 8552 2523 2525 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11070 2523 2524 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11069 2521 2531 2523 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11068 8552 3705 2531 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11067 2530 2531 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11066 8552 2527 2529 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11065 2528 2529 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11064 2522 2520 2521 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11063 8552 4977 2522 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11062 4977 2521 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11061 8552 2521 4977 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11060 1574 1576 1424 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11059 1423 1578 1574 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11058 8552 1570 1423 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11057 1570 1574 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11056 1568 1578 1570 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11055 8552 2028 1578 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11054 1576 1578 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11053 8552 3005 1577 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11052 1424 1577 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11051 1422 1435 1568 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11050 8552 1567 1422 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11049 1567 1568 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11048 8552 1568 1567 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11047 8552 2320 1839 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11046 1840 2325 1973 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11045 1838 2555 1840 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11044 1839 1976 1838 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11043 3980 5703 3807 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11042 3807 4157 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11041 8552 3978 3980 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11040 3979 3980 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11039 802 1980 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11038 802 800 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11037 8552 1552 802 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11036 4682 4688 4612 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11035 4611 4689 4682 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11034 8552 4680 4611 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11033 4680 4682 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11032 4679 4689 4680 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11031 8552 6232 4689 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11030 4688 4689 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11029 8552 4683 4687 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11028 4612 4687 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11027 4610 4609 4679 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11026 8552 6250 4610 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11025 6250 4679 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11024 8552 4679 6250 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11023 5082 5851 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11022 8552 5843 5082 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11021 5083 6708 5082 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11020 5082 5844 5083 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11019 5083 5158 5160 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11018 5160 8329 5083 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11017 2534 2535 2940 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11016 2533 2532 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11015 8552 2533 2534 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11014 3509 3512 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11013 8552 6092 3509 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11012 1980 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11011 1980 3753 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11010 8552 5465 1980 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11009 7534 7538 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11008 7538 7535 7539 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11007 8552 7887 7539 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11006 7539 7884 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11005 7537 7536 7538 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11004 7539 7533 7537 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11003 988 2734 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11002 8552 1123 988 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11001 2475 2499 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11000 2478 3066 2474 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10999 2474 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10998 8552 2473 2480 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10997 2480 2476 2477 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10996 2477 2475 2478 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10995 2478 2499 2479 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10994 8552 3414 2473 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10993 2645 2478 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10992 2479 2923 2480 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10991 8134 8132 8037 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10990 8037 8359 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10989 8552 8131 8134 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10988 8356 8134 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10987 3285 2334 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10986 3285 2305 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10985 8552 4530 3285 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10984 6032 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10983 6032 6037 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10982 8552 6043 6032 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10981 8552 5851 6032 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10980 8552 1702 1698 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10979 1700 1702 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10978 2103 1710 1700 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10977 1700 1698 2103 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10976 8552 1699 1700 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10975 1699 1710 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10974 4826 8478 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10973 4826 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10972 8552 5280 4826 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10971 8552 8480 4826 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10970 3972 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10969 3972 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10968 8552 6040 3972 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10967 8552 5562 3972 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10966 3849 3851 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10965 3782 4947 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10964 8552 4075 3853 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10963 8552 8168 3781 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10962 3781 3853 3851 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10961 3851 4075 3782 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10960 5025 5043 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10959 5030 8202 5024 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10958 5024 6307 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10957 8552 5026 5028 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10956 5028 5270 5027 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10955 5027 5025 5030 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10954 5030 5043 5029 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10953 8552 6307 5026 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10952 5023 5030 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10951 5029 6288 5028 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10950 3843 3844 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10949 3780 4481 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10948 8552 4075 3847 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10947 8552 7326 3779 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10946 3779 3847 3844 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10945 3844 4075 3780 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10944 2718 2720 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10943 2604 7723 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10942 8552 4530 2722 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10941 8552 6027 2605 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10940 2605 2722 2720 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10939 2720 4530 2604 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10938 8552 3648 3649 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10937 3647 3648 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10936 3822 3646 3647 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10935 3647 3649 3822 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10934 8552 3645 3647 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10933 3645 3646 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10932 7105 7307 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10931 7106 7308 7105 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10930 8552 7142 7106 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10929 2897 2774 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10928 2629 2772 2774 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10927 2630 2773 2629 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10926 8552 3163 2630 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10925 3009 3008 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10924 2901 3544 3008 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10923 2899 3538 2901 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10922 2900 2898 2899 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10921 8552 3525 2900 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10920 7074 7075 7073 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10919 8552 8135 7075 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10918 7072 7257 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10917 7073 8135 7072 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10916 8552 7071 7074 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10915 5173 5175 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10914 5091 5174 5175 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10913 5092 7880 5091 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10912 5090 7881 5092 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10911 8552 7877 5090 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10910 4969 5153 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10909 8552 5161 4969 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10908 4968 4969 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10907 1183 2986 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10906 8552 1567 1183 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10905 2586 1183 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10904 7474 8350 7476 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10903 7473 7472 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10902 8552 7473 7474 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10901 5152 5408 5081 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10900 5081 6843 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10899 8552 6259 5152 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10898 5150 5152 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10897 4560 4557 4559 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10896 4559 4754 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10895 8552 4558 4560 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10894 8010 4560 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10893 2959 2960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10892 8552 4999 2959 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10891 2962 2959 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10890 8552 3723 3129 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10889 3129 3290 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10888 8552 3126 3129 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10887 3125 3129 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10886 8552 8450 7581 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10885 7581 8781 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10884 7581 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10883 8552 8215 7581 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10882 7582 7581 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10881 8410 8677 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10880 6910 7553 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10879 8552 3960 2581 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10878 2581 2784 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10877 8552 3767 2581 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10876 2781 2581 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10875 1080 1084 1051 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10874 1050 1085 1080 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10873 8552 1077 1050 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10872 1077 1080 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10871 1076 1085 1077 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10870 8552 1302 1085 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10869 1084 1085 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10868 8552 1292 1083 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10867 1051 1083 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10866 1049 1048 1076 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10865 8552 1297 1049 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10864 1297 1076 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10863 8552 1076 1297 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10862 4060 4059 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10861 4061 4062 4060 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10860 8552 8627 4061 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10859 5048 5284 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10858 4046 4583 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10857 8472 8461 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10856 1910 1738 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10855 8552 1737 1910 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10854 3259 3258 3260 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10853 8552 3257 3260 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10852 3260 3670 3259 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10851 3415 3259 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10850 6799 6801 6680 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10849 6679 6838 6799 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10848 8552 6798 6679 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10847 6798 6799 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10846 6833 6838 6798 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10845 8552 8596 6838 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10844 6801 6838 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10843 8552 7475 6836 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10842 6680 6836 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10841 6678 6773 6833 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10840 8552 7472 6678 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10839 7472 6833 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10838 8552 6833 7472 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10837 1479 1489 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10836 8552 1496 1479 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10835 4931 5586 4932 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10834 4932 5130 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10833 8552 5119 4931 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10832 4934 4931 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10831 1364 1363 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10830 8552 4792 1364 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10829 1362 1159 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10828 8552 1768 1362 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10827 8060 8062 7924 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10826 7925 8113 8060 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10825 8552 8058 7925 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10824 8058 8060 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10823 8109 8113 8058 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10822 8552 8596 8113 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10821 8062 8113 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10820 8552 8061 8115 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10819 7924 8115 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10818 7922 8033 8109 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10817 8552 8110 7922 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10816 8110 8109 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10815 8552 8109 8110 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10814 7620 8065 7675 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10813 7674 7947 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10812 8552 7674 7620 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10811 2884 1765 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10810 8552 1766 2884 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10809 606 1016 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10808 794 7536 606 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10807 8552 6077 794 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10806 2922 3082 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10805 2922 3092 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10804 8552 3102 2922 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10803 8552 3083 2922 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10802 6132 6378 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10801 6132 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10800 8552 7185 6132 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10799 8097 7312 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10798 7214 7311 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10797 8552 8430 7314 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10796 8552 7547 7213 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10795 7213 7314 7312 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10794 7312 8430 7214 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10793 8217 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10792 8217 8781 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10791 8552 8450 8217 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10790 8552 8215 8217 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10789 8552 6715 6712 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10788 6712 6713 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10787 8552 6714 6712 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10786 7283 6712 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10785 4147 4577 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10784 4147 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10783 8552 6029 4147 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10782 8552 5013 4147 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10781 8236 7712 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10780 7609 7713 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10779 8552 8430 7715 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10778 8552 7895 7608 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10777 7608 7715 7712 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10776 7712 8430 7609 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10775 3358 6859 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10774 3433 5408 3358 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10773 8552 6265 3433 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10772 2174 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10771 2174 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10770 8552 3490 2174 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10769 8552 5465 2174 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10768 4770 5011 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10767 8552 8433 4770 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10766 4768 4770 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10765 7186 8487 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10764 8552 7404 7186 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10763 7588 7186 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10762 6550 6553 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10761 8552 6672 6550 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10760 6549 6550 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10759 8552 2305 1764 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10758 1764 4530 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10757 8552 2334 1764 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10756 1763 1764 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10755 2984 3160 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10754 8552 4139 2984 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10753 2983 2984 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10752 8552 6644 6535 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10751 6535 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10750 6535 8246 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10749 8552 8237 6535 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10748 6537 6535 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10747 8552 2764 1589 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10746 1589 2586 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10745 8552 4139 1589 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10744 1590 1589 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10743 8552 5471 5012 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10742 5012 5465 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10741 5012 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10740 8552 6312 5012 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10739 5011 5012 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10738 8003 8001 7903 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10737 7901 8007 8003 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10736 8552 8002 7901 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10735 8002 8003 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10734 7998 8007 8002 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10733 8552 8728 8007 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10732 8001 8007 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10731 8552 8004 8005 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10730 7903 8005 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10729 7900 7999 7998 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10728 8552 8000 7900 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10727 8000 7998 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10726 8552 7998 8000 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10725 1727 1862 1728 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10724 1728 2511 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10723 8552 2936 1727 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10722 1902 1727 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10721 8552 4795 4189 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10720 4334 4333 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10719 4189 4219 4333 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10718 770 767 662 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10717 662 1128 770 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10716 661 1129 662 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10715 662 764 661 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10714 1758 770 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10713 8552 1123 661 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10712 661 765 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10711 8552 5440 5442 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10710 5443 5851 5638 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10709 5441 6311 5443 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10708 5442 6283 5441 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10707 1835 1973 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10706 2301 1972 1835 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10705 8552 2151 2301 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10704 5381 5378 5380 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10703 5382 5385 5381 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10702 8552 5379 5382 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10701 5379 5381 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10700 5377 5385 5379 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10699 8552 6232 5385 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10698 5378 5385 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10697 8552 5383 5384 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10696 5380 5384 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10695 5376 5375 5377 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10694 8552 6290 5376 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10693 6290 5377 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10692 8552 5377 6290 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10691 4063 4065 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10690 8552 5371 4063 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10689 4062 4063 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10688 7595 8487 7596 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10687 7596 7913 7595 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10686 8552 7594 7596 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10685 4564 4563 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10684 4564 5244 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10683 8552 7315 4564 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10682 2958 3494 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10681 8552 3300 2958 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10680 1525 2734 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10679 8552 5214 1525 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10678 3806 4157 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10677 3977 5703 3806 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10676 8552 3978 3977 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10675 8454 8780 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10674 8454 8450 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10673 8552 8483 8454 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10672 8744 8018 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10671 8744 8487 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10670 8552 8019 8744 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10669 5859 7315 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10668 5861 6062 5858 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10667 5858 5856 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10666 8552 5857 5863 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10665 5863 6294 5862 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10664 5862 5859 5861 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10663 5861 7315 5860 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10662 8552 5856 5857 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10661 6052 5861 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10660 5860 7718 5863 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10659 1535 1203 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10658 1535 6285 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10657 8552 3753 1535 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10656 2328 2961 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10655 2328 3767 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10654 8552 3956 2328 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10653 5702 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10652 5702 7592 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10651 8552 6940 5702 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10650 8552 8490 5702 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10649 5703 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10648 5703 7353 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10647 8552 7592 5703 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10646 8552 8490 5703 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10645 2746 2747 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10644 2620 3144 2747 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10643 2621 4768 2620 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10642 8552 2745 2621 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10641 1732 2508 1731 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10640 1731 3269 1732 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10639 8552 1956 1731 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10638 2787 2345 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10637 2230 2343 2345 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10636 2231 2344 2230 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10635 8552 3156 2231 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10634 6719 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10633 6719 6043 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10632 8552 6040 6719 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10631 8552 8661 6719 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10630 5896 8030 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10629 8552 6940 5896 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10628 5895 5896 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10627 8552 418 419 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10626 1046 419 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10625 8552 419 1046 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10624 8552 419 1046 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10623 1046 419 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10622 8552 1046 1043 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10621 3898 1043 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10620 8552 1043 3898 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10619 8552 1043 3898 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10618 3898 1043 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10617 8552 1046 1047 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10616 4109 1047 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10615 8552 1047 4109 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10614 8552 1047 4109 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10613 4109 1047 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10612 1093 5214 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10611 8552 1092 1093 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10610 1462 1093 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10609 394 4346 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10608 8552 2974 394 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10607 614 394 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10606 8552 8027 7402 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10605 7402 8488 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10604 8552 8240 7402 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10603 7400 7402 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10602 5882 5886 5884 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10601 5883 5887 5882 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10600 8552 5881 5883 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10599 5881 5882 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10598 5879 5887 5881 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10597 8552 6512 5887 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10596 5886 5887 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10595 8552 5889 5885 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10594 5884 5885 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10593 5880 5878 5879 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10592 8552 6072 5880 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10591 6072 5879 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10590 8552 5879 6072 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10589 2356 2354 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10588 8552 4148 2356 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10587 2359 2356 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10586 8552 5563 5682 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10585 5682 5562 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10584 5682 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10583 8552 8065 5682 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10582 8019 5682 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10581 1883 1702 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10580 8552 1447 1883 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10579 8552 6717 4110 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10578 4110 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10577 4110 4577 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10576 8552 5263 4110 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10575 5643 4110 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10574 8552 4529 2948 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10573 2948 4750 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10572 2948 6878 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10571 8552 4530 2948 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10570 3471 2948 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10569 6908 7140 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10568 7895 8399 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10567 2961 5470 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10566 8735 8742 8543 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10565 8542 8743 8735 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10564 8552 8734 8542 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10563 8734 8735 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10562 8733 8743 8734 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10561 8552 8758 8743 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10560 8742 8743 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10559 8552 8747 8740 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10558 8543 8740 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10557 8541 8540 8733 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10556 8552 8731 8541 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10555 8731 8733 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10554 8552 8733 8731 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10553 1455 1456 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10552 8552 1496 1455 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10551 8552 2173 1796 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10550 1796 1794 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10549 1796 1795 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10548 8552 1793 1796 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10547 3061 1796 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10546 8552 1390 196 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10545 196 2566 195 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10544 8552 2986 184 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10543 184 1567 185 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10542 5996 6251 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10541 5143 5998 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10540 1928 2277 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10539 8552 2937 1928 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10538 8552 3150 2557 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10537 2555 2558 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10536 2557 2556 2558 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10535 4976 6860 4975 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10534 4975 6288 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10533 8552 4974 4976 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10532 4973 4976 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10531 6458 8661 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10530 6458 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10529 8552 7315 6458 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10528 8683 8687 8526 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10527 8527 8689 8683 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10526 8552 8679 8527 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10525 8679 8683 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10524 8678 8689 8679 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10523 8552 8728 8689 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10522 8687 8689 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10521 8552 8684 8686 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10520 8526 8686 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10519 8525 8524 8678 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10518 8552 8677 8525 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10517 8677 8678 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10516 8552 8678 8677 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10515 1755 5183 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10514 8552 1951 1755 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10513 3141 2544 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10512 2544 4300 2545 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10511 8552 3964 2545 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10510 2545 3295 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10509 2543 2542 2544 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10508 2545 3133 2543 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10507 4972 7880 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10506 4971 6007 4972 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10505 8552 5440 4971 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10504 5460 4994 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10503 4995 7142 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10502 8552 4997 4996 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10501 8552 6271 4993 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10500 4993 4996 4994 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10499 4994 4997 4995 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10498 1945 2139 1830 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10497 1830 3275 1945 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10496 8552 1956 1830 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10495 3078 3400 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10494 3078 3082 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10493 8552 3083 3078 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10492 8552 3429 3078 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10491 6715 7514 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10490 6715 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10489 8552 7315 6715 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10488 8220 8237 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10487 8220 8781 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10486 8552 8450 8220 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10485 2572 2784 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10484 8552 3964 2572 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10483 6303 6306 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10482 6305 7326 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10481 8552 6307 6308 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10480 8552 6309 6304 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10479 6304 6308 6306 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10478 6306 6307 6305 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10477 5165 5171 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10476 8552 5166 5165 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10475 7066 5165 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10474 8552 3677 3098 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10473 3098 3678 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10472 8552 8168 3098 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10471 3095 3098 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10470 4138 6716 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10469 4138 5465 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10468 8552 5563 4138 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10467 8552 4833 4138 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10466 8552 6691 6415 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10465 8552 8065 6416 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10464 6415 6416 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10463 8344 8343 8345 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10462 8345 8348 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10461 8552 8350 8344 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10460 8603 8344 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10459 3102 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10458 3102 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10457 8552 5013 3102 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10456 8552 7472 3102 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10455 189 2566 190 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10454 188 1390 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10453 8552 188 189 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10452 8772 8771 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10451 8552 8770 8772 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10450 8769 8772 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10449 8552 5789 5792 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10448 5791 5789 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10447 5974 5790 5791 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10446 5791 5792 5974 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10445 8552 5788 5791 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10444 5788 5790 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10443 8552 3750 3751 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10442 3748 3750 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10441 3749 5790 3748 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10440 3748 3751 3749 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10439 8552 3747 3748 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10438 3747 5790 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10437 4090 4091 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10436 4036 4289 4091 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10435 4035 7880 4036 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10434 4034 7881 4035 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10433 8552 7877 4034 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10432 6661 6964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10431 6661 8030 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10430 8552 7367 6661 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10429 8552 8240 6661 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10428 8552 4715 4706 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10427 8552 8350 4708 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10426 4706 4708 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10425 3466 4750 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10424 8552 4529 3466 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10423 3463 3466 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10422 3906 4027 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10421 8552 4533 3906 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10420 5010 3906 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10419 4980 5179 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10418 8552 5173 4980 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10417 4979 4980 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10416 7495 7497 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10415 7497 7535 7498 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10414 8552 7655 7498 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10413 7498 7648 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10412 7496 7536 7497 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10411 7498 7533 7496 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10410 8552 4488 4266 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10409 4173 4488 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10408 4279 6288 4173 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10407 4173 4266 4279 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10406 8552 4265 4173 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10405 4265 6288 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10404 2679 2934 2612 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10403 2612 2931 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10402 8552 3673 2679 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10401 2678 2679 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10400 5846 6290 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10399 8552 5843 5846 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10398 5847 8572 5846 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10397 5846 5844 5847 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10396 5847 5845 5848 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10395 5848 8363 5847 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10394 2580 2764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10393 8552 2586 2580 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10392 3165 2580 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10391 8437 8441 8439 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10390 8438 8442 8437 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10389 8552 8436 8438 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10388 8436 8437 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10387 8434 8442 8436 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10386 8552 8728 8442 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10385 8441 8442 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10384 8552 8444 8440 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10383 8439 8440 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10382 8435 8432 8434 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10381 8552 8433 8435 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10380 8433 8434 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10379 8552 8434 8433 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10378 512 515 511 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10377 513 516 512 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10376 8552 509 513 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10375 509 512 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10374 510 516 509 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10373 8552 1302 516 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10372 515 516 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10371 8552 715 514 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10370 511 514 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10369 508 507 510 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10368 8552 925 508 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10367 925 510 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10366 8552 510 925 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10365 8552 5790 4646 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10364 8552 8350 4647 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10363 4646 4647 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10362 8624 8625 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10361 8552 8623 8624 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10360 2221 2251 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10359 3846 2252 2221 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10358 8552 7877 3846 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10357 3691 3695 3690 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10356 3692 3696 3691 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10355 8552 3689 3692 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10354 3689 3691 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10353 3688 3696 3689 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10352 8552 3705 3696 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10351 3695 3696 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10350 8552 3693 3694 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10349 3690 3694 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10348 3687 3686 3688 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10347 8552 4501 3687 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10346 4501 3688 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10345 8552 3688 4501 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10344 2682 3254 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10343 2682 2933 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10342 8552 2927 2682 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10341 7587 8246 7586 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10340 7586 8235 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10339 8552 8247 7587 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10338 7761 7587 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10337 2933 7723 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10336 2933 3677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10335 8552 3678 2933 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10334 3703 3706 3702 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10333 3701 3707 3703 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10332 8552 3700 3701 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10331 3700 3703 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10330 3698 3707 3700 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10329 8552 3705 3707 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10328 3706 3707 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10327 8552 3863 3704 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10326 3702 3704 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10325 3699 3697 3698 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10324 8552 6005 3699 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10323 6005 3698 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10322 8552 3698 6005 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10321 3407 5580 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10320 3410 3637 3350 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10319 3350 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10318 8552 3403 3352 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10317 3352 3405 3351 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10316 3351 3407 3410 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10315 3410 5580 3353 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10314 8552 3414 3403 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10313 3832 3410 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10312 3353 3670 3352 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10311 5269 7353 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10310 8552 7184 5269 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10309 2318 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10308 2318 6037 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10307 8552 4109 2318 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10306 779 2734 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10305 8552 1128 779 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10304 6950 8030 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10303 6950 7391 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10302 8552 7593 6950 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10301 6258 6257 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10300 8552 6878 6258 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10299 6858 6258 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10298 3067 3066 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10297 3070 5580 3016 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10296 3016 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10295 8552 3063 3019 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10294 3019 3065 3018 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10293 3018 3067 3070 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10292 3070 3066 3017 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10291 8552 3414 3063 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10290 3644 3070 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10289 3017 3662 3019 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10288 7168 8020 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10287 7353 8235 7168 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10286 8552 8237 7353 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10285 8320 8326 8319 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10284 8319 8323 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10283 8552 8627 8320 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10282 8570 8320 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10281 8327 8323 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10280 8327 8324 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10279 8552 8325 8327 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10278 8552 8326 8327 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10277 8552 6635 6442 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10276 6442 6438 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10275 8552 6439 6442 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10274 7099 6442 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10273 6287 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10272 6287 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10271 8552 6282 6287 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10270 8552 7969 6287 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10269 8552 815 816 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10268 1173 816 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10267 8552 816 1173 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10266 8552 816 1173 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10265 1173 816 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10264 8552 1173 1174 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10263 3767 1174 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10262 8552 1174 3767 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10261 8552 1174 3767 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10260 3767 1174 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10259 8552 1173 1023 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10258 3753 1023 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10257 8552 1023 3753 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10256 8552 1023 3753 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10255 3753 1023 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10254 8552 1173 1024 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10253 4577 1024 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10252 8552 1024 4577 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10251 8552 1024 4577 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10250 4577 1024 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10249 8552 2672 2468 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10248 2467 2672 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10247 3639 2662 2467 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10246 2467 2468 3639 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10245 8552 2466 2467 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10244 2466 2662 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10243 5094 5643 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10242 5196 5644 5094 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10241 8552 5872 5196 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10240 2211 3048 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10239 2210 2559 2341 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10238 2579 2341 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10237 2341 2760 2211 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10236 8552 2890 2210 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10235 8552 190 187 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10234 621 187 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10233 8552 187 621 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10232 8552 187 621 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10231 621 187 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10230 8552 621 400 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10229 3490 400 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10228 8552 400 3490 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10227 8552 400 3490 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10226 3490 400 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10225 8552 621 622 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10224 5013 622 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10223 8552 622 5013 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10222 8552 622 5013 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10221 5013 622 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10220 8552 621 620 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10219 3956 620 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10218 8552 620 3956 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10217 8552 620 3956 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10216 3956 620 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10215 8552 396 182 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10214 398 182 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10213 8552 182 398 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10212 8552 182 398 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10211 398 182 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10210 8552 398 183 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10209 5192 183 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10208 8552 183 5192 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10207 8552 183 5192 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10206 5192 183 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10205 8552 398 397 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10204 3964 397 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10203 8552 397 3964 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10202 8552 397 3964 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10201 3964 397 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10200 8552 398 399 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10199 3531 399 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10198 8552 399 3531 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10197 8552 399 3531 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10196 3531 399 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10195 8137 8630 8038 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10194 8038 8361 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10193 8552 8135 8137 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10192 8368 8137 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10191 4285 4284 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10190 4180 5428 4284 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10189 4181 7880 4180 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10188 4179 7881 4181 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10187 8552 7877 4179 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10186 8552 8020 7580 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10185 7580 8235 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10184 8552 8237 7580 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10183 7593 7580 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10182 6764 7171 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10181 8552 6765 6764 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10180 6946 6764 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10179 5098 5363 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10178 5218 5214 5098 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10177 8552 5215 5218 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10176 1800 2784 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10175 8552 3964 1800 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10174 2017 1800 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10173 5429 5428 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10172 8324 8132 5429 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10171 8552 5426 8324 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10170 1509 1517 1419 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10169 1418 1518 1509 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10168 8552 1508 1418 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10167 1508 1509 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10166 1506 1518 1508 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10165 8552 1516 1518 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10164 1517 1518 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10163 8552 1513 1514 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10162 1419 1514 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10161 1417 1432 1506 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10160 8552 1505 1417 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10159 1505 1506 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10158 8552 1506 1505 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10157 8552 805 377 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10156 377 2974 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10155 8552 4358 377 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10154 374 377 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10153 2957 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10152 8552 3956 2957 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10151 3137 2957 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10150 6971 8222 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10149 8552 8215 6971 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10148 6970 6971 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10147 2163 2890 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10146 2165 2315 2164 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10145 2570 2164 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10144 2164 2305 2163 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10143 8552 3048 2165 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10142 6280 6279 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10141 6818 6873 6280 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10140 8552 6462 6818 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10139 1900 1911 1816 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10138 1816 1898 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10137 8552 1901 1900 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10136 2105 1900 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10135 3667 3666 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10134 3665 3685 3667 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10133 8552 3673 3665 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10132 5612 4977 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10131 6006 6005 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10130 8552 8209 7738 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10129 7738 7735 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10128 7738 8782 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10127 8552 8780 7738 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10126 7734 7738 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10125 4794 5031 4635 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10124 4635 5023 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10123 8552 4792 4794 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10122 4791 4794 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10121 5485 6316 5484 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10120 5483 5907 5485 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10119 8552 5565 5483 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10118 1004 1005 1003 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10117 1000 1007 1004 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10116 8552 1002 1000 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10115 1002 1004 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10114 1001 1007 1002 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10113 8552 1516 1007 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10112 1005 1007 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10111 8552 1141 1006 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10110 1003 1006 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10109 999 998 1001 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10108 8552 1140 999 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10107 1140 1001 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10106 8552 1001 1140 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10105 1709 2255 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10104 8552 2127 1709 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10103 8552 6286 1040 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10102 1040 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10101 1040 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10100 8552 5563 1040 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10099 1592 1040 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10098 8128 8605 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10097 7521 8363 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10096 4963 4501 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10095 1837 2320 1972 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10094 1836 1975 1837 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10093 8552 2551 1836 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10092 1716 3854 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10091 8552 1308 1716 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10090 6227 5783 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10089 5787 5785 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10088 8552 6934 5786 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10087 8552 6223 5784 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10086 5784 5786 5783 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10085 5783 6934 5787 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10084 4822 7347 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10083 8552 4580 4822 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10082 3741 3744 8552 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_10081 4985 3745 3741 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_10080 3740 3739 4985 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_10079 8552 3753 3740 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_10078 7053 7058 7055 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10077 7054 7057 7053 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10076 8552 7052 7054 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10075 7052 7053 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10074 7050 7057 7052 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10073 8552 8596 7057 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10072 7058 7057 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10071 8552 7060 7056 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10070 7055 7056 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10069 7051 7048 7050 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10068 8552 7049 7051 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10067 7049 7050 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10066 8552 7050 7049 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10065 2120 2119 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10064 8552 2509 2120 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10063 6309 6313 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10062 6314 6311 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10061 8552 6312 6315 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10060 8552 6489 6310 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10059 6310 6315 6313 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10058 6313 6312 6314 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10057 6281 7969 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10056 6281 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10055 8552 7315 6281 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10054 5917 8480 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10053 5917 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10052 8552 8478 5917 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10051 4634 4787 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10050 4789 4788 4634 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10049 8552 5015 4789 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10048 5496 5499 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10047 5502 6526 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10046 8552 7347 5503 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10045 8552 5498 5500 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10044 5500 5503 5499 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10043 5499 7347 5502 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10042 6655 6757 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10041 6657 6760 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10040 8552 8764 6759 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10039 8552 6758 6656 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10038 6656 6759 6757 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10037 6757 8764 6657 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10036 5666 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10035 5666 6073 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10034 8552 5465 5666 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10033 8552 6021 5666 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10032 5425 5427 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10031 5833 7066 5425 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10030 8552 5548 5833 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10029 4839 6378 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10028 4839 6674 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10027 8552 5280 4839 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10026 7749 8223 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10025 7749 8235 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10024 8552 8450 7749 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10023 8552 8780 7749 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10022 6781 6872 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10021 6874 6873 6781 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10020 8552 6879 6874 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10019 5947 6078 6075 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10018 8552 6077 6078 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10017 5946 6319 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10016 6075 6077 5946 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10015 8552 6307 5947 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10014 7062 7252 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10013 7063 7246 7062 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10012 8552 8350 7063 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10011 8552 8236 8031 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10010 8031 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10009 8552 8247 8031 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10008 8029 8031 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10007 5633 6276 5524 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10006 5524 8202 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10005 8552 6287 5633 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10004 5631 5633 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10003 2929 2931 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10002 2930 2934 2929 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10001 8552 3673 2930 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10000 6485 6487 6385 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09999 6384 6490 6485 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09998 8552 6481 6384 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09997 6481 6485 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09996 6479 6490 6481 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09995 8552 6512 6490 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09994 6487 6490 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09993 8552 6648 6488 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09992 6385 6488 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09991 6383 6403 6479 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09990 8552 6739 6383 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09989 6739 6479 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09988 8552 6479 6739 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09987 8552 2179 2181 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09986 2181 2180 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09985 8552 2178 2181 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09984 3178 2181 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09983 3038 3049 3527 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09982 3037 3305 3038 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09981 8552 3307 3037 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09980 5493 5489 5491 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09979 5492 5495 5493 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09978 8552 5490 5492 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09977 5490 5493 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09976 5488 5495 5490 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09975 8552 6361 5495 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09974 5489 5495 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09973 8552 5685 5494 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09972 5491 5494 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09971 5487 5486 5488 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09970 8552 5565 5487 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09969 5565 5488 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09968 8552 5488 5565 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09967 6629 6872 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09966 7068 6860 6629 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09965 8552 6699 7068 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09964 4053 4050 4052 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09963 4054 4058 4053 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09962 8552 4051 4054 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09961 4051 4053 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09960 4049 4058 4051 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09959 8552 4057 4058 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09958 4050 4058 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09957 8552 4055 4056 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09956 4052 4056 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09955 4048 4047 4049 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09954 8552 6027 4048 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09953 6027 4049 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09952 8552 4049 6027 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09951 8552 6352 5943 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09950 6292 6071 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09949 5943 6070 6071 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09948 1334 1489 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09947 8552 1496 1334 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09946 1333 1334 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09945 3482 3483 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09944 3371 4324 3483 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09943 3369 3485 3371 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09942 3370 3484 3369 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09941 8552 4330 3370 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09940 8544 8746 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09939 8747 8744 8544 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09938 8552 8745 8747 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09937 6295 6292 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09936 6294 6293 6295 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09935 8552 6291 6294 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09934 7926 8347 7858 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09933 7858 8346 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09932 8552 8065 7926 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09931 7857 7926 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09930 8552 3092 2472 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09929 2472 3102 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09928 8552 3657 2472 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09927 2471 2472 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09926 6134 8030 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09925 8552 8240 6134 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09924 2334 5013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09923 2334 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09922 8552 4577 2334 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09921 5892 8478 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09920 5892 5891 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09919 8552 7349 5892 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09918 5877 6312 5876 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09917 5876 6307 5877 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09916 8552 7115 5876 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09915 8552 6458 6457 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09914 6457 6455 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09913 8552 6453 6457 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09912 7300 6457 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09911 2159 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09910 2159 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09909 8552 5562 2159 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09908 6462 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09907 6462 6286 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09906 8552 6282 6462 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09905 8552 8160 6462 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09904 1037 624 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09903 501 498 624 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09902 500 499 501 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09901 8552 625 500 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09900 3467 2950 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09899 2888 2887 2950 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09898 2885 7127 2888 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09897 2886 2884 2885 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09896 8552 7126 2886 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09895 4089 4703 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09894 8552 4090 4089 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09893 4088 4089 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09892 1601 1599 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09891 8552 1793 1601 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09890 2183 1601 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09889 800 611 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09888 497 2566 611 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09887 495 5470 497 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09886 496 1203 495 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09885 8552 1390 496 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09884 8552 7593 7410 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09883 7410 7592 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09882 8552 8490 7410 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09881 7594 7410 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09880 1847 2890 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09879 1846 2159 1986 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09878 2563 1986 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09877 1986 3717 1847 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09876 8552 3048 1846 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09875 8243 8488 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09874 8552 8240 8243 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09873 8479 8243 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09872 8552 8020 7352 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09871 7352 8098 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09870 8552 8780 7352 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09869 7349 7352 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09868 7915 7852 7851 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09867 8552 7850 7851 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09866 7851 8327 7915 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09865 8055 7915 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09864 5005 5007 5004 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09863 5006 5009 5005 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09862 8552 5003 5006 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09861 5003 5005 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09860 5002 5009 5003 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09859 8552 6512 5009 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09858 5007 5009 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09857 8552 5555 5008 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09856 5004 5008 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09855 5001 5000 5002 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09854 8552 5466 5001 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09853 5466 5002 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09852 8552 5002 5466 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09851 8552 4579 4581 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09850 4830 4581 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09849 8552 4581 4830 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09848 8552 4581 4830 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09847 4830 4581 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09846 8552 4830 4582 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09845 7347 4582 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09844 8552 4582 7347 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09843 8552 4582 7347 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09842 7347 4582 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09841 8552 4830 4831 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09840 8764 4831 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09839 8552 4831 8764 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09838 8552 4831 8764 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09837 8764 4831 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09836 7658 8329 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09835 5428 8103 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09834 4319 7329 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09833 7864 7933 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09832 8346 8132 7864 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09831 8552 7932 8346 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09830 8752 8759 8548 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09829 8547 8760 8752 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09828 8552 8751 8547 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09827 8751 8752 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09826 8750 8760 8751 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09825 8552 8758 8760 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09824 8759 8760 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09823 8552 8763 8756 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09822 8548 8756 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09821 8546 8545 8750 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09820 8552 8761 8546 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09819 8761 8750 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09818 8552 8750 8761 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09817 2910 2672 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09816 8552 2662 2910 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09815 4957 8553 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09814 3860 7472 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09813 1978 2986 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09812 8552 1567 1978 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09811 6877 7115 6782 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09810 6782 7118 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09809 8552 7514 6877 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09808 7092 6877 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09807 1324 3110 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09806 8552 1323 1324 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09805 1325 1324 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09804 7535 2784 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09803 8552 4577 7535 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09802 8745 8764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09801 8552 8731 8745 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09800 1862 2508 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09799 8552 3269 1862 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09798 556 560 558 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09797 558 1128 556 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09796 557 1129 558 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09795 558 554 557 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09794 1113 556 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09793 8552 1123 557 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09792 557 555 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09791 8552 8350 2890 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09790 8552 3158 1565 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09789 2890 1565 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09788 6256 6255 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09787 8552 6254 6256 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09786 6417 6256 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09785 1939 2138 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_09784 1942 1952 1825 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09783 1825 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09782 8552 1935 1827 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09781 1827 1937 1826 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09780 1826 1939 1942 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09779 1942 2138 1828 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09778 8552 3414 1935 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_09777 2268 1942 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09776 1828 1946 1827 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09775 6975 3874 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09774 8552 3872 6975 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09773 5529 5643 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09772 5645 5644 5529 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09771 8552 6060 5645 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09770 7579 8020 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09769 8552 8247 7579 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09768 7731 8490 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09767 7731 7593 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09766 8552 8019 7731 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09765 8552 8240 7731 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09764 8235 7143 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09763 7144 7142 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09762 8552 8430 7145 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09761 8552 7140 7141 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09760 7141 7145 7143 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09759 7143 8430 7144 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09758 4625 6077 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09757 4624 6878 4745 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09756 4990 4745 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09755 4745 4748 4625 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09754 8552 4758 4624 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09753 8552 4523 4297 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09752 4297 4302 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09751 8552 4295 4297 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09750 5176 4297 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09749 2535 6878 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09748 2535 4750 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09747 8552 3716 2535 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09746 8552 3717 2535 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09745 3036 3154 8552 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_09744 3156 4984 3036 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_09743 3035 3155 3156 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_09742 8552 4988 3035 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_09741 7275 7276 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09740 7203 7277 7276 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09739 7201 7880 7203 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09738 7202 7881 7201 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09737 8552 7499 7202 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09736 5034 7347 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09735 8552 5033 5034 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09734 5260 5034 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09733 1014 3531 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09732 1013 3753 1014 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09731 8552 1154 1013 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09730 174 378 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09729 172 181 173 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09728 1129 173 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09727 173 175 174 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09726 8552 374 172 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09725 5992 6245 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09724 8552 5989 5992 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09723 5990 5992 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09722 7174 7593 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09721 8552 7184 7174 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09720 7227 7174 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09719 6369 6541 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09718 8552 7315 6369 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09717 6374 6369 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09716 668 783 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09715 667 786 785 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09714 2302 785 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09713 785 1149 668 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09712 8552 793 667 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09711 6693 6695 6627 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09710 6628 6698 6693 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09709 8552 6696 6628 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09708 6696 6693 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09707 6692 6698 6696 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09706 8552 8596 6698 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09705 6695 6698 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09704 8552 7718 6697 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09703 6627 6697 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09702 6625 6694 6692 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09701 8552 6691 6625 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09700 6691 6692 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09699 8552 6692 6691 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09698 142 143 141 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09697 138 145 142 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09696 8552 139 138 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09695 139 142 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09694 137 145 139 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09693 8552 1516 145 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09692 143 145 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09691 8552 333 144 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09690 141 144 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09689 136 135 137 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09688 8552 764 136 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09687 764 137 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09686 8552 137 764 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09685 8552 3158 673 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09684 673 8350 836 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09683 8552 5790 5138 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09682 5079 5790 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09681 5139 5466 5079 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09680 5079 5138 5139 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09679 8552 5135 5079 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09678 5135 5466 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09677 7639 8572 7616 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09676 7616 7643 7639 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09675 8552 7641 7616 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09674 97 99 96 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09673 98 101 97 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09672 8552 93 98 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09671 93 97 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09670 94 101 93 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09669 8552 1302 101 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09668 99 101 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09667 8552 543 100 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09666 96 100 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09665 92 91 94 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09664 8552 542 92 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09663 542 94 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09662 8552 94 542 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09661 8552 3977 3770 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09660 3768 3771 3772 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09659 3769 3773 3768 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09658 3770 4152 3769 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09657 2503 2505 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09656 3265 2504 2503 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09655 8552 7877 3265 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09654 7114 7116 7541 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09653 7113 7111 7114 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09652 8552 7112 7113 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09651 5420 5418 5423 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09650 5421 5424 5420 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09649 8552 5419 5421 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09648 5419 5420 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09647 5416 5424 5419 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09646 8552 5835 5424 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09645 5418 5424 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09644 8552 5647 5422 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09643 5423 5422 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09642 5417 5414 5416 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09641 8552 5415 5417 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09640 5415 5416 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09639 8552 5416 5415 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09638 3398 3429 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09637 3398 3657 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09636 8552 3400 3398 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09635 4999 5562 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09634 4999 6282 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09633 8552 3767 4999 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09632 4720 6040 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09631 4720 4539 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09630 8552 4536 4720 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09629 8552 6021 4720 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09628 5383 5114 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09627 5061 5112 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09626 8552 6934 5115 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09625 8552 6290 5060 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09624 5060 5115 5114 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09623 5114 6934 5061 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09622 6760 6765 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09621 6760 7170 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09620 8552 7171 6760 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09619 5041 5042 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09618 5041 5043 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09617 8552 5048 5041 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09616 1017 1015 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09615 3314 1016 1017 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09614 8552 2151 3314 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09613 8552 3498 3495 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09612 3495 3494 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09611 8552 3493 3495 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09610 4321 3495 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09609 7885 7961 8175 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09608 8552 8135 7961 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09607 7886 8383 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09606 8175 8135 7886 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09605 8552 8566 7885 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09604 4288 4712 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09603 8552 4538 4288 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09602 4286 4288 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09601 4142 4137 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09600 4045 5036 4137 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09599 4044 5790 4045 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09598 8552 8731 4044 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09597 3024 3271 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09596 3388 3262 3024 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09595 8552 3261 3388 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09594 176 2976 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09593 8552 807 176 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09592 382 176 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09591 7859 7927 8202 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09590 8552 8135 7927 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09589 7860 7937 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09588 8202 8135 7860 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09587 8552 7928 7859 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09586 8552 8098 7387 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09585 7387 8246 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09584 8552 8237 7387 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09583 8227 7387 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09582 8552 8020 7375 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09581 7375 8236 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09580 8552 8247 7375 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09579 7373 7375 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09578 528 530 527 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09577 525 531 528 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09576 8552 526 525 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09575 526 528 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09574 524 531 526 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09573 8552 1302 531 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09572 530 531 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09571 8552 728 529 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09570 527 529 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09569 523 522 524 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09568 8552 726 523 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09567 726 524 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09566 8552 524 726 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09565 8552 2764 1041 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09564 1041 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09563 8552 4139 1041 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09562 1202 1041 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09561 1467 1902 1429 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09560 1429 1729 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09559 8552 1723 1467 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09558 1898 1467 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09557 4040 7228 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09556 5162 6708 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09555 8552 4109 3752 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09554 3752 3767 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09553 8552 3956 3752 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09552 3912 3752 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09551 8552 8329 8117 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09550 8552 8065 8067 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09549 8117 8067 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09548 8087 8088 7962 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09547 7963 8150 8087 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09546 8552 8085 7963 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09545 8085 8087 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09544 8145 8150 8085 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09543 8552 8674 8150 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09542 8088 8150 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09541 8552 8373 8152 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09540 7962 8152 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09539 7960 8040 8145 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09538 8552 8372 7960 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09537 8372 8145 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09536 8552 8145 8372 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09535 955 956 954 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09534 953 958 955 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09533 8552 952 953 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09532 952 955 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09531 951 958 952 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09530 8552 1516 958 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09529 956 958 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09528 8552 960 957 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09527 954 957 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09526 950 949 951 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09525 8552 959 950 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09524 959 951 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09523 8552 951 959 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09522 4289 4715 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09521 7905 8761 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09520 5042 5270 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09519 3759 3936 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09518 8552 3931 3759 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09517 4263 4485 4172 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09516 4172 4498 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09515 8552 4944 4263 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09514 4479 4263 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09513 8552 1798 1384 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09512 1385 1381 1793 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09511 1383 1382 1385 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09510 1384 1590 1383 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09509 1016 6718 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09508 8552 5563 1016 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09507 5831 5836 5830 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09506 5832 5837 5831 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09505 8552 5829 5832 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09504 5829 5831 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09503 5828 5837 5829 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09502 8552 5835 5837 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09501 5836 5837 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09500 8552 5833 5834 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09499 5830 5834 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09498 5827 5825 5828 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09497 8552 5826 5827 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09496 5826 5828 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09495 8552 5828 5826 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09494 8552 2566 1027 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09493 1028 5470 2764 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09492 1026 1203 1028 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09491 1027 1390 1026 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09490 8551 8781 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09489 8785 8782 8551 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09488 8552 8780 8785 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09487 5888 5469 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09486 8552 6072 5888 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09485 6660 6950 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09484 8552 6766 6660 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09483 7861 8327 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09482 8069 7930 7861 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09481 8552 7929 8069 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09480 3429 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09479 3429 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09478 8552 3956 3429 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09477 8552 8553 3429 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09476 7735 6733 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09475 6643 6735 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09474 8552 8430 6734 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09473 8552 6908 6642 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09472 6642 6734 6733 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09471 6733 8430 6643 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09470 7991 7725 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09469 7613 7723 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09468 8552 8423 7726 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09467 8552 7987 7612 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09466 7612 7726 7725 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09465 7725 8423 7613 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09464 7707 7549 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09463 7550 7718 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09462 8552 8423 7551 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09461 8552 7716 7548 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09460 7548 7551 7549 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09459 7549 8423 7550 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09458 5247 5484 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09457 8552 5246 5247 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09456 5244 5247 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09455 4523 4522 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09454 4523 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09453 8552 7315 4523 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09452 3405 3258 3256 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09451 3256 3670 3405 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09450 8552 3257 3256 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09449 3775 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09448 3775 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09447 8552 3960 3775 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09446 8552 5471 3775 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09445 8696 8418 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09444 8419 8417 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09443 8552 8423 8420 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09442 8552 8690 8416 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09441 8416 8420 8418 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09440 8418 8423 8419 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09439 8552 2153 2154 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09438 2154 2155 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09437 2154 2307 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09436 8552 2157 2154 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09435 3677 2154 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09434 7331 7333 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09433 7220 7575 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09432 8552 7347 7334 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09431 8552 7329 7219 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09430 7219 7334 7333 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09429 7333 7347 7220 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09428 8552 2305 2152 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09427 2152 6878 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09426 2152 4530 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09425 8552 4984 2152 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09424 3678 2152 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09423 8552 3822 3823 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09422 3790 3822 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09421 5112 3826 3790 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09420 3790 3823 5112 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09419 8552 3819 3790 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09418 3819 3826 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09417 1063 1463 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09416 1100 1462 1063 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09415 8552 2723 1100 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09414 1427 1462 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09413 3840 1463 1427 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09412 8552 7877 3840 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09411 5805 5809 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09410 5807 5810 5809 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09409 5808 7880 5807 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09408 5806 7881 5808 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09407 8552 7877 5806 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09406 7076 7079 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09405 7079 7535 7080 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09404 8552 7081 7080 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09403 7080 7077 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09402 7078 7536 7079 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09401 7080 7533 7078 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09400 7573 7167 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09399 7573 7362 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09398 8552 7358 7573 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09397 8552 7356 7573 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09396 8481 8776 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09395 8482 8479 8481 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09394 8552 8480 8482 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09393 6774 7065 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09392 6841 7066 6774 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09391 8552 8065 6841 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09390 1134 5214 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09389 8552 1140 1134 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09388 1339 1134 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09387 4151 5508 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09386 8552 5280 4151 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09385 4152 4151 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09384 7520 7879 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09383 8348 8132 7520 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09382 8552 7532 8348 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09381 159 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09380 8552 5563 159 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09379 602 159 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09378 8552 8098 7388 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09377 7388 8483 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09376 8552 8237 7388 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09375 7391 7388 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09374 7191 7245 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09373 7242 7480 7191 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09372 8552 7240 7242 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09371 1829 2274 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09370 2137 2273 1829 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09369 8552 2260 2137 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09368 1108 1113 1055 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09367 1055 1114 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09366 8552 2260 1108 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09365 1476 1108 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09364 8552 6134 5921 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09363 5921 5922 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09362 8552 6136 5921 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09361 5920 5921 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09360 2021 2026 1860 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09359 1859 2029 2021 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09358 8552 2022 1859 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09357 2022 2021 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09356 2020 2029 2022 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09355 8552 2028 2029 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09354 2026 2029 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09353 8552 2187 2027 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09352 1860 2027 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09351 1857 1858 2020 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09350 8552 2189 1857 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09349 2189 2020 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09348 8552 2020 2189 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09347 3643 3826 3642 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09346 3642 3641 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09345 8552 3827 3643 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09344 3814 3643 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09343 663 993 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09342 8552 1123 663 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09341 664 992 663 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09340 663 1129 664 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09339 664 775 1135 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09338 1135 994 664 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09337 279 532 237 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09336 237 1128 279 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09335 236 1129 237 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09334 237 276 236 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09333 1463 279 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09332 8552 1123 236 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09331 236 274 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09330 5903 5905 5902 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09329 5901 5906 5903 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09328 8552 5900 5901 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09327 5900 5903 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09326 5898 5906 5900 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09325 8552 6361 5906 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09324 5905 5906 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09323 8552 6106 5904 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09322 5902 5904 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09321 5899 5897 5898 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09320 8552 6316 5899 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09319 6316 5898 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09318 8552 5898 6316 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09317 8552 3960 1035 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09316 1035 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09315 1035 5013 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09314 8552 5192 1035 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09313 1034 1035 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09312 7123 7120 7693 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09311 7122 7121 7123 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09310 8552 7124 7122 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09309 6229 6230 6228 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09308 6224 6233 6229 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09307 8552 6225 6224 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09306 6225 6229 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09305 6226 6233 6225 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09304 8552 6232 6233 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09303 6230 6233 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09302 8552 6227 6231 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09301 6228 6231 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09300 6222 6221 6226 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09299 8552 6223 6222 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09298 6223 6226 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09297 8552 6226 6223 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09296 8552 3657 3659 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09295 3659 3658 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09294 5785 3654 3659 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09293 3656 3832 5785 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09292 3659 3655 3656 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09291 3655 2940 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09290 3655 3479 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09289 8552 2942 3655 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09288 2947 3885 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09287 2947 3478 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09286 8552 3471 2947 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09285 4145 6672 4146 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09284 4146 4157 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09283 8552 4144 4145 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09282 4143 4145 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09281 6899 7115 6790 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09280 6790 7118 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09279 8552 8661 6899 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09278 7120 6899 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09277 8552 8488 7591 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09276 7591 7759 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09275 7589 8479 7591 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09274 7590 7588 7589 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09273 7591 8027 7590 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09272 5782 5958 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09271 8552 5958 5780 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09270 5779 6223 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09269 8552 5779 5782 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09268 5782 5780 5781 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09267 5781 6223 5782 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09266 5789 5781 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09265 8552 5781 5789 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09264 4652 4658 4602 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09263 4601 4659 4652 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09262 8552 4651 4601 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09261 4651 4652 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09260 4650 4659 4651 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09259 8552 6232 4659 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09258 4658 4659 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09257 8552 4660 4657 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09256 4602 4657 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09255 4600 4599 4650 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09254 8552 5851 4600 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09253 5851 4650 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09252 8552 4650 5851 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09251 2776 2170 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09250 2776 2178 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09249 8552 2171 2776 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09248 8688 7541 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09247 8552 7540 8688 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09246 7757 8215 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09245 7757 8097 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09244 8552 8235 7757 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09243 4660 4664 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09242 4604 4662 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09241 8552 6934 4665 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09240 8552 5851 4603 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09239 4603 4665 4664 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09238 4664 6934 4604 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09237 4967 4966 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09236 8552 6432 4967 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09235 4965 4967 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09234 4326 4328 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09233 8552 5870 4326 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09232 4324 4326 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09231 2227 2301 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09230 8394 2302 2227 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09229 8552 8065 8394 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09228 4722 4720 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09227 8552 4978 4722 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09226 4974 4722 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09225 6775 6843 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09224 7641 6860 6775 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09223 8552 6844 7641 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09222 7637 7252 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09221 7637 7481 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09220 8552 7251 7637 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09219 8552 7246 7637 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09218 8552 5013 3101 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09217 3101 6029 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09216 3101 6021 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09215 8552 7472 3101 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09214 3100 3101 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09213 1965 7533 1834 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09212 1834 7536 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09211 8552 2334 1965 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09210 1967 1965 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09209 6632 6701 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09208 8552 8135 6632 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09207 8552 8731 3039 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09206 3160 3159 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09205 3039 3050 3159 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09204 8552 3158 1696 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09203 3048 1774 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09202 1696 1695 1774 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09201 6765 8490 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09200 6765 6954 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09199 8552 6673 6765 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09198 8244 8248 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09197 8552 8778 8244 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09196 8242 8244 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09195 8552 7252 7067 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09194 7067 7251 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09193 7067 7065 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09192 8552 7066 7067 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09191 7480 7067 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09190 8552 8325 8322 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09189 8322 8323 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09188 8552 8326 8322 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09187 8321 8322 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09186 8552 6728 6725 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09185 6725 6726 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09184 8552 6727 6725 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09183 7542 6725 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09182 7077 7071 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09181 8552 8135 7077 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09180 5279 5280 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09179 5279 6677 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09178 8552 8490 5279 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09177 8552 6378 5279 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09176 7888 7959 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09175 7882 7879 7959 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09174 7883 7880 7882 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09173 7878 7881 7883 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09172 8552 7877 7878 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09171 6948 7381 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09170 8552 6946 6948 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09169 6947 6948 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09168 5433 7307 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09167 5432 7308 5433 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09166 8552 8427 5432 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09165 2314 6878 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09164 8552 2315 2314 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09163 2727 2314 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09162 3555 3553 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09161 8552 3776 3555 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09160 3552 3555 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09159 5511 6118 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09158 8552 5920 5511 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09157 5510 5511 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09156 6962 8246 6796 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09155 6796 8222 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09154 8552 8780 6962 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09153 6961 6962 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09152 7648 7928 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09151 8552 8135 7648 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09150 5155 5611 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09149 8552 5411 5155 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09148 5153 5155 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09147 2924 3100 2925 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09146 2925 3095 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09145 8552 3673 2924 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09144 2923 2924 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09143 8552 8235 7179 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09142 7179 8097 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09141 7179 8246 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09140 8552 8780 7179 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09139 7178 7179 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09138 8552 3471 2724 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09137 2724 3885 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09136 8552 4999 2724 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09135 2723 2724 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09134 8552 2981 2590 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09133 2590 3012 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09132 2590 3335 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09131 8552 2589 2590 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09130 2588 2590 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09129 8552 6037 3524 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09128 3524 4109 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09127 8552 3753 3524 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09126 3944 3524 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09125 5478 5476 5480 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09124 5479 5482 5478 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09123 8552 5477 5479 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09122 5477 5478 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09121 5474 5482 5477 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09120 8552 6512 5482 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09119 5476 5482 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09118 8552 5677 5481 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09117 5480 5481 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09116 5475 5473 5474 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09115 8552 5676 5475 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09114 5676 5474 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09113 8552 5474 5676 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09112 8552 6543 6120 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09111 6120 6123 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09110 6120 6372 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09109 8552 5957 6120 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09108 6118 6120 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09107 8552 2359 2360 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09106 2360 2584 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09105 8552 3324 2360 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09104 2592 2360 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09103 8552 1592 1441 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09102 1441 1591 2185 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09101 6288 5851 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09100 6859 6027 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09099 4928 5790 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09098 2906 2644 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09097 8552 2645 2906 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09096 4502 5440 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09095 4929 5466 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09094 3307 2962 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09093 8552 2963 3307 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09092 2775 2756 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09091 2775 2569 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09090 8552 2570 2775 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09089 7104 7126 7103 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09088 7103 7127 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09087 8552 7718 7104 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09086 7102 7104 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09085 4997 4999 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09084 8552 6077 4997 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09083 4626 4747 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09082 4748 4755 4626 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09081 8552 5188 4748 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09080 6255 6000 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09079 6255 6889 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09078 8552 6272 6255 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09077 1101 3854 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09076 8552 1308 1101 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09075 1309 1101 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09074 5555 5890 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09073 8552 5554 5555 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09072 8552 1011 1012 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09071 1012 1009 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09070 1147 2542 1012 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09069 1010 3531 1147 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09068 1012 3753 1010 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09067 2649 3092 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09066 8552 3102 2649 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09065 2648 2649 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09064 2315 3767 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09063 2315 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09062 8552 6285 2315 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09061 5554 5469 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09060 8552 5466 5554 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09059 6253 6252 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09058 8552 6878 6253 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09057 6408 6253 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09056 1327 1755 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_09055 1332 1325 1326 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09054 1326 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09053 8552 1328 1330 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09052 1330 1333 1329 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09051 1329 1327 1332 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09050 1332 1755 1331 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09049 8552 3414 1328 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_09048 1923 1332 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09047 1331 1744 1330 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09046 3023 3095 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09045 3090 3100 3023 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09044 8552 3673 3090 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09043 8552 4795 1542 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09042 1542 1538 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09041 8552 1539 1542 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09040 1537 1542 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09039 8552 2754 2624 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09038 2966 2755 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09037 2624 2753 2755 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09036 8450 8187 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09035 7997 8185 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09034 8552 8430 8189 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09033 8552 8191 7996 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09032 7996 8189 8187 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09031 8187 8430 7997 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09030 8552 6864 6633 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09029 8552 8135 6705 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09028 6633 6705 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09027 6323 6325 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09026 6327 7164 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09025 8552 7347 6328 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09024 8552 6324 6326 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09023 6326 6328 6325 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09022 6325 7347 6327 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09021 2670 2682 2609 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09020 2609 2930 2670 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09019 8552 3257 2609 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09018 8552 3956 2935 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09017 2935 6043 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09016 2935 6284 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09015 8552 7228 2935 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09014 2934 2935 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09013 8483 8193 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09012 8008 8417 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09011 8552 8430 8197 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09010 8552 8690 8006 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09009 8006 8197 8193 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09008 8193 8430 8008 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09007 8552 6852 6420 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09006 8552 8135 6421 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09005 6420 6421 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09004 8552 8769 8476 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09003 8476 8475 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09002 8552 8482 8476 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09001 8474 8476 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09000 8552 3832 3348 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08999 3348 3828 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08998 3390 3827 3348 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08997 3347 3825 3390 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08996 3348 3826 3347 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08995 4141 4142 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08994 8552 4139 4141 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08993 4140 4141 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08992 4553 3158 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08991 5231 6758 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08990 7619 8128 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08989 8625 8132 7619 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08988 8552 8127 8625 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08987 8552 382 385 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08986 385 388 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08985 385 614 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08984 8552 612 385 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08983 1128 385 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08982 8445 8717 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08981 5365 5565 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08980 4759 4758 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08979 2585 2584 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08978 8552 3324 2585 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08977 2589 2585 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08976 2626 2890 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08975 2625 3717 2757 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08974 2756 2757 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08973 2757 4530 2626 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08972 8552 3048 2625 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08971 6779 6859 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08970 6861 6860 6779 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08969 8552 6858 6861 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08968 6814 6815 6709 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08967 6710 6869 6814 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08966 8552 6812 6710 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08965 6812 6814 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08964 6863 6869 6812 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08963 8552 8674 6869 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08962 6815 6869 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08961 8552 7723 6871 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08960 6709 6871 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08959 6707 6780 6863 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08958 8552 6864 6707 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08957 6864 6863 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08956 8552 6863 6864 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08955 8552 6029 3952 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08954 3952 5046 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08953 3952 5471 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08952 8552 4300 3952 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08951 3950 3952 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08950 8552 8731 4134 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08949 4134 5790 4135 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08948 1152 7533 1058 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08947 1058 7536 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08946 8552 2161 1152 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08945 1151 1152 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08944 71 73 70 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08943 66 74 71 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08942 8552 68 66 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08941 68 71 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08940 67 74 68 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08939 8552 1302 74 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08938 73 74 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08937 8552 75 72 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08936 70 72 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08935 65 64 67 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08934 8552 276 65 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08933 276 67 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08932 8552 67 276 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08931 8552 7680 7621 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08930 8361 7681 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08929 7621 7679 7681 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08928 6793 6820 7545 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08927 6792 6821 6793 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08926 8552 6819 6792 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08925 7636 8553 7484 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08924 7484 7643 7636 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08923 8552 7485 7484 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08922 6055 6057 5938 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08921 5937 6059 6055 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08920 8552 6050 5937 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08919 6050 6055 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08918 6048 6059 6050 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08917 8552 6512 6059 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08916 6057 6059 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08915 8552 6052 6058 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08914 5938 6058 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08913 5936 5935 6048 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08912 8552 6062 5936 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08911 6062 6048 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08910 8552 6048 6062 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08909 5455 5453 5454 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08908 5451 5456 5455 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08907 8552 5452 5451 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08906 5452 5455 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08905 5450 5456 5452 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08904 8552 6512 5456 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08903 5453 5456 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08902 8552 5651 5457 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08901 5454 5457 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08900 5449 5448 5450 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08899 8552 6060 5449 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08898 6060 5450 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08897 8552 5450 6060 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08896 2244 2664 2197 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08895 8552 3257 2197 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08894 2197 3090 2244 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08893 2476 2244 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08892 3258 3254 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08891 3258 3400 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08890 8552 3429 3258 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08889 4534 4532 4535 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08888 8552 6735 4535 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08887 4535 4533 4534 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08886 4966 4534 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08885 8716 7693 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08884 8552 7888 8716 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08883 1498 1500 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08882 1416 3254 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08881 8552 2263 1502 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08880 8552 3673 1415 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08879 1415 1502 1500 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08878 1500 2263 1416 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08877 8552 2255 1887 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08876 1887 2127 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08875 8552 3657 1887 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08874 1886 1887 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08873 7289 7288 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08872 8552 7291 7289 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08871 8127 7289 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08870 2763 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08869 2763 2764 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08868 8552 3960 2763 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08867 6428 6431 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08866 6431 7535 6399 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08865 8552 6633 6399 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08864 6399 6632 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08863 6398 7536 6431 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08862 6399 7533 6398 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08861 7906 8237 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08860 7906 8020 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08859 8552 8235 7906 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08858 5639 5638 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08857 8552 5637 5639 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08856 5662 5639 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08855 6376 8480 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08854 6376 8478 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08853 8552 8240 6376 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08852 7571 7574 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08851 7572 7731 7571 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08850 8552 7570 7572 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08849 7907 8247 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08848 7907 8236 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08847 8552 8483 7907 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08846 7631 7907 8552 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_08845 7759 7757 7631 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_08844 7630 7758 7759 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_08843 8552 7906 7630 8552 sg13_lv_pmos L=0.13U W=3.24U AS=0.7776P AD=0.7776P PS=6.97U PD=6.97U 
Mtr_08842 5438 4984 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08841 5438 4987 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08840 8552 4985 5438 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08839 8552 4986 5438 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08838 8552 2105 2106 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08837 2104 2105 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08836 5978 2103 2104 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08835 2104 2106 5978 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08834 8552 2102 2104 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08833 2102 2103 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08832 3006 3956 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08831 3006 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08830 8552 6718 3006 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08829 8552 6284 3006 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08828 7881 5010 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08827 7881 3903 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08826 8552 6873 7881 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08825 8552 4999 7881 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08824 7746 8247 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08823 7746 8020 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08822 8552 8236 7746 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08821 8552 3278 1096 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08820 1095 1096 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08819 8552 1096 1095 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08818 8552 1096 1095 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08817 1095 1096 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08816 8552 3278 1301 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08815 1300 1301 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08814 8552 1301 1300 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08813 8552 1301 1300 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08812 1300 1301 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08811 8552 3278 1303 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08810 1302 1303 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08809 8552 1303 1302 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08808 8552 1303 1302 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08807 1302 1303 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08806 4144 4577 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08805 4144 3960 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08804 8552 4109 4144 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08803 8552 3956 4144 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08802 5161 5163 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08801 5086 5162 5163 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08800 5084 7273 5086 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08799 5085 7881 5084 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08798 8552 7877 5085 8552 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08797 8552 8010 8009 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08796 8207 8009 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08795 8552 8009 8207 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08794 8552 8009 8207 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08793 8207 8009 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08792 8552 8207 8206 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08791 8215 8206 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08790 8552 8206 8215 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08789 8552 8206 8215 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08788 8215 8206 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08787 8552 8207 8013 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08786 8237 8013 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08785 8552 8013 8237 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08784 8552 8013 8237 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08783 8237 8013 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08782 8552 8207 8014 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08781 8247 8014 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08780 8552 8014 8247 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08779 8552 8014 8247 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08778 8247 8014 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08777 8552 8207 8208 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08776 8780 8208 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08775 8552 8208 8780 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08774 8552 8208 8780 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08773 8780 8208 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08772 8552 1897 1894 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08771 1815 1897 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08770 4662 1911 1815 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08769 1815 1894 4662 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08768 8552 1893 1815 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08767 1893 1911 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08766 3323 3325 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08765 3324 6365 3323 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08764 8552 3333 3324 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08763 8552 4943 4489 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08762 4489 5466 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08761 8552 5415 4489 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08760 4488 4489 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08759 8552 198 197 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08758 416 197 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08757 8552 197 416 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08756 8552 197 416 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08755 416 197 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08754 8552 416 411 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08753 5465 411 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08752 8552 411 5465 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08751 8552 411 5465 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08750 5465 411 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08749 8552 416 417 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08748 5562 417 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08747 8552 417 5562 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08746 8552 417 5562 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08745 5562 417 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08744 8552 3278 1122 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08743 1121 1122 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08742 8552 1122 1121 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08741 8552 1122 1121 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08740 1121 1122 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08739 8552 3278 1336 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08738 1335 1336 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08737 8552 1336 1335 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08736 8552 1336 1335 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08735 1335 1336 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08734 8552 3278 1337 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08733 1516 1337 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08732 8552 1337 1516 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08731 8552 1337 1516 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08730 1516 1337 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08729 8552 3278 3077 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08728 3076 3077 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08727 8552 3077 3076 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08726 8552 3077 3076 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08725 3076 3077 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08724 8552 3278 3252 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08723 3251 3252 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08722 8552 3252 3251 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08721 8552 3252 3251 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08720 3251 3252 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08719 8552 3278 3253 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08718 4057 3253 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08717 8552 3253 4057 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08716 8552 3253 4057 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08715 4057 3253 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08714 8552 3278 3114 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08713 3113 3114 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08712 8552 3114 3113 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08711 8552 3114 3113 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08710 3113 3114 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08709 1097 1463 1054 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08708 1054 1462 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08707 8552 2260 1097 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08706 2121 1097 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08705 8552 4139 1856 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08704 1856 2017 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08703 2795 3960 1856 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08702 1855 2015 2795 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08701 1856 2016 1855 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08700 8552 5440 2706 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08699 8552 8627 2708 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08698 2706 2708 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08697 8552 3880 3876 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08696 3876 3875 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08695 8552 3881 3876 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08694 3874 3876 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08693 8552 2564 2565 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08692 2565 2769 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08691 8552 2563 2565 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08690 2972 2565 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08689 8552 6873 4992 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08688 4992 5010 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08687 8552 4999 4992 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08686 6246 4992 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08685 8552 3278 3277 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08684 3276 3277 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08683 8552 3277 3276 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08682 8552 3277 3276 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08681 3276 3277 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08680 8552 3278 3279 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08679 3705 3279 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08678 8552 3279 3705 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08677 8552 3279 3705 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08676 3705 3279 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08675 8552 3330 1167 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08674 1166 1167 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08673 8552 1167 1166 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08672 8552 1167 1166 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08671 1166 1167 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08670 8552 3330 1366 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08669 1365 1366 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08668 8552 1366 1365 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08667 8552 1366 1365 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08666 1365 1366 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08665 8552 3330 1368 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08664 1367 1368 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08663 8552 1368 1367 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08662 8552 1368 1367 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08661 1367 1368 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08660 8552 3330 1200 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08659 1199 1200 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08658 8552 1200 1199 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08657 8552 1200 1199 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08656 1199 1200 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08655 8552 3330 1387 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08654 1386 1387 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08653 8552 1387 1386 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08652 8552 1387 1386 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08651 1386 1387 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08650 8552 3330 1388 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08649 2028 1388 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08648 8552 1388 2028 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08647 8552 1388 2028 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08646 2028 1388 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08645 594 597 593 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08644 595 598 594 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08643 8552 592 595 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08642 592 594 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08641 591 598 592 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08640 8552 1367 598 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08639 597 598 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08638 8552 777 596 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08637 593 596 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08636 590 589 591 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08635 8552 994 590 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08634 994 591 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08633 8552 591 994 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08632 8552 4109 1370 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08631 1370 6037 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08630 1370 4577 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08629 8552 4139 1370 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08628 1564 1370 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08627 8552 4937 4938 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08626 4936 4937 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08625 4935 4934 4936 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08624 4936 4938 4935 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08623 8552 4933 4936 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08622 4933 4934 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08621 2595 3338 2596 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08620 2594 3015 2595 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08619 8552 2593 2594 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08618 8552 1596 1440 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08617 1440 1602 2179 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08616 5945 6072 6073 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08615 5944 6352 5945 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08614 8552 6316 5944 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08613 8552 3330 3149 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08612 3148 3149 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08611 8552 3149 3148 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08610 8552 3149 3148 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08609 3148 3149 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08608 8552 3330 3303 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08607 3302 3303 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08606 8552 3303 3302 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08605 8552 3303 3302 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08604 3302 3303 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08603 8552 3330 3304 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08602 4121 3304 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08601 8552 3304 4121 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08600 8552 3304 4121 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08599 4121 3304 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08598 8552 3330 3173 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08597 3172 3173 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08596 8552 3173 3172 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08595 8552 3173 3172 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08594 3172 3173 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08593 8552 3330 3328 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08592 3327 3328 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08591 8552 3328 3327 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08590 8552 3328 3327 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08589 3327 3328 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08588 8552 3330 3331 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08587 3329 3331 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08586 8552 3331 3329 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08585 8552 3331 3329 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08584 3329 3331 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08583 8669 8672 8523 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08582 8522 8675 8669 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08581 8552 8664 8522 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08580 8664 8669 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08579 8663 8675 8664 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08578 8552 8674 8675 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08577 8672 8675 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08576 8552 8670 8673 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08575 8523 8673 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08574 8521 8520 8663 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08573 8552 8661 8521 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08572 8661 8663 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08571 8552 8663 8661 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08570 7167 8030 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08569 8552 7353 7167 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08568 7358 8030 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08567 8552 6940 7358 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08566 4130 5036 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08565 4342 6077 4130 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08564 8552 6307 4342 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08563 8552 7684 5387 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08562 5386 5387 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08561 8552 5387 5386 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08560 8552 5387 5386 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08559 5386 5387 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08558 1956 1961 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08557 1833 1959 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08556 8552 2949 1963 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08555 8552 6324 1832 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08554 1832 1963 1961 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08553 1961 2949 1833 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08552 8552 2781 2634 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08551 2635 2782 2783 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08550 2633 2787 2635 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08549 2634 3001 2633 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08548 3717 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08547 3717 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08546 8552 6285 3717 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08545 4530 3964 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08544 4530 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08543 8552 6040 4530 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08542 6364 8487 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08541 8552 8227 6364 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08540 4565 5031 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08539 8552 4754 4565 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08538 7211 7307 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08537 7305 7308 7211 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08536 8552 8417 7305 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08535 8552 7684 5591 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08534 5590 5591 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08533 8552 5591 5590 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08532 8552 5591 5590 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08531 5590 5591 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08530 8552 7684 5592 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08529 6232 5592 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08528 8552 5592 6232 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08527 8552 5592 6232 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08526 6232 5592 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08525 8552 7684 5431 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08524 5430 5431 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08523 8552 5431 5430 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08522 8552 5431 5430 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08521 5430 5431 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08520 8552 7684 5629 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08519 5628 5629 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08518 8552 5629 5628 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08517 8552 5629 5628 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08516 5628 5629 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08515 7667 7671 7600 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08514 7601 7672 7667 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08513 8552 7664 7601 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08512 7664 7667 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08511 7662 7672 7664 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08510 8552 8674 7672 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08509 7671 7672 8552 8552 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08508 8552 7669 7670 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08507 7600 7670 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08506 7599 7618 7662 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08505 8552 7660 7599 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08504 7660 7662 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08503 8552 7662 7660 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08502 1715 1716 8552 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08501 1718 1922 1714 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08500 1714 3414 8552 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08499 8552 1711 1720 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08498 1720 1712 1713 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08497 1713 1715 1718 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08496 1718 1716 1719 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08495 8552 3414 1711 8552 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08494 1710 1718 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08493 1719 1717 1720 8552 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08492 8552 7684 5630 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08491 5835 5630 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08490 8552 5630 5835 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08489 8552 5630 5835 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08488 5835 5630 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08487 8552 7684 7489 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08486 7488 7489 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08485 8552 7489 7488 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08484 8552 7489 7488 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08483 7488 7489 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08482 8552 7684 7646 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08481 7645 7646 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08480 8552 7646 7645 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08479 8552 7646 7645 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08478 7645 7646 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08477 8552 7684 7647 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08476 8596 7647 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08475 8552 7647 8596 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08474 8552 7647 8596 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08473 8596 7647 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08472 2667 2682 2608 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08471 8552 3257 2608 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08470 2608 2930 2667 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08469 2666 2667 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08468 6436 6711 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08467 8552 6878 6436 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08466 6714 6436 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08465 3716 4300 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08464 3716 4536 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08463 8552 5013 3716 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08462 8222 7147 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08461 7148 7326 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08460 8552 8430 7149 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08459 8552 7553 7146 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08458 7146 7149 7147 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08457 7147 8430 7148 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08456 3927 3756 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08455 3757 3755 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08454 8552 4747 3758 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08453 8552 4792 3754 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08452 3754 3758 3756 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08451 3756 4747 3757 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08450 6648 6738 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08449 6649 7151 8552 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08448 8552 6934 6740 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08447 8552 6739 6647 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08446 6647 6740 6738 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08445 6738 6934 6649 8552 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08444 8028 8029 7914 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08443 7914 8486 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08442 8552 8030 8028 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08441 7913 8028 8552 8552 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08440 2317 2315 8552 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08439 8552 3717 2317 8552 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08438 2321 2317 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08437 4970 5162 8552 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08436 7065 5169 4970 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08435 8552 4973 7065 8552 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08434 8787 7684 7527 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08433 7526 7527 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08432 8787 7527 7526 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08431 8787 7527 7526 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08430 7526 7527 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08429 4055 3811 3813 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08428 3813 3812 4055 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08427 8787 3809 3813 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08426 8246 7565 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08425 8787 8430 7567 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08424 7439 7723 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08423 7565 7567 7439 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08422 7438 8430 7565 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08421 8787 7987 7438 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08420 3491 4577 3492 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08419 3492 4111 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08418 3494 3490 3491 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08417 708 710 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08416 8787 988 713 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08415 712 4073 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08414 710 713 712 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08413 709 988 710 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08412 8787 926 709 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08411 6034 6032 6033 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08410 6033 6281 6035 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08409 8787 6273 6034 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08408 7297 6035 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08407 8787 7684 7683 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08406 7682 7683 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08405 8787 7683 7682 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08404 8787 7683 7682 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08403 7682 7683 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08402 8787 7684 7685 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08401 8674 7685 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08400 8787 7685 8674 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08399 8787 7685 8674 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08398 8674 7685 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08397 8787 7765 5468 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08396 5467 5468 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08395 8787 5468 5467 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08394 8787 5468 5467 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08393 5467 5468 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08392 8787 7765 5674 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08391 5673 5674 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08390 8787 5674 5673 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08389 8787 5674 5673 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08388 5673 5674 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08387 8787 7765 5675 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08386 6512 5675 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08385 8787 5675 6512 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08384 8787 5675 6512 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08383 6512 5675 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08382 8787 7765 5507 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08381 5506 5507 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08380 8787 5507 5506 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08379 8787 5507 5506 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08378 5506 5507 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08377 3427 3956 3428 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08376 3428 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08375 3426 4300 3427 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08374 3672 3425 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08373 3425 3424 3426 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08372 4085 3859 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08371 3859 3860 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08370 8787 7880 3859 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08369 3859 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08368 8787 7499 3859 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08367 8787 7757 7383 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08366 7383 7582 7384 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08365 7382 7384 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08364 3817 3835 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08363 8787 3835 3818 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08362 5371 3816 3817 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08361 3815 3818 5371 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08360 8787 3814 3815 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08359 3816 3814 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08358 8787 5180 5182 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08357 5182 5434 5181 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08356 5179 5181 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08355 8787 7765 5695 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08354 5694 5695 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08353 8787 5695 5694 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08352 8787 5695 5694 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08351 5694 5695 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08350 8787 7765 5696 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08349 6361 5696 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08348 8787 5696 6361 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08347 8787 5696 6361 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08346 6361 5696 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08345 8787 7765 7569 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08344 7568 7569 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08343 8787 7569 7568 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08342 8787 7569 7568 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08341 7568 7569 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08340 8787 7765 7728 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08339 7727 7728 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08338 8787 7728 7727 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08337 8787 7728 7727 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08336 7727 7728 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08335 8787 7765 7729 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08334 8728 7729 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08333 8787 7729 8728 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08332 8787 7729 8728 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08331 8728 7729 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08330 8787 7765 7585 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08329 7584 7585 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08328 8787 7585 7584 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08327 8787 7585 7584 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08326 7584 7585 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08325 8787 7765 7764 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08324 7763 7764 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08323 8787 7764 7763 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08322 8787 7764 7763 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08321 7763 7764 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08320 8787 7765 7766 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08319 8758 7766 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08318 8787 7766 8758 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08317 8787 7766 8758 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08316 8758 7766 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08315 8787 5465 789 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08314 789 6282 790 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08313 1011 790 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08312 8787 5471 814 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08311 814 6718 813 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08310 3295 813 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08309 808 1558 809 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08308 809 1020 810 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08307 8787 1769 808 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08306 807 810 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08305 2797 2847 2796 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08304 2796 2795 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08303 2794 4230 2797 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08302 3343 2793 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08301 2793 2792 2794 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08300 8787 8237 6216 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08299 6216 8246 6379 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08298 6378 6379 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08297 5724 6717 5725 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08296 5725 6029 5838 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08295 8787 6026 5724 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08294 6007 5838 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08293 8787 3006 2791 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08292 2791 5279 2790 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08291 2789 2790 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08290 6008 7880 6009 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08289 6009 6007 6008 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08288 8787 6027 6009 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08287 492 372 370 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08286 370 369 492 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08285 8787 1641 370 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08284 8787 6763 2258 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08283 3278 2258 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08282 8787 2258 3278 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08281 8787 2258 3278 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08280 3278 2258 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08279 8787 6763 2342 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08278 3330 2342 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08277 8787 2342 3330 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08276 8787 2342 3330 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08275 3330 2342 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08274 2469 2471 2379 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08273 2379 2482 2469 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08272 8787 2639 2379 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08271 2907 2469 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08270 481 5465 482 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08269 482 3753 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08268 480 5471 481 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08267 824 623 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08266 623 479 480 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08265 6943 7735 6942 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08264 6942 8020 6941 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08263 8787 8247 6943 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08262 6940 6941 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08261 702 700 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08260 8787 702 675 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08259 675 707 700 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08258 700 706 703 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08257 8787 1302 706 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08256 707 706 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08255 8787 704 705 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08254 703 701 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08253 699 707 702 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08252 674 706 699 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08251 8787 926 674 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08250 926 699 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08249 8787 699 926 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08248 8231 8025 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08247 7844 8490 8025 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08246 8025 8479 7845 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08245 7845 8027 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08244 8787 8242 7844 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08243 7844 8026 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08242 8358 8602 8269 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08241 8269 8355 8358 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08240 8787 8356 8269 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08239 861 994 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08238 996 1128 861 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08237 860 1129 996 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08236 8787 992 860 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08235 1338 996 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08234 8787 1123 859 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08233 859 993 996 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08232 3195 4087 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08231 5146 3265 3195 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08230 8080 8082 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08229 8787 8080 8081 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08228 8081 8083 8082 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08227 8082 8143 8140 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08226 8787 8674 8143 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08225 8083 8143 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08224 8787 8141 8142 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08223 8140 8139 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08222 8138 8083 8080 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08221 8079 8143 8138 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08220 8787 8363 8079 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08219 8363 8138 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08218 8787 8138 8363 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08217 2462 2591 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08216 2593 2592 2462 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08215 7431 7545 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08214 8741 7546 7431 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08213 7125 7127 7002 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08212 7002 7126 7125 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08211 8787 7326 7002 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08210 7124 7125 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08209 2695 2701 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08208 8787 2695 2696 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08207 2696 2703 2701 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08206 2701 2704 2702 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08205 8787 3705 2704 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08204 2703 2704 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08203 8787 2697 2700 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08202 2702 2698 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08201 2693 2703 2695 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08200 2694 2704 2693 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08199 8787 5440 2694 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08198 5440 2693 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08197 8787 2693 5440 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08196 8787 2936 2676 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08195 2676 2685 2677 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08194 2675 2677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08193 1794 1783 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_08192 8787 1988 1794 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_08191 1794 2343 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_08190 8787 1781 1794 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_08189 1466 2255 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08188 1465 2127 1466 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08187 8787 1956 1465 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08186 1717 1465 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08185 8787 2481 2033 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08184 2033 5150 2111 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08183 2235 2111 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08182 8225 8222 8224 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08181 8224 8223 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08180 8226 8780 8225 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08179 5461 5211 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08178 5210 5215 5211 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08177 5211 5209 5213 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08176 5213 5212 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08175 8787 5363 5210 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08174 5210 5214 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08173 2445 2576 2444 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08172 2444 2771 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08171 2773 3317 2445 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08170 7365 7579 7366 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08169 7366 7734 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08168 7364 7367 7365 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08167 7012 7573 7013 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08166 7013 7357 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08165 7164 7167 7012 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08164 6554 7404 6555 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08163 6555 8487 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08162 6552 8030 6554 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08161 6553 8240 6552 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08160 8234 8231 8233 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08159 8233 8232 8234 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08158 8787 8473 8233 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08157 8467 8234 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08156 3338 3339 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08155 8787 3551 3339 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08154 3339 3544 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08153 8787 3525 3339 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08152 7448 8098 7449 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08151 7449 8020 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08150 7578 8780 7448 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08149 8787 8019 7039 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08148 7039 7770 7183 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08147 7182 7183 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08146 8787 185 186 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08145 3320 186 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08144 8787 186 3320 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08143 8787 186 3320 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08142 3320 186 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08141 8787 3320 3321 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08140 6026 3321 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08139 8787 3321 6026 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08138 8787 3321 6026 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08137 6026 3321 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08136 8787 3320 1029 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08135 6021 1029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08134 8787 1029 6021 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08133 8787 1029 6021 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08132 6021 1029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08131 8787 3320 3161 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08130 6716 3161 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08129 8787 3161 6716 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08128 8787 3161 6716 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08127 6716 3161 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08126 8787 3320 3162 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08125 6284 3162 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08124 8787 3162 6284 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08123 8787 3162 6284 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08122 6284 3162 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08121 8787 3320 819 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08120 4300 819 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08119 8787 819 4300 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08118 8787 819 4300 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08117 4300 819 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08116 6937 7353 6939 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08115 6939 7576 6938 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08114 8787 7592 6937 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08113 6936 6938 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08112 8787 8455 8295 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08111 8295 8454 8456 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08110 8746 8456 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08109 8787 638 635 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08108 1044 635 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08107 8787 635 1044 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08106 8787 635 1044 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08105 1044 635 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08104 8787 1044 1045 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08103 3333 1045 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08102 8787 1045 3333 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08101 8787 1045 3333 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08100 3333 1045 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08099 8787 1044 634 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08098 4139 634 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08097 8787 634 4139 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08096 8787 634 4139 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08095 4139 634 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08094 7240 7228 6802 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08093 8787 8350 6803 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08092 6802 6803 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08091 6333 6335 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08090 8787 6333 6190 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08089 6190 6336 6335 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08088 6335 6338 6192 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08087 8787 6512 6338 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08086 6336 6338 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08085 8787 6191 6337 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08084 6192 6218 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08083 6332 6336 6333 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08082 6189 6338 6332 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08081 8787 6514 6189 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08080 6514 6332 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08079 8787 6332 6514 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08078 2095 2182 2096 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08077 2096 2183 2184 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08076 8787 2789 2095 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08075 2582 2184 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08074 3217 3297 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_08073 6873 3531 3217 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_08072 3216 6021 6873 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_08071 8787 3294 3216 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_08070 3216 3295 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_08069 6493 6494 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08068 8787 6493 6495 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08067 6495 6501 6494 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08066 6494 6500 6496 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08065 8787 6512 6500 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08064 6501 6500 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08063 8787 6497 6499 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08062 6496 6498 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08061 6492 6501 6493 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08060 6491 6500 6492 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08059 8787 6925 6491 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08058 6925 6492 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08057 8787 6492 6925 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08056 2711 2713 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08055 2712 2942 2713 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08054 2713 2949 2714 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08053 2714 5676 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08052 8787 2947 2712 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08051 2712 2715 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08050 1269 4109 1270 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08049 1270 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08048 1268 3964 1269 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08047 1591 1380 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08046 1380 1278 1268 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08045 1873 6717 1872 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08044 1872 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08043 1871 3964 1873 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08042 2008 2006 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08041 2006 2007 1871 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08040 2863 2949 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08039 2944 5220 2863 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08038 3773 4157 3632 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08037 3632 5915 3773 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08036 8787 3775 3632 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08035 4981 6279 4866 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08034 4866 6860 4981 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08033 8787 4990 4866 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08032 5170 4981 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08031 3558 3648 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08030 3827 3644 3558 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08029 5623 8110 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08028 5625 5621 5623 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08027 8787 5843 5620 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08026 5620 6283 5625 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08025 8787 5826 5622 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08024 5622 5844 5625 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08023 392 2974 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08022 391 6077 392 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08021 2375 2596 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08020 2376 2374 2375 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08019 2882 3342 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08018 3015 3181 2882 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08017 6772 8478 6605 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08016 6605 6972 6772 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08015 8787 6970 6605 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08014 6674 6772 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08013 5354 7404 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08012 5505 6940 5354 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08011 5277 8764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08010 5275 5284 5277 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08009 8787 3275 2047 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08008 2047 2139 2136 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08007 2270 2136 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08006 8787 7294 7287 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08005 7287 7285 7286 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08004 8131 7286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08003 6832 8235 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08002 6964 8780 6832 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08001 1255 3898 1254 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08000 1254 6037 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07999 1772 3531 1255 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07998 7121 6720 6574 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07997 6574 6873 7121 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07996 8787 6719 6574 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07995 8787 1496 1104 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07994 1104 1318 1103 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07993 1310 1103 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07992 6024 6286 6025 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07991 6025 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07990 6023 6021 6024 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07989 6883 6022 6023 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07988 1168 2964 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07987 1215 2723 1168 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07986 307 310 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07985 8787 988 311 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07984 309 3680 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07983 310 311 309 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07982 308 988 310 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07981 8787 555 308 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07980 986 989 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07979 8787 988 991 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07978 772 2718 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07977 989 991 772 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07976 771 988 989 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07975 8787 993 771 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07974 3074 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07973 3648 3073 3074 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07972 3072 3246 3648 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07971 8787 3655 3072 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07970 3072 3646 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07969 4898 5562 4897 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07968 4897 5013 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07967 4896 6284 4898 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07966 5014 6758 4896 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07965 3011 2777 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07964 8787 3000 2777 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07963 2777 2775 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07962 8787 2776 2777 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07961 6601 7752 6670 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07960 6670 6770 6601 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07959 8787 6769 6601 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07958 6601 6955 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07957 4852 4943 4851 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07956 4851 5851 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07955 4850 5466 4852 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07954 4944 5415 4850 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07953 944 947 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07952 8787 1525 948 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07951 739 3849 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07950 947 948 739 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07949 738 1525 947 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07948 8787 1105 738 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07947 1286 1086 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07946 8787 1525 1089 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07945 1088 4073 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07944 1086 1089 1088 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07943 1087 1525 1086 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07942 8787 1280 1087 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07941 975 976 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07940 8787 988 978 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07939 756 2284 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07938 976 978 756 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07937 754 988 976 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07936 8787 1125 754 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07935 7304 7307 7303 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07934 7303 7308 7304 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07933 8787 7326 7303 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07932 8787 3414 1474 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07931 1472 1716 1470 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07930 1475 1915 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_07929 1470 1469 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07928 1474 1477 1471 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07927 1471 1915 1472 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07926 1472 1475 1473 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07925 2119 1472 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07924 8787 3414 1469 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_07923 1473 1732 1474 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07922 2339 2337 2344 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07921 2344 2890 2339 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07920 8787 2338 2339 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07919 2339 6307 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07918 8787 1138 1136 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07917 1136 1135 1137 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07916 3469 1137 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07915 8787 5645 5627 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07914 5627 5625 5626 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07913 5624 5626 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07912 8485 8782 8306 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07911 8306 8483 8485 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07910 8787 8780 8306 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07909 6267 7320 6159 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07908 6159 6276 6267 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07907 8787 6721 6159 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07906 6265 6267 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07905 434 548 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07904 540 1128 434 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07903 433 1129 540 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07902 8787 542 433 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07901 2504 540 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07900 8787 1123 432 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07899 432 538 540 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07898 6241 6243 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07897 6148 7535 6243 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07896 6243 6242 6147 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07895 6147 6420 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07894 8787 7536 6148 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07893 6148 7533 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07892 4394 4943 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07891 8787 4943 4497 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07890 4499 4495 4394 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07889 4393 4497 4499 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07888 8787 5466 4393 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07887 4495 5466 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07886 8787 8247 7007 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07885 7007 8020 7150 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07884 7151 7150 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07883 8465 8466 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07882 8787 8465 8298 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07881 8298 8470 8466 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07880 8466 8471 8300 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07879 8787 8758 8471 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07878 8470 8471 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07877 8787 8299 8468 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07876 8300 8313 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07875 8463 8470 8465 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07874 8297 8471 8463 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07873 8787 8461 8297 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07872 8461 8463 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07871 8787 8463 8461 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07870 2261 2274 2262 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07869 2262 2273 2261 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07868 8787 2260 2262 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07867 3262 2261 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07866 418 5470 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07865 8787 1203 418 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07864 6235 6237 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07863 6145 7535 6237 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07862 6237 6238 6146 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07861 6146 6415 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07860 8787 7536 6145 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07859 6145 7533 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07858 7087 6433 6434 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07857 6434 6873 7087 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07856 8787 6432 6434 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07855 3913 3912 3914 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07854 3914 3915 3913 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07853 8787 8627 3914 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07852 4217 3913 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07851 1560 4530 1559 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07850 1559 2305 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07849 1557 2159 1560 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07848 1558 1556 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07847 1556 1555 1557 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07846 6106 6107 6105 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07845 6105 6115 6106 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07844 8787 6104 6105 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07843 7939 7940 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07842 8787 7939 7789 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07841 7789 7942 7940 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07840 7940 7944 7791 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07839 8787 8674 7944 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07838 7942 7944 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07837 8787 7790 7943 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07836 7791 7867 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07835 7934 7942 7939 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07834 7788 7944 7934 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07833 8787 7937 7788 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07832 7937 7934 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07831 8787 7934 7937 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07830 8787 8341 8599 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07829 8341 8586 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07828 8599 8350 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07827 7701 7705 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07826 8787 7701 7704 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07825 7704 7709 7705 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07824 7705 7710 7703 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07823 8787 8728 7710 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07822 7709 7710 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07821 8787 7706 7708 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07820 7703 7702 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07819 7700 7709 7701 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07818 7699 7710 7700 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07817 8787 7716 7699 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07816 7716 7700 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07815 8787 7700 7716 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07814 3841 5388 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07813 5601 3840 3841 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07812 8004 7904 7733 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07811 7733 7731 8004 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07810 8787 7732 7733 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07809 8050 8049 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07808 8315 8627 8050 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07807 6469 6474 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07806 8787 6469 6470 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07805 6470 6476 6474 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07804 6474 6478 6475 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07803 8787 6512 6478 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07802 6476 6478 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07801 8787 6471 6477 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07800 6475 6472 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07799 6467 6476 6469 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07798 6468 6478 6467 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07797 8787 6466 6468 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07796 6466 6467 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07795 8787 6467 6466 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07794 8787 4469 3556 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07793 3556 3639 3640 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07792 3812 3640 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07791 3857 6720 3858 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07790 3858 5408 3857 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07789 8787 6268 3858 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07788 8787 6077 1631 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07787 1631 2151 1762 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07786 1959 1762 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07785 8787 4799 4332 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07784 4332 4773 4331 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07783 4330 4331 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07782 8787 6254 6017 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07781 6017 6432 6016 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07780 6439 6016 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07779 8290 8764 8723 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07778 8787 8764 8449 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07777 8291 8446 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07776 8723 8449 8291 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07775 8787 8445 8290 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07774 2826 3956 2827 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07773 2827 6718 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07772 2825 6716 2826 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07771 2937 5826 2825 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07770 8130 8128 8129 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07769 8129 8132 8130 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07768 8787 8127 8129 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07767 8355 8130 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07766 8787 631 632 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07765 631 2566 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07764 632 1390 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07763 1997 822 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07762 822 823 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07761 8787 824 822 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07760 8787 8775 8777 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07759 8777 8778 8779 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07758 8776 8779 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07757 1460 1725 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07756 8787 1725 1461 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07755 1897 1458 1460 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07754 1459 1461 1897 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07753 8787 1723 1459 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07752 1458 1723 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07751 5186 2248 2249 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07750 2249 2247 5186 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07749 8787 2723 2249 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07748 4008 5563 4009 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07747 4009 5562 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07746 6077 6716 4008 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07745 3005 3004 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07744 8787 2897 3004 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07743 3004 3539 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07742 8787 3535 3004 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07741 7786 8627 8185 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07740 8787 8627 7931 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07739 7785 8121 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07738 8185 7931 7785 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07737 8787 8585 7786 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07736 8787 4971 4705 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07735 4705 4961 4704 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07734 4703 4704 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07733 4095 4094 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07732 4094 4040 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07731 8787 7880 4094 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07730 4094 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07729 8787 7877 4094 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07728 8787 4085 3994 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07727 3994 5606 4086 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07726 4087 4086 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07725 8787 2572 2431 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07724 2431 2548 2549 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07723 2550 2549 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07722 8787 5641 5635 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07721 5635 5848 5636 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07720 5634 5636 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07719 8787 4109 2428 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07718 2428 6037 2546 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07717 3133 2546 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07716 3244 3552 3245 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07715 3245 3343 3344 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07714 8787 4237 3244 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07713 3342 3344 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07712 4317 6282 4316 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07711 4316 4536 4315 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07710 8787 6716 4317 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07709 5644 4315 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07708 8787 4158 4159 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07707 4374 4159 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07706 8787 4159 4374 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07705 8787 4159 4374 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07704 4374 4159 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07703 8787 4374 3908 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07702 8135 3908 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07701 8787 3908 8135 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07700 8787 3908 8135 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07699 8135 3908 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07698 8787 4374 3909 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07697 8627 3909 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07696 8787 3909 8627 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07695 8787 3909 8627 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07694 8627 3909 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07693 8787 4374 4375 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07692 8350 4375 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07691 8787 4375 8350 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07690 8787 4375 8350 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07689 8350 4375 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07688 8787 4374 4136 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07687 8065 4136 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07686 8787 4136 8065 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07685 8787 4136 8065 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07684 8065 4136 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07683 2989 2992 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07682 8787 2989 2842 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07681 2842 2994 2992 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07680 2992 2995 2843 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07679 8787 3329 2995 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07678 2994 2995 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07677 8787 2876 2993 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07676 2843 2892 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07675 2988 2994 2989 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07674 2841 2995 2988 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07673 8787 2986 2841 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07672 2986 2988 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07671 8787 2988 2986 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07670 3651 3389 3391 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07669 3391 3390 3651 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07668 8787 3388 3391 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07667 6269 7073 6160 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07666 6160 6276 6269 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07665 8787 6719 6160 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07664 6268 6269 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07663 8787 5470 52 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07662 52 1203 199 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07661 198 199 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07660 4849 5124 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07659 8787 5124 4942 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07658 4941 4939 4849 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07657 4848 4942 4941 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07656 8787 5130 4848 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07655 4939 5130 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07654 127 128 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07653 8787 127 28 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07652 28 133 128 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07651 128 134 30 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07650 8787 1516 134 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07649 133 134 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07648 8787 29 132 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07647 30 130 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07646 125 133 127 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07645 27 134 125 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07644 8787 560 27 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07643 560 125 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07642 8787 125 560 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07641 1646 3717 1777 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07640 1777 2890 1646 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07639 8787 1775 1646 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07638 1646 2159 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07637 1599 1202 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07636 8787 1201 1599 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07635 903 3898 904 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07634 904 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07633 902 5013 903 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07632 1201 1042 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07631 1042 901 902 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07630 2130 2517 2044 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07629 2044 2707 2130 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07628 8787 2129 2044 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07627 2128 2130 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07626 1266 3753 1267 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07625 1267 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07624 1265 5471 1266 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07623 1790 1377 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07622 1377 1277 1265 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07621 8090 8091 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07620 8787 8090 8092 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07619 8092 8093 8091 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07618 8091 8159 8157 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07617 8787 8674 8159 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07616 8093 8159 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07615 8787 8155 8158 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07614 8157 8156 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07613 8154 8093 8090 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07612 8089 8159 8154 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07611 8787 8160 8089 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07610 8160 8154 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07609 8787 8154 8160 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07608 4231 6537 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07607 4230 5280 4231 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07606 3507 3750 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07605 8787 3750 3506 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07604 8787 5790 3504 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07603 3505 3503 3507 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07602 3504 3506 3505 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07601 3502 3505 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07600 8787 3505 3502 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07599 3503 5790 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07598 7348 7347 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07597 7570 7345 7348 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07596 5553 6307 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07595 5668 6077 5553 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07594 4398 7315 4399 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07593 4399 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07592 4503 4501 4398 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07591 2271 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07590 2272 2270 2271 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07589 2269 2267 2272 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07588 8787 3655 2269 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07587 2269 2268 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07586 1951 1757 1629 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07585 1629 1758 1951 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07584 8787 2260 1629 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07583 8787 2127 1891 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07582 1891 2255 1892 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07581 1890 1892 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07580 3586 3716 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07579 3715 3717 3586 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07578 8787 3860 3715 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07577 3875 3715 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07576 3680 3682 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07575 8787 4075 3684 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07574 3575 4281 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07573 3682 3684 3575 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07572 3574 4075 3682 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07571 8787 8417 3574 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07570 4870 5557 4869 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07569 4869 5438 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07568 7643 4988 4870 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07567 8787 8364 8366 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07566 8364 8363 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07565 8366 8627 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07564 7043 8781 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07563 7185 8780 7043 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07562 2332 6717 2333 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07561 2333 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07560 2337 3753 2332 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07559 4757 6029 4756 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07558 4756 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07557 4988 6026 4757 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07556 3910 6717 3911 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07555 3911 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07554 4984 6026 3910 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07553 1141 1144 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07552 8787 1525 1146 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07551 1143 2718 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07550 1144 1146 1143 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07549 1142 1525 1144 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07548 8787 1140 1142 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07547 5427 5171 5167 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07546 5167 5166 5427 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07545 8787 8065 5167 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07544 8787 3414 2394 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07543 2497 2500 2392 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07542 2492 2498 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_07541 2392 2493 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07540 2394 2670 2393 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07539 2393 2498 2497 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07538 2497 2492 2395 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07537 2671 2497 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07536 8787 3414 2493 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_07535 2395 2930 2394 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07534 2343 2004 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07533 2004 2005 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07532 8787 2008 2004 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07531 1633 3956 1632 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07530 1632 6718 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07529 4532 6284 1633 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07528 937 734 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07527 8787 779 735 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07526 733 4073 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07525 734 735 733 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07524 732 779 734 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07523 8787 931 732 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07522 1513 1343 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07521 8787 1525 1345 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07520 1244 2284 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07519 1343 1345 1244 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07518 1243 1525 1343 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07517 8787 1505 1243 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07516 960 963 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07515 8787 1525 964 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07514 750 3680 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07513 963 964 750 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07512 748 1525 963 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07511 8787 959 748 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07510 5769 7184 5770 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07509 5770 7353 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07508 5768 6677 5769 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07507 5919 8490 5768 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07506 5336 7592 5335 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07505 5335 6673 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07504 5334 6940 5336 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07503 5915 8490 5334 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07502 1642 3767 1643 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07501 1643 4109 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07500 2160 3956 1642 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07499 550 551 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07498 8787 779 552 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07497 438 3849 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07496 551 552 438 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07495 437 779 551 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07494 8787 548 437 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07493 4762 4999 4761 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07492 4761 6307 4760 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07491 8787 6077 4762 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07490 5212 4760 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07489 1666 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07488 1738 1741 1666 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07487 1665 1926 1738 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07486 8787 3655 1665 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07485 1665 1923 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07484 7540 7109 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07483 7109 8128 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07482 8787 7880 7109 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07481 7109 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07480 8787 7877 7109 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07479 8787 8135 2736 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07478 2736 2746 2735 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07477 2734 2735 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07476 8787 8019 5756 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07475 5756 6368 5913 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07474 5912 5913 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07473 8787 3460 3461 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07472 3861 3461 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07471 8787 3461 3861 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07470 8787 3461 3861 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07469 3861 3461 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07468 8787 3861 3862 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07467 7499 3862 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07466 8787 3862 7499 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07465 8787 3862 7499 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07464 7499 3862 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07463 8787 3861 3708 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07462 7877 3708 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07461 8787 3708 7877 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07460 8787 3708 7877 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07459 7877 3708 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07458 8787 6095 6096 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07457 6096 8764 6097 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07456 6761 6097 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07455 6850 7228 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07454 6849 7643 6850 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07453 8787 6861 6849 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07452 7251 6849 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07451 8787 5465 3487 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07450 3487 3956 3486 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07449 3744 3486 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07448 319 322 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07447 8787 319 320 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07446 320 327 322 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07445 322 326 321 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07444 8787 1516 326 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07443 327 326 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07442 8787 323 325 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07441 321 324 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07440 318 327 319 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07439 317 326 318 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07438 8787 765 317 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07437 765 318 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07436 8787 318 765 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07435 1661 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07434 1725 1907 1661 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07433 1660 1902 1725 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07432 8787 3655 1660 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07431 1660 1723 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07430 8620 8622 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07429 8621 8624 8620 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07428 8787 8618 8621 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07427 8619 8621 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07426 49 2974 50 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07425 50 805 180 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07424 8787 5033 49 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07423 179 180 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07422 1673 2572 1674 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07421 1674 4792 1770 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07420 8787 2334 1673 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07419 1769 1770 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07418 7644 8572 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07417 7642 7643 7644 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07416 8787 7641 7642 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07415 8323 7642 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07414 282 285 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07413 8787 282 286 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07412 286 288 285 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07411 285 290 284 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07410 8787 1302 290 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07409 288 290 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07408 8787 287 289 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07407 284 283 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07406 281 288 282 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07405 280 290 281 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07404 8787 538 280 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07403 538 281 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07402 8787 281 538 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07401 2908 2907 2808 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07400 2808 2911 2908 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07399 8787 2906 2808 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07398 3826 2908 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07397 3240 5471 3241 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07396 3241 5562 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07395 3239 4300 3240 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07394 5280 3332 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07393 3332 3238 3239 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07392 4914 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07391 5044 5043 4914 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07390 4913 5280 5044 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07389 8787 6957 4913 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07388 4913 8023 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07387 8608 8609 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07386 8787 8608 8610 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07385 8610 8615 8609 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07384 8609 8616 8613 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07383 8787 8674 8616 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07382 8615 8616 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07381 8787 8611 8614 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07380 8613 8612 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07379 8607 8615 8608 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07378 8606 8616 8607 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07377 8787 8605 8606 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07376 8605 8607 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07375 8787 8607 8605 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07374 1529 1771 1530 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07373 1530 1537 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07372 2260 1763 1529 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07371 7536 2986 367 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07370 8787 1567 368 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07369 367 368 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07368 8251 8323 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07367 8569 8326 8251 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07366 4025 4061 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07365 4206 4646 4025 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07364 2042 3490 2043 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07363 2043 6718 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07362 2041 4300 2042 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07361 2127 7049 2041 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07360 8787 2936 2810 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07359 2810 3085 2914 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07358 3246 2914 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07357 372 1567 371 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07356 8787 2986 373 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07355 371 373 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07354 4026 4690 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07353 4083 4079 4026 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07352 7974 7697 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07351 8787 8394 7698 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07350 7696 8741 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07349 7697 7698 7696 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07348 7695 8394 7697 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07347 8787 7969 7695 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07346 8655 8379 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07345 8787 8394 8381 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07344 8153 8688 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07343 8379 8381 8153 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07342 8149 8394 8379 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07341 8787 8648 8149 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07340 7515 7517 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07339 8787 8394 7519 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07338 7424 8646 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07337 7517 7519 7424 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07336 7423 8394 7517 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07335 8787 7514 7423 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07334 8787 6878 6451 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07333 6451 6719 6452 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07332 6453 6452 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07331 4432 4577 4433 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07330 4433 6717 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07329 4431 5562 4432 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07328 4787 4561 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07327 4561 4430 4431 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07326 8787 414 415 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07325 414 5470 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07324 415 1203 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07323 5407 6872 5306 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07322 5306 5408 5407 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07321 8787 6262 5306 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07320 5406 5407 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07319 8787 5036 3517 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07318 3517 4139 3518 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07317 3516 3518 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07316 5286 5290 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07315 8787 5286 5289 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07314 5289 5294 5290 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07313 5290 5295 5288 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07312 8787 6361 5295 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07311 5294 5295 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07310 8787 5291 5293 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07309 5288 5287 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07308 5285 5294 5286 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07307 5283 5295 5285 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07306 8787 5284 5283 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07305 5284 5285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07304 8787 5285 5284 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07303 2348 2346 2347 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07302 2347 2567 2349 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07301 8787 3317 2348 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07300 2587 2349 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07299 7117 7118 7001 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07298 7001 7115 7117 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07297 8787 8648 7001 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07296 7116 7117 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07295 8787 7921 7855 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07294 7921 8110 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07293 7855 8135 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07292 5961 5965 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07291 8787 5961 5964 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07290 5964 5968 5965 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07289 5965 5970 5963 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07288 8787 6232 5970 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07287 5968 5970 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07286 8787 5967 5969 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07285 5963 5962 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07284 5960 5968 5961 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07283 5959 5970 5960 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07282 8787 5958 5959 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07281 5958 5960 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07280 8787 5960 5958 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07279 6823 6825 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07278 8787 6823 6824 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07277 6824 6826 6825 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07276 6825 6918 6915 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07275 8787 8728 6918 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07274 6826 6918 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07273 8787 6916 6917 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07272 6915 6914 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07271 6911 6826 6823 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07270 6822 6918 6911 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07269 8787 7329 6822 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07268 7329 6911 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07267 8787 6911 7329 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07266 1234 3254 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07265 1496 3673 1234 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07264 7676 7875 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07263 7677 7874 7676 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07262 8787 7675 7677 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07261 7951 7677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07260 3243 3553 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07259 3341 3776 3243 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07258 4218 4217 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07257 8423 4553 4218 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07256 4412 4529 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07255 5776 4530 4412 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07254 8774 8782 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07253 8775 8780 8774 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07252 3607 6029 3606 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07251 3606 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07250 6307 3753 3607 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07249 333 336 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07248 8787 983 337 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07247 335 3709 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07246 336 337 335 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07245 334 983 336 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07244 8787 764 334 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07243 5264 8764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07242 5265 5263 5264 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07241 5566 8764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07240 5684 5565 5566 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07239 6030 6029 6031 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07238 6031 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07237 6028 6026 6030 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07236 6446 6027 6028 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07235 8787 1951 1953 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07234 1953 5183 1955 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07233 1952 1955 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07232 8787 3269 1909 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07231 1909 2508 1908 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07230 1907 1908 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07229 3540 4153 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07228 3539 4148 3540 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07227 7655 7937 7654 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07226 8787 8135 7656 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07225 7654 7656 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07224 4951 4698 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07223 4696 7535 4698 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07222 4698 4697 4699 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07221 4699 4723 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07220 8787 7536 4696 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07219 4696 7533 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07218 980 982 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07217 8787 983 984 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07216 763 2284 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07215 982 984 763 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07214 762 983 982 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07213 8787 1124 762 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07212 7271 7658 7272 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07211 7272 8132 7271 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07210 8787 7657 7272 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07209 7929 7271 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07208 8266 8349 8267 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07207 8267 8348 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07206 8265 8346 8266 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07205 8602 8347 8265 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07204 2853 3678 2852 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07203 2852 3677 2932 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07202 8787 7723 2853 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07201 2931 2932 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07200 6163 6286 6162 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07199 6162 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07198 6161 6284 6163 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07197 6438 6271 6161 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07196 1753 1758 1628 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07195 1628 1757 1753 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07194 8787 2723 1628 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07193 2844 3326 2845 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07192 2845 2999 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07191 3000 2998 2844 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07190 5180 7880 5168 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07189 5168 6007 5180 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07188 8787 6283 5168 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07187 2075 4530 2074 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07186 2074 4792 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07185 2073 2572 2075 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07184 2745 2159 2073 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07183 680 565 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07182 8787 779 567 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07181 445 2284 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07180 565 567 445 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07179 444 779 565 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07178 8787 1127 444 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07177 559 563 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07176 8787 779 564 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07175 443 3680 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07174 563 564 443 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07173 442 779 563 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07172 8787 560 442 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07171 7081 7257 6994 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07170 8787 8065 7082 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07169 6994 7082 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07168 715 718 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07167 8787 983 719 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07166 717 4073 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07165 718 719 717 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07164 716 983 718 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07163 8787 925 716 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07162 4406 4714 4407 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07161 4407 4520 4521 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07160 8787 4518 4406 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07159 4519 4521 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07158 8787 4095 3996 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07157 3996 5824 4093 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07156 4092 4093 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07155 5120 5790 5121 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07154 5121 6290 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07153 5118 5466 5120 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07152 5119 5415 5118 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07151 8457 8226 8221 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07150 8221 8220 8457 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07149 8787 8454 8221 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07148 8787 1522 1519 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07147 1519 5214 1520 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07146 1757 1520 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07145 7741 7743 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07144 7742 8220 7743 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07143 7743 8235 7744 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07142 7744 8247 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07141 8787 8455 7742 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07140 7742 7746 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07139 8787 4792 2434 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_07138 2434 3048 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_07137 2569 2562 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07136 2434 6878 2562 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_07135 2562 2890 2434 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_07134 3271 4502 3200 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07133 3200 5408 3271 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07132 8787 4096 3200 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07131 3888 6040 3890 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07130 3890 4536 3889 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07129 8787 3964 3888 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07128 4075 3889 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07127 364 1016 365 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07126 365 7536 364 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07125 8787 6077 365 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07124 363 364 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07123 4227 4229 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07122 8787 4227 4228 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07121 4228 4362 4229 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07120 4229 4364 4360 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07119 8787 6361 4364 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07118 4362 4364 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07117 8787 4361 4363 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07116 4360 4359 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07115 4357 4362 4227 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07114 4226 4364 4357 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07113 8787 4358 4226 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07112 4358 4357 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07111 8787 4357 4358 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07110 724 726 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07109 725 1128 724 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07108 723 1129 725 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07107 8787 720 723 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07106 2252 725 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07105 8787 1123 722 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07104 722 721 725 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07103 6958 8490 6959 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07102 6959 7761 6960 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07101 8787 8240 6958 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07100 6957 6960 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07099 5357 6940 5358 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07098 5358 6673 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07097 5356 7184 5357 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07096 5508 5509 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07095 5509 5355 5356 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07094 7326 7073 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07093 8417 8202 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07092 404 3490 405 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07091 405 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07090 403 5192 404 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07089 499 402 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07088 402 401 403 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07087 6249 6247 6149 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07086 6149 6246 6249 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07085 8787 7076 6149 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07084 6245 6249 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07083 3866 3469 3464 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07082 3464 3462 3866 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07081 8787 4092 3464 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07080 6891 7127 6892 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07079 6892 7126 6891 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07078 8787 7142 6892 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07077 7088 6891 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07076 8075 8077 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07075 8787 8075 8076 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07074 8076 8078 8077 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07073 8077 8126 8125 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07072 8787 8674 8126 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07071 8078 8126 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07070 8787 8122 8124 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07069 8125 8123 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07068 8120 8078 8075 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07067 8074 8126 8120 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07066 8787 8121 8074 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07065 8121 8120 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07064 8787 8120 8121 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07063 1497 1498 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07062 1747 1496 1497 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07061 4098 8185 3997 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07060 3997 6276 4098 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07059 8787 4099 3997 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07058 4096 4098 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07057 7826 3472 3470 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07056 3470 3469 7826 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07055 8787 3718 3470 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07054 1145 3898 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07053 7533 6717 1145 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07052 1865 4979 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07051 2148 1954 1865 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07050 7989 7988 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07049 8787 7989 7807 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07048 7807 7993 7988 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07047 7988 7995 7809 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07046 8787 8728 7995 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07045 7993 7995 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07044 8787 7808 7992 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07043 7809 7898 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07042 7984 7993 7989 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07041 7806 7995 7984 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07040 8787 7987 7806 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07039 7987 7984 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07038 8787 7984 7987 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07037 1637 4577 1636 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07036 1636 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07035 1966 2566 1637 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07034 6888 7315 6890 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07033 6890 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07032 6887 8372 6888 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07031 3335 5510 3242 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07030 3242 3334 3335 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07029 8787 3333 3242 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07028 2686 2927 2687 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07027 2687 2933 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07026 2684 3082 2686 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07025 2685 3083 2684 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07024 8787 3429 3402 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07023 3402 3400 3401 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07022 3658 3401 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07021 4389 5466 4390 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07020 4390 4943 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07019 4487 5415 4389 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07018 5600 5604 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07017 8787 8394 5605 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07016 5603 5601 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07015 5604 5605 5603 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07014 5602 8394 5604 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07013 8787 6000 5602 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07012 5402 5147 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07011 8787 8394 5149 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07010 5148 5146 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07009 5147 5149 5148 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07008 5145 8394 5147 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07007 8787 6251 5145 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07006 4215 4082 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07005 8787 8394 4084 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07004 3993 4083 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07003 4082 4084 3993 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07002 3992 8394 4082 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07001 8787 5998 3992 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07000 1933 2937 1932 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06999 1932 2277 1934 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06998 8787 3657 1933 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06997 1931 1934 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06996 1662 3269 1663 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06995 1663 2508 1730 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06994 8787 3657 1662 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06993 1729 1730 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06992 1532 6718 1531 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06991 1531 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06990 1768 3136 1532 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06989 1256 3753 1257 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06988 1257 4109 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06987 1546 1369 1256 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06986 8787 2334 2335 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06985 2335 2890 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06984 3318 2336 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06983 2335 2337 2336 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06982 2336 3048 2335 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06981 2881 5279 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06980 3007 3006 2881 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06979 5142 7880 5144 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06978 5144 6007 5142 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06977 8787 6271 5144 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06976 2293 2147 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06975 8787 8394 2150 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06974 1962 2148 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06973 2147 2150 1962 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06972 1958 8394 2147 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06971 8787 5188 1958 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06970 3199 3956 3198 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06969 3198 6286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06968 3197 6284 3199 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06967 3269 6708 3197 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06966 3049 2971 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06965 8787 2890 2971 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06964 2971 3314 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06963 8787 3315 2971 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06962 8787 1297 1222 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06961 1222 5214 1298 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06960 2251 1298 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06959 8787 3956 2737 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06958 2737 6286 2738 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06957 3297 2738 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06956 8787 4577 2768 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06955 2768 2784 2767 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06954 3164 2767 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06953 8787 8780 6974 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06952 6974 8483 6973 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06951 6972 6973 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06950 5994 5996 5995 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06949 5995 6246 5994 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06948 8787 6241 5995 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06947 5993 5994 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06946 3723 7118 3591 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06945 3591 7115 3723 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06944 8787 4522 3591 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06943 1206 1210 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06942 8787 1206 1207 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06941 1207 1212 1210 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06940 1210 1214 1211 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06939 8787 2028 1214 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06938 1212 1214 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06937 8787 1208 1213 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06936 1211 1209 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06935 1204 1212 1206 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06934 1205 1214 1204 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06933 8787 1203 1205 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06932 1203 1204 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06931 8787 1204 1203 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06930 5766 5915 5767 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06929 5767 5919 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06928 5765 5916 5766 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06927 6123 5918 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06926 5918 5764 5765 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06925 2171 1995 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06924 8787 1996 2171 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06923 5672 5669 5671 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06922 5671 5668 5672 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06921 8787 5666 5671 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06920 5856 5672 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06919 753 752 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06918 8787 753 679 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06917 679 759 752 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06916 752 761 757 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06915 8787 1516 761 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06914 759 761 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06913 8787 758 760 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06912 757 755 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06911 751 759 753 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06910 678 761 751 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06909 8787 1127 678 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06908 1127 751 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06907 8787 751 1127 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06906 2265 2511 2264 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06905 2264 2263 2265 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06904 8787 2936 2264 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06903 2267 2265 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06902 3234 6286 3235 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06901 3235 3749 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06900 3233 6282 3234 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06899 3334 3322 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06898 3322 3232 3233 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06897 2170 1791 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06896 8787 1790 2170 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06895 1178 5470 1179 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06894 1179 1203 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06893 1176 1390 1178 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06892 2784 1177 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06891 1177 1175 1176 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06890 5545 5547 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06889 8787 5545 5546 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06888 5546 5598 5547 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06887 5547 5599 5596 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06886 8787 6232 5599 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06885 5598 5599 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06884 8787 5594 5597 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06883 5596 5595 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06882 5593 5598 5545 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06881 5544 5599 5593 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06880 8787 6000 5544 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06879 6000 5593 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06878 8787 5593 6000 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06877 1866 2151 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06876 2537 6077 1866 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06875 3839 4693 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06874 5580 3838 3839 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06873 2099 2372 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06872 2191 2374 2099 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06871 362 360 361 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06870 361 363 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06869 599 609 362 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06868 4212 4213 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06867 8787 4212 4214 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06866 4214 4275 4213 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06865 4213 4276 4273 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06864 8787 6232 4276 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06863 4275 4276 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06862 8787 4271 4274 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06861 4273 4272 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06860 4268 4275 4212 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06859 4211 4276 4268 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06858 8787 5998 4211 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06857 5998 4268 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06856 8787 4268 5998 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06855 2122 3857 2040 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06854 2040 2121 2122 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06853 8787 3261 2040 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06852 3537 3765 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06851 3538 5044 3537 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06850 6103 8764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06849 6104 6316 6103 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06848 5171 5174 5172 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06847 5172 5169 5171 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06846 8787 5170 5172 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06845 8349 7658 7659 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06844 7659 8132 8349 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06843 8787 7657 7659 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06842 2276 3678 2278 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06841 2278 3677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06840 2277 8412 2276 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06839 4000 4529 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06838 4104 4530 4000 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06837 8787 8359 4104 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06836 4105 4104 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06835 6298 6300 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06834 8787 6739 6302 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06833 6181 6299 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06832 6300 6302 6181 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06831 6180 6739 6300 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06830 8787 6296 6180 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06829 7846 8246 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06828 8480 8215 7846 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06827 2433 5562 2432 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06826 2432 6717 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06825 2559 6716 2433 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06824 8787 6878 6575 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06823 6575 6721 6722 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06822 6637 6722 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06821 8274 8362 8275 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06820 8275 8361 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06819 8273 8625 8274 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06818 8369 8623 8273 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06817 2331 5563 2330 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06816 2330 3753 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06815 2548 5470 2331 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06814 6296 6063 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06813 8787 6920 6065 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06812 6064 6062 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06811 6063 6065 6064 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06810 6061 6920 6063 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06809 8787 6060 6061 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06808 5760 6940 5759 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06807 5759 6673 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06806 5758 7184 5760 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06805 5916 8490 5758 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06804 7173 8222 7027 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06803 7027 8246 7173 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06802 8787 8247 7027 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06801 1172 3964 1171 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06800 1171 6717 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06799 2161 5562 1172 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06798 1444 1702 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06797 8787 1702 1445 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06796 1879 1443 1444 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06795 1442 1445 1879 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06794 8787 1447 1442 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06793 1443 1447 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06792 3219 4533 3220 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06791 3220 4027 3301 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06790 8787 3300 3219 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06789 4327 3301 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06788 3500 6286 3499 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06787 3499 3749 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06786 3501 6282 3500 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06785 3498 6716 3501 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06784 6010 6717 6012 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06783 6012 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06782 6011 6026 6010 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06781 6711 7514 6011 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06780 4068 4070 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06779 8787 4075 4072 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06778 3989 4941 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06777 4070 4072 3989 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06776 3988 4075 4070 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06775 8787 7718 3988 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06774 4307 8350 6735 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06773 8787 8350 4306 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06772 4308 4727 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06771 6735 4306 4308 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06770 8787 4305 4307 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06769 3809 6027 3808 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06768 8787 8627 3810 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06767 3808 3810 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06766 3384 3648 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06765 8787 3648 3385 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06764 3825 3382 3384 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06763 3383 3385 3825 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06762 8787 3644 3383 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06761 3382 3644 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06760 7295 7529 7296 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06759 7296 7528 7295 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06758 8787 7947 7296 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06757 7523 7295 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06756 8787 6466 5648 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06755 5648 6072 5649 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06754 5647 5649 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06753 8787 4577 1653 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06752 1653 2764 1802 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06751 2015 1802 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06750 8787 8240 7462 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06749 7462 8030 7583 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06748 8023 7583 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06747 6619 8222 6618 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06746 6618 8483 6771 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06745 8787 8237 6619 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06744 6673 6771 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06743 7245 7251 7244 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06742 7244 7243 7245 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06741 8787 8350 7244 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06740 7411 7478 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06739 7477 7637 7411 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06738 8787 7476 7477 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06737 7475 7477 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06736 1283 1288 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06735 8787 1283 1217 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06734 1217 1290 1288 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06733 1288 1291 1219 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06732 8787 1302 1291 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06731 1290 1291 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06730 8787 1218 1289 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06729 1219 1285 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06728 1281 1290 1283 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06727 1216 1291 1281 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06726 8787 1280 1216 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06725 1280 1281 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06724 8787 1281 1280 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06723 1550 1552 1554 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06722 1554 1553 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06721 1551 1772 1550 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06720 2974 1549 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06719 1549 1548 1551 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06718 3163 3168 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06717 3166 5046 3168 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06716 3168 6111 3167 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06715 3167 5280 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06714 8787 3164 3166 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06713 3166 3165 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06712 3611 3767 3612 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06711 3612 6282 3760 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06710 8787 5562 3611 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06709 7115 3760 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06708 1885 2105 1884 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06707 1884 1882 1885 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06706 8787 1883 1884 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06705 2108 1885 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06704 6724 7118 6577 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06703 6577 7115 6724 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06702 8787 8160 6577 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06701 6817 6724 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06700 8575 8580 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06699 8787 8575 8576 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06698 8576 8582 8580 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06697 8580 8584 8581 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06696 8787 8596 8584 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06695 8582 8584 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06694 8787 8578 8583 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06693 8581 8579 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06692 8573 8582 8575 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06691 8574 8584 8573 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06690 8787 8572 8574 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06689 8572 8573 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06688 8787 8573 8572 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06687 57 59 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06686 8787 57 3 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06685 3 61 59 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06684 59 63 2 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06683 8787 1302 63 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06682 61 63 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06681 8787 4 62 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06680 2 56 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06679 55 61 57 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06678 1 63 55 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06677 8787 274 1 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06676 274 55 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06675 8787 55 274 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06674 2051 2139 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06673 2263 3275 2051 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06672 4716 7643 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06671 4714 4715 4716 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06670 2050 3445 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06669 2138 2137 2050 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06668 3047 3502 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06667 3154 4139 3047 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06666 5237 5239 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06665 8787 6312 5240 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06664 5238 5440 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06663 5239 5240 5238 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06662 5236 6312 5239 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06661 8787 5365 5236 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06660 8333 8334 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06659 8787 8333 8259 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06658 8259 8339 8334 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06657 8334 8338 8261 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06656 8787 8596 8338 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06655 8339 8338 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06654 8787 8260 8336 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06653 8261 8309 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06652 8330 8339 8333 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06651 8258 8338 8330 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06650 8787 8329 8258 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06649 8329 8330 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06648 8787 8330 8329 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06647 8787 6955 6545 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06646 6545 6668 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06645 6543 6544 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06644 6545 7752 6544 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06643 6544 6770 6545 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06642 4395 5415 4396 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06641 4396 4499 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06640 4498 6283 4395 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06639 4584 4587 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06638 8787 8764 4588 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06637 4366 6125 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06636 4587 4588 4366 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06635 4365 8764 4587 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06634 8787 4583 4365 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06633 8787 2159 1252 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06632 1252 4027 1361 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06631 1539 1361 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06630 1318 1320 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06629 8787 1862 1322 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06628 1233 3254 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06627 1320 1322 1233 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06626 1232 1862 1320 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06625 8787 3673 1232 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06624 2690 3956 2689 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06623 2689 6043 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06622 2688 6284 2690 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06621 2927 7228 2688 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06620 8787 7106 6997 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06619 6997 7099 7100 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06618 7522 7100 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06617 5641 5643 5642 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06616 5642 5644 5641 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06615 8787 6062 5642 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06614 3937 6718 3938 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06613 3938 4135 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06612 3935 3964 3937 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06611 3936 5471 3935 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06610 6137 8490 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06609 6136 8240 6137 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06608 7917 8324 7779 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06607 7779 8321 7917 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06606 8787 8627 7779 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06605 7852 7917 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06604 8787 6878 6461 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06603 6461 6462 6463 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06602 6727 6463 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06601 5274 6115 5273 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06600 5273 5505 5274 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06599 8787 5272 5273 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06598 8787 6878 6425 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06597 6425 6426 6427 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06596 6699 6427 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06595 877 1553 876 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06594 876 4750 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06593 875 4529 877 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06592 1019 1552 875 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06591 1323 1114 1111 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06590 1111 1113 1323 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06589 8787 2260 1111 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06588 844 931 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06587 927 1128 844 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06586 843 1129 927 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06585 8787 925 843 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06584 2248 927 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06583 8787 1123 842 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06582 842 926 927 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06581 8787 4744 4702 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06580 4702 5160 4701 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06579 4700 4701 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06578 3630 5471 3631 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06577 3631 5562 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06576 3629 4300 3630 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06575 4157 4139 3629 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06574 7059 7049 6804 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06573 8787 8065 6805 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06572 6804 6805 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06571 3515 5013 3514 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06570 3514 6286 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06569 3513 6026 3515 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06568 3512 3511 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06567 3511 3510 3513 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06566 1264 6040 1263 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06565 1263 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06564 1262 4577 1264 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06563 1566 1371 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06562 1371 1276 1262 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06561 7337 7342 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06560 8787 7337 7338 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06559 7338 7344 7342 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06558 7342 7346 7341 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06557 8787 8728 7346 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06556 7344 7346 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06555 8787 7339 7343 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06554 7341 7340 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06553 7335 7344 7337 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06552 7336 7346 7335 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06551 8787 7345 7336 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06550 7345 7335 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06549 8787 7335 7345 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06548 2090 2176 2091 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06547 2091 2571 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06546 2089 2350 2090 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06545 2173 2175 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06544 2175 2088 2089 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06543 8787 2373 2372 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06542 2373 2592 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06541 2372 3009 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06540 8787 3049 2979 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06539 2979 2968 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06538 8787 3307 2979 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06537 2452 4143 2453 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06536 2453 2582 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06535 2451 2587 2452 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06534 2591 2583 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06533 2583 2464 2451 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06532 6897 7127 6896 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06531 6896 7126 6897 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06530 8787 7723 6896 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06529 7112 6897 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06528 5540 5542 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06527 8787 5540 5541 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06526 5541 5577 5542 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06525 5542 5578 5574 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06524 8787 6232 5578 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06523 5577 5578 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06522 8787 5575 5576 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06521 5574 5573 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06520 5572 5577 5540 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06519 5539 5578 5572 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06518 8787 6271 5539 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06517 6271 5572 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06516 8787 5572 6271 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06515 6278 8175 6167 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06514 6167 6276 6278 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06513 8787 6462 6167 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06512 6275 6278 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06511 2742 6284 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06510 2743 2741 2742 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06509 8787 3531 2739 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06508 2739 3297 2743 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06507 8787 3133 2740 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06506 2740 3767 2743 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06505 4505 4502 4400 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06504 4400 6860 4505 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06503 8787 4503 4400 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06502 4520 4505 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06501 2256 3678 2254 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06500 2254 3677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06499 2255 7326 2256 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06498 3214 5465 3215 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06497 3215 3490 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06496 3300 4300 3214 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06495 2997 2996 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06494 2996 2893 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06493 8787 3171 2996 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06492 2785 2784 2786 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06491 2786 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06490 2998 4577 2785 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06489 6542 6644 6540 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06488 6540 8483 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06487 6541 8237 6542 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06486 8787 4320 4293 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06485 4293 4292 4294 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06484 4518 4294 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06483 1619 2508 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06482 1733 3269 1619 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06481 8787 1956 1733 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06480 1916 1733 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06479 6968 8488 6967 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06478 6967 7592 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06477 6965 6964 6968 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06476 6966 8240 6965 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06475 4216 4305 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06474 4697 8350 4216 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06473 6572 6717 6573 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06472 6573 6718 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06471 6571 6716 6572 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06470 6879 8372 6571 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06469 75 77 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06468 8787 983 79 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06467 10 3843 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06466 77 79 10 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06465 9 983 77 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06464 8787 276 9 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06463 338 340 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06462 8787 983 342 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06461 341 2718 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06460 340 342 341 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06459 339 983 340 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06458 8787 992 339 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06457 8787 817 818 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06456 1180 818 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06455 8787 818 1180 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06454 8787 818 1180 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06453 1180 818 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06452 8787 1180 1181 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06451 6037 1181 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06450 8787 1181 6037 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06449 8787 1181 6037 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06448 6037 1181 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06447 8787 1180 1025 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06446 6285 1025 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06445 8787 1025 6285 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06444 8787 1025 6285 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06443 6285 1025 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06442 2013 3898 2014 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06441 2014 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06440 2012 6282 2013 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06439 2180 6021 2012 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06438 8787 8785 8786 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06437 8784 8786 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06436 8787 8786 8784 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06435 8787 8786 8784 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06434 8784 8786 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06433 8787 8784 8489 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06432 8488 8489 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06431 8787 8489 8488 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06430 8787 8489 8488 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06429 8488 8489 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06428 8787 8784 8491 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06427 8490 8491 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06426 8787 8491 8490 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06425 8787 8491 8490 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06424 8490 8491 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06423 8787 5196 5190 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06422 5190 5841 5191 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06421 5189 5191 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06420 8787 3180 3182 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06419 3182 3541 3183 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06418 3181 3183 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06417 8787 8455 7753 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06416 7753 8220 7754 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06415 7752 7754 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06414 8787 4826 3971 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06413 3971 3969 3970 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06412 3968 3970 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06411 6367 6664 6202 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06410 6202 6370 6367 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06409 8787 7315 6202 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06408 6365 6367 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06407 878 4750 879 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06406 879 1021 1022 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06405 8787 2161 878 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06404 1020 1022 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06403 8100 8098 8101 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06402 8101 8097 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06401 8099 8235 8100 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06400 8778 8230 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06399 8230 8096 8099 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06398 8199 8690 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06397 4233 4235 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06396 8787 4233 4234 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06395 4234 4371 4235 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06394 4235 4373 4370 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06393 8787 6361 4373 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06392 4371 4373 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06391 8787 4368 4372 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06390 4370 4369 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06389 4367 4371 4233 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06388 4232 4373 4367 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06387 8787 4583 4232 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06386 4583 4367 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06385 8787 4367 4583 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06384 4380 6934 4471 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06383 8787 6934 4472 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06382 4381 4469 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06381 4471 4472 4381 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06380 8787 4473 4380 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06379 1929 2511 1930 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06378 1930 1928 1929 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06377 8787 2936 1930 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06376 1926 1929 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06375 1112 3110 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06374 1915 1323 1112 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06373 3670 3676 3570 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06372 3570 3672 3670 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06371 8787 3673 3570 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06370 1998 1997 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06369 8787 2344 1998 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06368 5033 4350 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06367 4580 4358 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06366 8191 8703 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06365 5685 6115 5686 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06364 5686 5683 5685 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06363 8787 5684 5686 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06362 8639 8632 8633 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06361 8633 8630 8639 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06360 8787 8631 8633 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06359 1009 2986 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06358 7847 8778 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06357 7912 8030 7847 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06356 6165 6272 6164 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06355 6164 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06354 6447 8648 6165 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06353 7097 7118 6996 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06352 6996 7115 7097 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06351 8787 7660 6996 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06350 7096 7097 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06349 6547 6549 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06348 6548 7767 6547 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06347 8301 8764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06346 8473 8472 8301 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06345 5651 5655 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06344 8787 5656 5659 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06343 5657 5660 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06342 5655 5659 5657 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06341 5654 5656 5655 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06340 8787 6060 5654 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06339 601 608 455 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06338 455 599 601 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06337 8787 793 455 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06336 783 601 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06335 5558 8237 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06334 5557 7315 5558 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06333 1251 4532 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06332 1358 1552 1251 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06331 8693 8694 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06330 8787 8693 8695 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06329 8695 8701 8694 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06328 8694 8702 8700 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06327 8787 8728 8702 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06326 8701 8702 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06325 8787 8697 8699 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06324 8700 8698 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06323 8692 8701 8693 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06322 8691 8702 8692 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06321 8787 8690 8691 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06320 8690 8692 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06319 8787 8692 8690 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06318 6570 7315 6569 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06317 6569 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06316 6635 7660 6570 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06315 8787 6878 6880 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06314 6880 6879 6881 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06313 6882 6881 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06312 2447 2579 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06311 2782 2578 2447 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06310 3891 4027 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06309 7118 4533 3891 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06308 5864 5867 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06307 8787 6307 5869 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06306 5663 8412 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06305 5867 5869 5663 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06304 5661 6307 5867 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06303 8787 5865 5661 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06302 8787 7304 7302 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06301 7302 7300 7301 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06300 7532 7301 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06299 6347 6100 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06298 8787 8764 6101 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06297 6099 6660 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06296 6100 6101 6099 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06295 6098 8764 6100 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06294 8787 6339 6098 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06293 8763 8766 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06292 8787 8764 8767 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06291 8765 8778 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06290 8766 8767 8765 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06289 8762 8764 8766 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06288 8787 8761 8762 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06287 8787 6878 6423 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06286 6423 6422 6424 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06285 6844 6424 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06284 8098 7979 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06283 8787 8430 7980 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06282 7805 8168 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06281 7979 7980 7805 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06280 7804 8430 7979 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06279 8787 8399 7804 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06278 5818 7273 5717 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06277 5717 6007 5818 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06276 8787 6290 5717 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06275 5116 5466 5117 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06274 5117 5790 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06273 5587 5415 5116 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06272 5743 5891 5744 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06271 5744 6320 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06270 5742 7349 5743 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06269 5890 8478 5742 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06268 5031 5043 4907 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06267 4907 5243 5031 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06266 8787 5041 4907 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06265 1158 6021 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06264 3903 1157 1158 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06263 8787 2784 1156 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06262 1156 4577 3903 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06261 8787 3531 1155 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06260 1155 1154 3903 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06259 5234 6284 5235 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06258 5235 5471 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06257 5233 5470 5234 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06256 5469 8350 5233 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06255 5973 5974 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06254 8787 5974 5975 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06253 6293 5971 5973 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06252 5972 5975 6293 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06251 8787 6433 5972 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06250 5971 6433 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06249 2352 5562 2353 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06248 2353 3531 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06247 2351 5471 2352 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06246 2350 3333 2351 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06245 7688 7689 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06244 7689 8359 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06243 8787 7880 7689 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06242 7689 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06241 8787 7877 7689 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06240 8049 7637 7638 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06239 7638 7639 8049 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06238 8787 7636 7638 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06237 2481 2251 2034 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06236 2034 2252 2481 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06235 8787 2260 2034 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06234 8787 6282 872 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06233 872 3898 1018 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06232 1154 1018 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06231 4282 4279 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06230 8787 4279 4277 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06229 4281 4280 4282 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06228 4278 4277 4281 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06227 8787 4498 4278 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06226 4280 4498 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06225 8248 8483 8249 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06224 8249 8246 8248 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06223 8787 8247 8249 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06222 8787 5280 2846 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06221 2846 6530 3002 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06220 3001 3002 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06219 4854 5137 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06218 8787 5137 4948 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06217 4947 4945 4854 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06216 4853 4948 4947 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06215 8787 6872 4853 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06214 4945 6872 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06213 7543 7307 7309 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06212 7309 7308 7543 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06211 8787 8412 7309 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06210 4116 4118 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06209 8787 4116 4004 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06208 4004 4115 4118 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06207 4118 4122 4005 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06206 8787 4121 4122 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06205 4115 4122 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06204 8787 4032 4120 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06203 4005 4043 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06202 4114 4115 4116 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06201 4003 4122 4114 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06200 8787 8430 4003 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06199 8430 4114 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06198 8787 4114 8430 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06197 2234 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06196 2644 2648 2234 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06195 2233 2482 2644 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06194 8787 3655 2233 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06193 2233 2639 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06192 3947 4109 3948 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06191 3948 6037 3949 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06190 8787 6284 3947 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06189 3946 3949 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06188 6830 8235 6831 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06187 6831 8020 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06186 6829 7394 6830 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06185 6954 6953 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06184 6953 6828 6829 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06183 5350 6284 5351 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06182 5351 5471 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06181 5349 5470 5350 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06180 5891 5472 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06179 5472 5348 5349 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06178 1393 1394 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06177 8787 1393 1272 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06176 1272 1399 1394 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06175 1394 1400 1274 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06174 8787 2028 1400 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06173 1399 1400 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06172 8787 1273 1398 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06171 1274 1396 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06170 1391 1399 1393 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06169 1271 1400 1391 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06168 8787 1390 1271 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06167 1390 1391 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06166 8787 1391 1390 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06165 1917 1476 1478 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06164 1478 3273 1917 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06163 8787 1477 1478 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06162 8270 8358 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06161 8632 8627 8270 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06160 1984 4529 1996 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06159 1996 2890 1984 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06158 8787 1983 1984 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06157 1984 3716 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06156 4882 5563 4881 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06155 4881 5562 4998 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06154 8787 6716 4882 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06153 5446 4998 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06152 6533 6644 6532 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06151 6532 8483 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06150 6531 7394 6533 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06149 6530 6529 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06148 6529 6528 6531 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06147 1187 6037 1188 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06146 1188 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06145 1185 3898 1187 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06144 1372 1186 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06143 1186 1184 1185 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06142 5637 6290 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_06141 8787 6271 5637 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_06140 5637 6022 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_06139 8787 6027 5637 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_06138 2291 2297 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06137 8787 2291 2292 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06136 2292 2299 2297 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06135 2297 2300 2296 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06134 8787 3705 2300 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06133 2299 2300 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06132 8787 2294 2298 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06131 2296 2295 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06130 2290 2299 2291 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06129 2289 2300 2290 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06128 8787 5188 2289 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06127 5188 2290 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06126 8787 2290 5188 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06125 5843 5263 4752 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06124 4752 4750 5843 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06123 8787 4999 4752 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06122 4954 5143 4856 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06121 4856 6246 4954 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06120 8787 4951 4856 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06119 4952 4954 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06118 4341 4338 4340 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06117 4340 4339 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06116 4562 5870 4341 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06115 5399 5400 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06114 8787 5399 5304 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06113 5304 5398 5400 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06112 5400 5405 5305 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06111 8787 6232 5405 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06110 5398 5405 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06109 8787 5343 5404 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06108 5305 5360 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06107 5396 5398 5399 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06106 5303 5405 5396 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06105 8787 6251 5303 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06104 6251 5396 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06103 8787 5396 6251 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06102 1547 1546 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06101 2748 4027 1547 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06100 6126 6128 6127 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06099 6127 7177 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06098 6125 6377 6126 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06097 8787 2937 1622 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06096 1622 2277 1742 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06095 1741 1742 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06094 2053 5013 2054 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06093 2054 3898 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06092 2151 6284 2053 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06091 2442 3295 2441 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06090 2441 2983 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06089 2571 3964 2442 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06088 1640 4792 1639 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06087 1639 1768 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06086 1976 1772 1640 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06085 2324 6307 2326 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06084 2326 2328 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06083 2325 2760 2324 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06082 8787 5432 5177 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06081 5177 5176 5178 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06080 5426 5178 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06079 8787 6878 6166 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06078 6166 6287 6274 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06077 6273 6274 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06076 2402 3678 2401 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06075 2401 3677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06074 2508 8417 2402 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06073 3627 3960 3628 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06072 3628 4111 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06071 3626 6282 3627 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06070 4154 3767 3626 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06069 6445 6717 6444 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06068 6444 6718 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06067 6443 6716 6445 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06066 6721 8648 6443 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06065 6176 6286 6175 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06064 6175 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06063 6174 6284 6176 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06062 6726 6283 6174 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06061 3811 3639 3381 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06060 3381 4469 3811 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06059 8787 8627 3381 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06058 1989 4530 1988 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06057 1988 2890 1989 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06056 8787 1987 1989 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06055 1989 3717 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06054 8072 8349 8073 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06053 8073 8348 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06052 8071 8346 8072 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06051 8623 8119 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06050 8119 8070 8071 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06049 8787 168 158 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06048 1760 158 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06047 8787 158 1760 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06046 8787 158 1760 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06045 1760 158 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06044 8787 1760 1761 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06043 6043 1761 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06042 8787 1761 6043 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06041 8787 1761 6043 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06040 6043 1761 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06039 8787 1760 1357 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06038 6286 1357 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06037 8787 1357 6286 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06036 8787 1357 6286 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06035 6286 1357 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06034 8787 1760 1528 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06033 6029 1528 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06032 8787 1528 6029 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06031 8787 1528 6029 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06030 6029 1528 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06029 8787 1760 157 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06028 6718 157 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06027 8787 157 6718 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06026 8787 157 6718 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06025 6718 157 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06024 3480 6095 3481 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06023 3481 4327 3480 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06022 8787 3478 3481 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06021 3479 3480 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06020 6847 7049 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06019 6848 7643 6847 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06018 8787 6846 6848 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06017 7252 6848 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06016 6260 7311 6157 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06015 6157 6276 6260 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06014 8787 6711 6157 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06013 6259 6260 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06012 8787 4300 1652 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06011 1652 2764 1801 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06010 2016 1801 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06009 3588 4103 3589 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06008 3589 3721 3719 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06007 8787 3884 3588 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06006 3718 3719 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06005 2430 6718 2429 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06004 2429 6285 2547 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06003 8787 3136 2430 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06002 2749 2547 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06001 740 737 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06000 8787 740 677 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05999 677 746 737 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05998 737 745 743 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05997 8787 1302 745 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05996 746 745 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05995 8787 741 744 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05994 743 742 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05993 736 746 740 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05992 676 745 736 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05991 8787 1105 676 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05990 1105 736 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05989 8787 736 1105 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05988 7834 8782 7835 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05987 7835 8209 8015 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05986 8787 8780 7834 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05985 8478 8015 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05984 7547 7716 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05983 1369 1390 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05982 3136 1567 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05981 691 5192 692 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05980 692 4111 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05979 690 5563 691 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05978 1030 820 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05977 820 821 690 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05976 5988 6250 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05975 5363 8433 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05974 6902 7127 6901 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05973 6901 7126 6902 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05972 8787 8412 6901 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05971 6900 6902 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05970 7231 7232 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05969 8787 7231 7233 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05968 7233 7239 7232 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05967 7232 7238 7236 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05966 8787 8596 7238 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05965 7239 7238 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05964 8787 7234 7237 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05963 7236 7235 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05962 7230 7239 7231 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05961 7229 7238 7230 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05960 8787 7228 7229 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05959 7228 7230 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05958 8787 7230 7228 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05957 8362 8359 7796 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05956 7796 8132 8362 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05955 8787 8131 7796 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05954 1139 5214 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05953 1138 1140 1139 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05952 2551 2554 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05951 2554 2553 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05950 8787 3150 2554 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05949 850 5412 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05948 943 1100 850 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05947 2759 2784 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05946 2760 6716 2759 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05945 5459 5462 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05944 8787 5461 5464 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05943 5322 5460 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05942 5462 5464 5322 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05941 5321 5461 5462 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05940 8787 5872 5321 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05939 8052 8054 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05938 8787 8052 8053 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05937 8053 8056 8054 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05936 8054 8106 8105 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05935 8787 8596 8106 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05934 8056 8106 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05933 8787 8107 8108 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05932 8105 8104 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05931 8102 8056 8052 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05930 8051 8106 8102 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05929 8787 8103 8051 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05928 8103 8102 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05927 8787 8102 8103 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05926 6473 6068 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05925 8787 6075 6069 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05924 6067 6466 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05923 6068 6069 6067 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05922 6066 6075 6068 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05921 8787 6303 6066 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05920 8787 7315 7316 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05919 7316 8215 7317 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05918 7528 7317 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05917 8787 7066 6839 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05916 6839 7065 6840 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05915 7246 6840 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05914 8787 6763 6706 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05913 7684 6706 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05912 8787 6706 7684 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05911 8787 6706 7684 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05910 7684 6706 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05909 8787 6763 6762 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05908 7765 6762 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05907 8787 6762 7765 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05906 8787 6762 7765 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05905 7765 6762 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05904 8787 4311 4312 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05903 6763 4312 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05902 8787 4312 6763 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05901 8787 4312 6763 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05900 6763 4312 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05899 5133 6022 5132 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05898 5132 5139 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05897 5130 5415 5133 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05896 2850 3106 2851 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05895 2851 3668 2919 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05894 8787 3657 2850 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05893 3247 2919 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05892 4347 5471 4348 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05891 4348 5465 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05890 4345 6716 4347 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05889 4346 8461 4345 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05888 2457 2587 2458 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05887 2458 3180 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05886 2803 2783 2457 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05885 8787 4753 4755 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05884 4753 4751 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05883 4755 4754 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05882 8787 5609 5608 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05881 5608 5993 5607 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05880 5606 5607 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05879 6358 6115 6110 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05878 6110 6364 6358 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05877 8787 6109 6110 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05876 3111 6288 3112 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05875 3112 5408 3111 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05874 8787 5631 3112 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05873 3110 3111 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05872 8787 2566 466 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05871 466 1390 619 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05870 817 619 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05869 6747 6748 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05868 8787 6747 6587 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05867 6587 6746 6748 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05866 6748 6751 6588 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05865 8787 8728 6751 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05864 6746 6751 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05863 8787 6616 6749 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05862 6588 6652 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05861 6744 6746 6747 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05860 6586 6751 6744 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05859 8787 6920 6586 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05858 6920 6744 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05857 8787 6744 6920 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05856 3122 3125 3123 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05855 3123 3121 3124 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05854 8787 3120 3122 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05853 3280 3124 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05852 3264 3271 3194 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05851 3194 3262 3264 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05850 8787 3261 3194 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05849 3392 3264 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05848 2405 2940 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05847 2513 3479 2405 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05846 8787 2942 2513 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05845 2511 2513 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05844 8024 8098 7824 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05843 7824 8246 8024 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05842 8787 8247 7824 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05841 7908 8024 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05840 6113 6644 6112 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05839 6112 8483 6114 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05838 8787 8237 6113 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05837 6111 6114 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05836 4554 4759 4427 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05835 4427 7315 4554 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05834 8787 4553 4427 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05833 5568 5569 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05832 8787 5568 5570 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05831 5570 5693 5569 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05830 5569 5692 5690 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05829 8787 6361 5692 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05828 5693 5692 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05827 8787 5688 5691 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05826 5690 5689 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05825 5687 5693 5568 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05824 5567 5692 5687 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05823 8787 5907 5567 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05822 5907 5687 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05821 8787 5687 5907 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05820 5773 6674 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05819 5922 6378 5773 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05818 1583 5046 1582 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05817 1582 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05816 1581 3753 1583 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05815 1791 1580 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05814 1580 1579 1581 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05813 8787 7096 7091 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05812 7091 7087 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05811 8787 7088 7091 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05810 2259 2949 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05809 3414 5676 2259 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05808 2938 2273 2275 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05807 2275 2274 2938 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05806 8787 2723 2275 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05805 4460 4462 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05804 8787 4460 4378 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05803 4378 4466 4462 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05802 4462 4467 4377 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05801 8787 6232 4467 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05800 4466 4467 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05799 8787 4379 4465 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05798 4377 4452 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05797 4459 4466 4460 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05796 4376 4467 4459 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05795 8787 6022 4376 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05794 6022 4459 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05793 8787 4459 6022 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05792 7831 7957 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05791 7874 8369 7831 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05790 3231 3519 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05789 3526 3318 3231 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05788 682 2734 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05787 983 1129 682 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05786 8787 2927 2819 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05785 2819 2933 2928 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05784 2926 2928 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05783 8787 3414 3418 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05782 3420 3482 3413 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05781 3417 5580 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_05780 3413 3412 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05779 3418 3415 3416 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05778 3416 5580 3420 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05777 3420 3417 3419 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05776 3411 3420 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05775 8787 3414 3412 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_05774 3419 3671 3418 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05773 8787 3414 2654 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05772 2657 3660 2651 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05771 2655 3066 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_05770 2651 2652 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05769 2654 2659 2653 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05768 2653 3066 2657 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05767 2657 2655 2656 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05766 3646 2657 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05765 8787 3414 2652 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_05764 2656 3665 2654 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05763 3572 3678 3573 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05762 3573 3677 3679 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05761 8787 7142 3572 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05760 3676 3679 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05759 1116 1113 1110 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05758 1110 1114 1116 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05757 8787 2723 1110 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05756 3966 5046 3967 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05755 3967 4111 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05754 3965 6282 3966 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05753 3978 3964 3965 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05752 7887 8383 7833 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05751 8787 8627 7964 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05750 7833 7964 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05749 6522 8490 6523 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05748 6523 6954 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05747 6766 8240 6522 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05746 2761 2890 2762 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05745 2762 2760 2761 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05744 8787 2763 2762 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05743 2847 2761 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05742 8787 632 630 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05741 831 630 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05740 8787 630 831 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05739 8787 630 831 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05738 831 630 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05737 8787 831 830 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05736 6040 830 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05735 8787 830 6040 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05734 8787 830 6040 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05733 6040 830 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05732 8787 831 627 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05731 6717 627 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05730 8787 627 6717 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05729 8787 627 6717 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05728 6717 627 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05727 8787 831 832 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05726 6282 832 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05725 8787 832 6282 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05724 8787 832 6282 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05723 6282 832 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05722 3325 3311 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05721 8787 3307 3311 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05720 3311 3759 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05719 8787 3310 3311 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05718 2076 2161 2077 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05717 2077 2160 2162 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05716 8787 6077 2076 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05715 4127 2162 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05714 7690 7502 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05713 7502 7933 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05712 8787 7880 7502 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05711 7502 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05710 8787 7499 7502 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05709 8787 836 837 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05708 835 837 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05707 8787 837 835 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05706 8787 837 835 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05705 835 837 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05704 8787 835 833 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05703 3960 833 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05702 8787 833 3960 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05701 8787 833 3960 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05700 3960 833 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05699 8787 835 834 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05698 5046 834 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05697 8787 834 5046 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05696 8787 834 5046 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05695 5046 834 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05694 8787 2176 2092 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05693 2092 2571 2177 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05692 2354 2177 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05691 8787 2578 2446 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05690 2446 2579 2577 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05689 2999 2577 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05688 7405 8246 7407 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05687 7407 8236 7406 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05686 8787 8237 7405 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05685 7404 7406 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05684 8631 8634 8628 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05683 8787 8627 8629 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05682 8628 8629 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05681 1196 3531 1197 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05680 1197 2764 1198 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05679 8787 4139 1196 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05678 1381 1198 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05677 8720 8722 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05676 8787 8720 8721 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05675 8721 8729 8722 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05674 8722 8730 8726 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05673 8787 8728 8730 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05672 8729 8730 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05671 8787 8724 8727 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05670 8726 8725 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05669 8719 8729 8720 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05668 8718 8730 8719 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05667 8787 8717 8718 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05666 8717 8719 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05665 8787 8719 8717 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05664 6247 6000 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05663 5613 5612 5614 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05662 5614 6246 5613 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05661 8787 7495 5614 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05660 5611 5613 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05659 8787 6072 5246 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05658 5246 6758 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05657 8787 8717 5246 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05656 4802 4805 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05655 8787 4802 4806 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05654 4806 4810 4805 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05653 4805 4809 4804 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05652 8787 6361 4809 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05651 4810 4809 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05650 8787 4807 4808 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05649 4804 4803 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05648 4801 4810 4802 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05647 4800 4809 4801 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05646 8787 5036 4800 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05645 5036 4801 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05644 8787 4801 5036 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05643 1606 4577 1607 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05642 1607 3898 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05641 1604 5013 1606 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05640 1602 1605 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05639 1605 1603 1604 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05638 8359 8634 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05637 7277 7947 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05636 5436 5188 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05635 683 4027 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05634 792 2159 683 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05633 3880 3897 3879 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05632 3879 7115 3880 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05631 8787 6022 3879 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05630 4557 4751 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05629 4434 4789 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05628 4778 4562 4434 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05627 3824 3831 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05626 3829 3827 3831 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05625 3831 3828 3830 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05624 3830 3832 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05623 8787 3825 3829 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05622 3829 3826 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05621 1117 4700 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05620 1118 1116 1117 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05619 3237 6530 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05618 3326 5280 3237 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05617 8706 8710 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05616 8787 8706 8709 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05615 8709 8714 8710 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05614 8710 8715 8708 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05613 8787 8728 8715 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05612 8714 8715 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05611 8787 8712 8713 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05610 8708 8707 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05609 8705 8714 8706 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05608 8704 8715 8705 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05607 8787 8703 8704 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05606 8703 8705 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05605 8787 8705 8703 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05604 3477 6282 3476 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05603 3476 6286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05602 3475 6716 3477 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05601 3478 3750 3475 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05600 3207 4750 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05599 3288 4529 3207 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05598 5187 5189 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05597 5341 5186 5187 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05596 6515 6517 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05595 8787 8764 6519 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05594 6518 6936 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05593 6517 6519 6518 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05592 6516 8764 6517 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05591 8787 6514 6516 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05590 2859 3083 2860 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05589 2860 3479 2941 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05588 8787 2940 2859 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05587 3657 2941 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05586 8787 6767 6664 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05585 6767 7173 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05584 6664 7749 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05583 5677 5680 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05582 8787 7347 5681 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05581 5679 5895 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05580 5680 5681 5679 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05579 5678 7347 5680 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05578 8787 5676 5678 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05577 8787 7543 7430 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05576 7430 7542 7544 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05575 7932 7544 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05574 2964 2965 2837 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05573 2837 2966 2964 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05572 8787 8731 2837 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05571 3488 6282 3489 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05570 3489 3898 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05569 4750 4577 3488 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05568 3315 1977 1979 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05567 1979 1978 3315 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05566 8787 7535 1979 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05565 1783 1376 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05564 1376 1374 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05563 8787 1373 1376 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05562 1995 1032 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05561 1032 1031 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05560 8787 1030 1032 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05559 6927 6929 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05558 8787 8764 6930 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05557 6928 7573 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05556 6929 6930 6928 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05555 6926 8764 6929 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05554 8787 6925 6926 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05553 2046 2272 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05552 8787 2272 2135 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05551 2517 2132 2046 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05550 2045 2135 2517 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05549 8787 2133 2045 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05548 2132 2133 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05547 7255 7251 7254 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05546 7254 7481 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05545 7256 7252 7255 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05544 8326 7250 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05543 7250 7253 7256 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05542 8787 1992 1994 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05541 1994 3318 1993 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05540 2000 1993 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05539 8787 6718 3131 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05538 3131 6285 3130 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05537 3294 3130 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05536 117 119 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05535 8787 117 25 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05534 25 121 119 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05533 119 123 24 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05532 8787 1516 123 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05531 121 123 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05530 8787 26 122 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05529 24 116 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05528 115 121 117 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05527 23 123 115 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05526 8787 554 23 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05525 554 115 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05524 8787 115 554 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05523 4318 4747 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05522 8787 4751 4318 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05521 2097 3335 2098 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05520 2098 2981 2186 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05519 8787 2185 2097 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05518 2374 2186 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05517 7836 8450 7837 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05516 7837 8781 8016 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05515 8787 8237 7836 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05514 8030 8016 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05513 5821 6006 5718 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05512 5718 6246 5821 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05511 8787 6428 5718 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05510 5822 5821 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05509 795 604 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05508 472 602 604 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05507 604 4300 473 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05506 473 3295 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05505 8787 1009 472 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05504 472 5192 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05503 4729 4731 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05502 8787 4729 4733 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05501 4733 4735 4731 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05500 4731 4737 4732 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05499 8787 5835 4737 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05498 4735 4737 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05497 8787 4734 4736 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05496 4732 4730 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05495 4728 4735 4729 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05494 4726 4737 4728 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05493 8787 4727 4726 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05492 4727 4728 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05491 8787 4728 4727 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05490 7838 8222 7839 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05489 7839 8223 8017 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05488 8787 8780 7838 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05487 8240 8017 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05486 7380 8023 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05485 7381 7379 7380 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05484 8787 7579 7377 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05483 7377 7400 7381 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05482 8787 7593 7378 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05481 7378 7756 7381 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05480 265 269 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05479 8787 265 268 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05478 268 271 269 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05477 269 273 267 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05476 8787 1302 273 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05475 271 273 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05474 8787 270 272 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05473 267 266 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05472 264 271 265 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05471 263 273 264 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05470 8787 720 263 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05469 720 264 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05468 8787 264 720 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05467 8787 7092 7279 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05466 7279 7093 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05465 8787 7102 7279 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05464 3731 3733 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05463 8787 3731 3596 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05462 3596 3736 3733 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05461 3733 3738 3595 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05460 8787 4121 3738 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05459 3736 3738 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05458 8787 3597 3737 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05457 3595 3636 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05456 3730 3736 3731 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05455 3594 3738 3730 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05454 8787 3750 3594 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05453 3750 3730 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05452 8787 3730 3750 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05451 7184 8098 7036 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05450 7036 8246 7184 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05449 8787 8247 7036 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05448 6995 7091 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05447 8617 7275 6995 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05446 4886 4999 4887 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05445 4887 6307 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05444 5216 6077 4886 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05443 8787 4533 2063 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05442 2063 2328 2156 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05441 2155 2156 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05440 390 2974 389 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05439 389 805 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05438 388 4350 390 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05437 2836 3964 2835 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05436 2835 3956 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05435 2960 2961 2836 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05434 8787 5676 2400 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05433 2400 2949 2507 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05432 3261 2507 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05431 462 2974 463 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05430 463 805 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05429 616 5033 462 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05428 47 391 48 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05427 48 2976 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05426 613 807 47 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05425 8787 5231 4771 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05424 4771 5011 4772 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05423 5215 4772 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05422 4303 6029 4304 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05421 4304 6037 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05420 4301 4300 4303 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05419 4302 5440 4301 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05418 1869 4750 1868 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05417 1868 4027 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05416 1867 4529 1869 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05415 2153 1970 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05414 1970 1971 1867 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05413 8787 1016 40 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05412 40 1015 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05411 360 162 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05410 40 369 162 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05409 162 7536 40 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05408 8787 6008 5719 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05407 5719 5822 5823 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05406 5824 5823 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05405 7291 7307 7292 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05404 7292 7308 7291 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05403 8787 7723 7292 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05402 2642 2644 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05401 8787 2644 2643 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05400 2904 2640 2642 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05399 2641 2643 2904 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05398 8787 2639 2641 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05397 2640 2639 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05396 934 935 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05395 8787 934 846 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05394 846 941 935 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05393 935 940 848 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05392 8787 1302 940 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05391 941 940 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05390 8787 847 938 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05389 848 906 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05388 933 941 934 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05387 845 940 933 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05386 8787 931 845 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05385 931 933 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05384 8787 933 931 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05383 4442 4577 4443 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05382 4443 6718 4578 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05381 8787 5563 4442 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05380 5043 4578 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05379 408 3490 410 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05378 410 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05377 409 5465 408 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05376 498 407 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05375 407 406 409 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05374 6988 7472 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05373 7069 7643 6988 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05372 8787 7068 7069 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05371 7481 7069 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05370 913 914 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05369 8787 913 839 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05368 839 918 914 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05367 914 919 841 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05366 8787 1302 919 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05365 918 919 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05364 8787 840 916 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05363 841 905 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05362 911 918 913 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05361 838 919 911 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05360 8787 1092 838 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05359 1092 911 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05358 8787 911 1092 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05357 3999 4529 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05356 4102 4530 3999 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05355 8787 8128 4102 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05354 4103 4102 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05353 7879 8586 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05352 7933 8110 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05351 6095 5220 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05350 8787 5790 4132 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05349 4132 8731 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05348 8787 5036 4132 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05347 4220 4564 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05346 4339 4342 4220 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05345 3394 3824 3393 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05344 3393 3392 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05343 3650 3396 3394 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05342 3872 2504 2399 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05341 2399 2505 3872 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05340 8787 2723 2399 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05339 4713 8103 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05338 4712 4710 4713 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05337 8787 5843 4709 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05336 4709 5440 4712 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05335 8787 4715 4711 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05334 4711 5844 4712 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05333 2145 6324 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05332 5817 8572 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05331 5609 7880 5610 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05330 5610 6007 5609 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05329 8787 6022 5610 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05328 4718 4719 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05327 4719 4717 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05326 8787 5166 4719 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05325 6685 6682 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05324 8787 6685 6558 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05323 6558 6684 6682 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05322 6682 6687 6557 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05321 8787 8596 6687 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05320 6684 6687 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05319 8787 6607 6686 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05318 6557 6621 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05317 6681 6684 6685 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05316 6556 6687 6681 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05315 8787 6708 6556 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05314 6708 6681 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05313 8787 6681 6708 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05312 1231 1318 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05311 1477 1496 1231 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05310 1667 5624 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05309 1876 1753 1667 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05308 5910 6115 5754 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05307 5754 5911 5910 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05306 8787 5908 5754 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05305 7031 7178 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05304 7177 7582 7031 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05303 5552 5634 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05302 6138 5551 5552 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05301 6464 7315 6465 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05300 6465 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05299 6728 8160 6464 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05298 8787 3414 1626 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05297 1752 1755 1624 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05296 1748 2138 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_05295 1624 1746 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05294 1626 1747 1625 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05293 1625 2138 1752 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05292 1752 1748 1627 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05291 2133 1752 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05290 8787 3414 1746 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_05289 1627 1945 1626 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05288 3087 3106 3086 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05287 3086 3668 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05286 3084 3082 3087 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05285 3085 3083 3084 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05284 3395 3832 3075 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05283 3075 3655 3395 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05282 8787 3654 3075 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05281 4884 5465 4885 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05280 4885 5013 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05279 4883 6021 4884 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05278 5209 6514 4883 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05277 8787 5557 5316 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05276 5316 5438 5439 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05275 8132 5439 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05274 3652 4662 3562 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05273 3562 4258 3652 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05272 8787 4064 3562 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05271 3438 3490 3439 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05270 3439 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05269 3437 6026 3438 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05268 3685 3436 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05267 3436 3435 3437 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05266 5982 8065 7311 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05265 8787 8065 5984 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05264 5983 6691 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05263 7311 5984 5983 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05262 8787 6234 5982 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05261 7041 8030 7042 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05260 7042 7593 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05259 7040 7184 7041 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05258 7770 8240 7040 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05257 8787 8487 7393 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05256 7393 7391 7392 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05255 8026 7392 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05254 4291 4320 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05253 5166 4292 4291 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05252 4290 4520 5166 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05251 8787 4289 4290 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05250 4290 5169 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05249 8787 3509 2838 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05248 2838 2972 2973 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05247 2978 2973 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05246 4539 4747 4422 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05245 8787 4758 4540 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05244 4422 4540 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05243 7156 7157 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05242 8787 7156 7009 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05241 7009 7163 7157 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05240 7157 7162 7011 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05239 8787 8728 7162 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05238 7163 7162 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05237 8787 7010 7161 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05236 7011 7047 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05235 7154 7163 7156 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05234 7008 7162 7154 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05233 8787 7153 7008 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05232 7153 7154 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05231 8787 7154 7153 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05230 1488 2277 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05229 1487 2937 1488 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05228 8787 1956 1487 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05227 3053 6286 3054 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05226 3054 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05225 3052 3767 3053 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05224 3171 3169 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05223 3169 3051 3052 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05222 7397 8235 7399 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05221 7399 8236 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05220 7398 7394 7397 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05219 8027 7396 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05218 7396 7395 7398 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05217 7414 8553 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05216 7486 7643 7414 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05215 8787 7485 7486 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05214 8325 7486 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05213 8787 6816 7686 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05212 7686 6874 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05211 8787 6893 7686 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05210 4203 4205 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05209 8787 4203 4204 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05208 4204 4243 4205 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05207 4205 4244 4240 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05206 8787 6232 4244 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05205 4243 4244 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05204 8787 4241 4242 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05203 4240 4239 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05202 4238 4243 4203 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05201 4202 4244 4238 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05200 8787 5790 4202 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05199 5790 4238 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05198 8787 4238 5790 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05197 4813 4816 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05196 8787 4813 4814 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05195 4814 4820 4816 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05194 4816 4821 4817 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05193 8787 6361 4821 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05192 4820 4821 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05191 8787 4818 4819 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05190 4817 4815 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05189 4811 4820 4813 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05188 4812 4821 4811 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05187 8787 5263 4812 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05186 5263 4811 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05185 8787 4811 5263 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05184 4773 5010 4774 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05183 4774 5893 4773 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05182 8787 5014 4774 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05181 3012 3341 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_05180 8787 3011 3012 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_05179 3012 3544 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_05178 8787 3551 3012 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_05177 2501 2505 2257 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05176 2257 2504 2501 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05175 8787 2260 2257 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05174 2824 3083 2823 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05173 2823 3479 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05172 2936 2940 2824 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05171 7284 7283 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05170 7680 7282 7284 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05169 6546 6673 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05168 6668 8490 6546 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05167 7281 7279 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05166 8646 7280 7281 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05165 8068 8069 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05164 8116 8350 8068 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05163 5796 5798 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05162 8787 5796 5713 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05161 5713 5801 5798 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05160 5798 5802 5712 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05159 8787 6232 5802 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05158 5801 5802 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05157 8787 5714 5800 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05156 5712 5774 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05155 5795 5801 5796 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05154 5711 5802 5795 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05153 8787 6311 5711 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05152 6311 5795 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05151 8787 5795 6311 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05150 2699 2515 2407 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05149 2407 2518 2699 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05148 8787 2706 2407 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05147 2663 3102 2665 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05146 2665 3092 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05145 2664 3254 2663 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05144 2965 2955 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05143 2873 6021 2955 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05142 2955 3297 2872 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05141 2872 3531 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05140 8787 3295 2873 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05139 2873 3137 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05138 3545 3968 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05137 3544 3973 3545 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05136 7355 7353 7354 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05135 7354 7576 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05134 7356 7592 7355 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05133 5966 5584 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05132 8787 6934 5585 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05131 5583 5580 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05130 5584 5585 5583 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05129 5582 6934 5584 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05128 8787 5958 5582 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05127 5543 5372 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05126 8787 6934 5374 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05125 5297 5371 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05124 5372 5374 5297 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05123 5296 6934 5372 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05122 8787 6271 5296 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05121 3093 3678 3094 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05120 3094 3677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05119 3092 8168 3093 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05118 8787 3106 2814 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05117 2814 3668 2921 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05116 3073 2921 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05115 2865 3471 2864 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05114 2864 3478 2946 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05113 8787 3885 2865 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05112 2945 2946 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05111 3520 6092 3521 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05110 3521 3762 3520 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05109 8787 3761 3521 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05108 3519 3520 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05107 7023 7169 7024 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05106 7024 7373 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05105 7170 8478 7023 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05104 8787 7305 7299 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05103 7299 7297 7298 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05102 7657 7298 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05101 4464 4246 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05100 8787 6934 4248 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05099 4249 4247 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05098 4246 4248 4249 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05097 4245 6934 4246 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05096 8787 6022 4245 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05095 461 2974 460 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05094 460 805 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05093 612 4358 461 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05092 6597 8030 6596 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05091 6596 7391 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05090 6662 6964 6597 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05089 6143 6234 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05088 6238 8065 6143 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05087 3871 6282 3870 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05086 3870 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05085 3869 4300 3871 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05084 4099 4522 3869 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05083 6144 6410 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05082 6242 8065 6144 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05081 5989 7880 5716 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05080 5716 6007 5989 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05079 8787 6311 5716 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05078 7280 7278 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05077 7278 7521 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05076 8787 7880 7278 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05075 7278 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05074 8787 7877 7278 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05073 8787 4530 2052 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05072 2052 4529 2144 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05071 2532 2144 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05070 5812 5814 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05069 5814 5817 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05068 8787 7273 5814 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05067 5814 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05066 8787 7877 5814 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05065 8787 4955 4692 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05064 4692 4949 4691 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05063 4690 4691 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05062 4843 4929 4844 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05061 4844 4928 4930 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05060 8787 5415 4843 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05059 4927 4930 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05058 7371 7394 7370 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05057 7370 8098 7372 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05056 8787 8247 7371 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05055 7592 7372 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05054 6504 6507 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05053 8787 6504 6505 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05052 6505 6511 6507 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05051 6507 6513 6508 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05050 8787 6512 6513 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05049 6511 6513 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05048 8787 6509 6510 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05047 6508 6506 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05046 6502 6511 6504 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05045 6503 6513 6502 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05044 8787 6758 6503 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05043 6758 6502 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05042 8787 6502 6758 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05041 1308 1462 849 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05040 849 1463 1308 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05039 8787 2260 849 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05038 5810 7049 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05037 889 6285 890 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05036 890 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05035 888 4109 889 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05034 1189 1036 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05033 1036 887 888 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05032 6343 6345 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05031 8787 6343 6195 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05030 6195 6349 6345 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05029 6345 6350 6194 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05028 8787 6361 6350 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05027 6349 6350 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05026 8787 6196 6348 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05025 6194 6219 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05024 6342 6349 6343 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05023 6193 6350 6342 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05022 8787 6339 6193 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05021 6339 6342 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05020 8787 6342 6339 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05019 5174 5826 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05018 4799 5498 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05017 6654 7153 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05016 6153 7315 6152 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05015 6152 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05014 6426 6251 6153 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05013 2858 4286 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05012 2939 2938 2858 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05011 6433 6271 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05010 6003 7315 6004 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05009 6004 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05008 6257 6005 6003 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05007 8787 6925 2828 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05006 2828 2949 2943 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05005 2942 2943 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05004 7840 8098 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05003 8018 8247 7840 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05002 5741 5888 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05001 5889 5892 5741 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05000 793 791 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04999 791 802 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04998 8787 794 791 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04997 791 795 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04996 8787 792 791 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04995 685 4027 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04994 684 1363 685 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04993 7560 7325 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04992 8787 8423 7328 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04991 7327 7326 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04990 7325 7328 7327 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04989 7324 8423 7325 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04988 8787 7553 7324 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04987 8404 8171 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04986 8787 8423 8172 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04985 8170 8168 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04984 8171 8172 8170 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04983 8169 8423 8171 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04982 8787 8399 8169 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04981 7135 6905 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04980 8787 8423 6906 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04979 6904 7142 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04978 6905 6906 6904 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04977 6903 8423 6905 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04976 8787 7140 6903 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04975 3109 3490 3108 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04974 3108 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04973 3107 6716 3109 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04972 3106 8572 3107 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04971 7282 7307 6998 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04970 6998 7308 7282 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04969 8787 7718 6998 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04968 5292 6115 5276 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04967 5276 5914 5292 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04966 8787 5275 5276 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04965 8684 8413 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04964 8787 8423 8415 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04963 8182 8412 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04962 8413 8415 8182 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04961 8179 8423 8413 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04960 8787 8677 8179 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04959 8781 8181 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04958 8787 8430 8183 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04957 8180 8412 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04956 8181 8183 8180 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04955 8178 8430 8181 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04954 8787 8677 8178 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04953 4874 4988 4875 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04952 4875 6878 4989 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04951 8787 6077 4874 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04950 4987 4989 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04949 2002 1998 2003 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04948 2003 2172 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04947 2001 1999 2002 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04946 2772 2000 2001 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04945 4411 4527 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04944 8787 4527 4528 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04943 4526 4524 4411 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04942 4410 4528 4526 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04941 8787 6279 4410 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04940 4524 6279 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04939 3273 6288 3201 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04938 3201 5408 3273 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04937 8787 5631 3201 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04936 7142 6735 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04935 2438 2570 2437 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04934 2437 2569 2568 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04933 8787 2756 2438 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04932 2567 2568 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04931 572 575 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04930 8787 572 447 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04929 447 576 575 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04928 575 578 448 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04927 8787 1516 578 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04926 576 578 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04925 8787 469 577 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04924 448 489 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04923 571 576 572 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04922 446 578 571 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04921 8787 1124 446 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04920 1124 571 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04919 8787 571 1124 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04918 5656 6514 5219 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04917 5219 5218 5656 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04916 8787 5216 5219 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04915 6807 6809 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04914 8787 6807 6808 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04913 6808 6810 6809 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04912 6809 6855 6854 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04911 8787 8596 6855 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04910 6810 6855 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04909 8787 6856 6857 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04908 6854 6853 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04907 6851 6810 6807 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04906 6806 6855 6851 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04905 8787 6852 6806 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04904 6852 6851 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04903 8787 6851 6852 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04902 688 1558 689 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04901 689 1020 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04900 687 1769 688 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04899 805 804 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04898 804 806 687 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04897 4569 4572 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04896 8787 4569 4440 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04895 4440 4575 4572 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04894 4572 4576 4439 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04893 8787 6361 4576 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04892 4575 4576 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04891 8787 4441 4574 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04890 4439 4455 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04889 4567 4575 4569 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04888 4438 4576 4567 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04887 8787 4754 4438 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04886 4754 4567 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04885 8787 4567 4754 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04884 150 152 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04883 8787 150 37 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04882 37 154 152 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04881 152 156 36 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04880 8787 1516 156 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04879 154 156 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04878 8787 38 155 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04877 36 149 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04876 148 154 150 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04875 35 156 148 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04874 8787 992 35 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04873 992 148 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04872 8787 148 992 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04871 4328 4799 4329 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04870 4329 4327 4328 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04869 8787 4334 4329 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04868 6821 6288 6177 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04867 6177 6873 6821 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04866 8787 6287 6177 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04865 5987 5988 5986 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04864 5986 6246 5987 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04863 8787 6235 5986 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04862 5985 5987 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04861 7687 7686 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04860 8665 7688 7687 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04859 4777 4781 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04858 8787 4777 4782 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04857 4782 4785 4781 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04856 4781 4786 4780 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04855 8787 6512 4786 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04854 4785 4786 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04853 8787 4783 4784 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04852 4780 4779 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04851 4776 4785 4777 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04850 4775 4786 4776 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04849 8787 5870 4775 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04848 5870 4776 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04847 8787 4776 5870 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04846 3550 4153 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04845 3551 3979 3550 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04844 5976 5980 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04843 8787 6934 5981 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04842 5979 5978 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04841 5980 5981 5979 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04840 5977 6934 5980 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04839 8787 6311 5977 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04838 3838 2247 2035 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04837 2035 2248 3838 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04836 8787 2260 2035 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04835 8353 8625 8268 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04834 8268 8623 8353 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04833 8787 8627 8268 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04832 8622 8353 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04831 4673 4260 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04830 8787 6934 4261 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04829 4259 4258 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04828 4260 4261 4259 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04827 4257 6934 4260 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04826 8787 6283 4257 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04825 3460 3283 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04824 3283 3282 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04823 8787 3285 3283 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04822 457 5471 458 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04821 458 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04820 1021 1009 457 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04819 7026 8490 7025 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04818 7025 7593 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04817 7171 7173 7026 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04816 3828 2916 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04815 2848 3654 2916 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04814 2916 3658 2849 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04813 2849 3657 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04812 8787 3832 2848 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04811 2848 3655 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04810 8787 166 168 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04809 166 1203 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04808 168 5470 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04807 8294 8474 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04806 8453 8459 8294 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04805 8787 8764 8453 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04804 8451 8453 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04803 5865 6316 5735 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04802 8787 6283 5855 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04801 5735 5855 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04800 2070 6307 2072 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04799 2072 2337 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04798 2071 2760 2070 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04797 2157 2158 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04796 2158 2069 2071 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04795 1616 2255 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04794 1722 2127 1616 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04793 8787 1956 1722 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04792 7093 6843 6566 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04791 6566 6873 7093 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04790 8787 6711 6566 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04789 8787 1105 1107 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04788 1107 5214 1106 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04787 2505 1106 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04786 8604 8603 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04785 8601 8602 8604 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04784 8787 8599 8601 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04783 8600 8601 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04782 298 301 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04781 8787 298 300 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04780 300 304 301 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04779 301 306 302 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04778 8787 1516 306 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04777 304 306 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04776 8787 303 305 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04775 302 299 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04774 297 304 298 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04773 296 306 297 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04772 8787 548 296 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04771 548 297 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04770 8787 297 548 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04769 6211 6373 6212 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04768 6212 6374 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04767 6210 6666 6211 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04766 6372 6375 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04765 6375 6209 6210 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04764 695 3753 694 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04763 694 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04762 693 3490 695 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04761 827 825 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04760 825 826 693 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04759 3916 3964 3918 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04758 3918 6717 3917 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04757 8787 5562 3916 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04756 3915 3917 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04755 8787 8000 6319 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04754 6319 7345 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04753 8787 6316 6319 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04752 8787 8317 8567 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04751 8317 8572 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04750 8567 8350 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04749 1349 1350 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04748 8787 1349 1246 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04747 1246 1355 1350 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04746 1350 1356 1248 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04745 8787 1367 1356 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04744 1355 1356 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04743 8787 1247 1354 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04742 1248 1352 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04741 1347 1355 1349 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04740 1245 1356 1347 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04739 8787 1522 1245 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04738 1522 1347 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04737 8787 1347 1522 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04736 1913 1924 1912 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04735 1912 2128 1913 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04734 8787 1910 1912 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04733 1911 1913 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04732 2498 2125 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04731 2125 2124 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04730 8787 3433 2125 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04729 6720 6311 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04728 6872 6022 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04727 6843 6290 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04726 8651 8652 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04725 8787 8651 8653 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04724 8653 8659 8652 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04723 8652 8660 8654 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04722 8787 8674 8660 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04721 8659 8660 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04720 8787 8656 8658 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04719 8654 8657 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04718 8650 8659 8651 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04717 8649 8660 8650 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04716 8787 8648 8649 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04715 8648 8650 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04714 8787 8650 8648 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04713 2182 1790 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04712 8787 1996 2182 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04711 2182 1791 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04710 8787 1995 2182 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04709 6279 6283 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04708 4473 4943 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04707 2346 1193 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04706 8787 1189 2346 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04705 2346 1373 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04704 8787 1372 2346 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04703 4509 4511 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04702 8787 4509 4403 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04701 4403 4514 4511 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04700 4511 4515 4402 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04699 8787 5835 4515 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04698 4514 4515 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04697 8787 4404 4513 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04696 4402 4453 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04695 4508 4514 4509 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04694 4401 4515 4508 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04693 8787 4715 4401 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04692 4715 4508 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04691 8787 4508 4715 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04690 7126 3140 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04689 3139 3745 3140 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04688 3140 3136 3138 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04687 3138 3137 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04686 8787 3531 3139 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04685 3139 3753 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04684 1672 4109 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04683 1977 3956 1672 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04682 4011 6285 4010 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04681 4010 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04680 4792 6716 4011 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04679 4001 6282 4002 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04678 4002 4111 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04677 4541 6716 4001 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04676 5551 2252 2250 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04675 2250 2251 5551 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04674 8787 2723 2250 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04673 1561 6282 1562 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04672 1562 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04671 2305 3767 1561 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04670 8711 8422 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04669 8787 8423 8425 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04668 8196 8427 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04667 8422 8425 8196 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04666 8194 8423 8422 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04665 8787 8703 8194 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04664 8787 6878 3998 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04663 3998 4099 4100 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04662 4295 4100 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04661 2674 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04660 2672 2926 2674 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04659 2673 2675 2672 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04658 8787 3655 2673 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04657 2673 2671 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04656 8209 8174 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04655 8787 8430 8177 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04654 8176 8175 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04653 8174 8177 8176 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04652 8173 8430 8174 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04651 8787 8410 8173 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04650 8782 8429 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04649 8787 8430 8431 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04648 8201 8427 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04647 8429 8431 8201 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04646 8198 8430 8429 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04645 8787 8703 8198 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04644 8787 637 638 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04643 637 8350 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04642 638 3158 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04641 4446 5563 4445 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04640 4445 5465 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04639 4444 6284 4446 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04638 4579 8065 4444 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04637 8787 3414 1485 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04636 1484 1915 1481 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04635 1486 1755 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_04634 1481 1480 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04633 1485 1479 1483 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04632 1483 1755 1484 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04631 1484 1486 1482 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04630 1737 1484 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04629 8787 3414 1480 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_04628 1482 1487 1485 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04627 8223 8203 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04626 8787 8430 8204 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04625 8205 8202 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04624 8203 8204 8205 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04623 8200 8430 8203 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04622 8787 8199 8200 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04621 8787 3286 3462 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04620 3286 3463 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04619 3462 3285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04618 8561 8315 8250 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04617 8250 8321 8561 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04616 8787 8314 8250 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04615 2807 2904 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04614 8787 2904 2902 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04613 4247 2903 2807 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04612 2806 2902 4247 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04611 8787 2911 2806 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04610 2903 2911 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04609 1914 1919 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04608 1920 1917 1919 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04607 1919 5676 1918 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04606 1918 2949 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04605 8787 1915 1920 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04604 1920 1916 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04603 7955 7957 7797 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04602 7797 8369 7955 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04601 8787 8065 7797 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04600 7875 7955 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04599 5618 8586 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04598 5619 5617 5618 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04597 8787 5843 5616 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04596 5616 6311 5619 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04595 8787 7049 5615 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04594 5615 5844 5619 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04593 7546 7274 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04592 7274 7658 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04591 8787 7273 7274 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04590 7274 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04589 8787 7877 7274 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04588 6489 8000 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04587 6934 8065 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04586 4563 5036 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04585 8787 6717 867 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04584 867 6718 1008 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04583 2542 1008 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04582 8787 5812 5302 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04581 5302 5803 5392 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04580 5390 5392 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04579 6690 6708 6608 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04578 8787 8065 6689 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04577 6608 6689 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04576 5728 7947 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04575 5841 5839 5728 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04574 8787 5843 5726 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04573 5726 6271 5841 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04572 8787 8553 5727 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04571 5727 5844 5841 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04570 6312 6316 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04569 4558 4747 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04568 8571 8570 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04567 8568 8569 8571 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04566 8787 8567 8568 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04565 8577 8568 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04564 3921 3925 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04563 8787 3921 3924 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04562 3924 3929 3925 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04561 3925 3930 3923 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04560 8787 4121 3930 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04559 3929 3930 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04558 8787 3926 3928 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04557 3923 3922 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04556 3920 3929 3921 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04555 3919 3930 3920 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04554 8787 4747 3919 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04553 4747 3920 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04552 8787 3920 4747 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04551 3561 3650 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04550 4059 3651 3561 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04549 1686 6285 1687 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04548 1687 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04547 1685 6718 1686 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04546 1870 1797 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04545 1797 1684 1685 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04544 7127 3134 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04543 3132 5192 3134 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04542 3134 3133 3135 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04541 3135 6021 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04540 8787 3294 3132 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04539 3132 3295 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04538 8787 7635 7850 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04537 7635 8103 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04536 7850 8627 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04535 8787 2980 2981 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04534 2980 2978 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04533 2981 2979 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04532 7949 7950 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04531 8787 7949 7793 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04530 7793 7948 7950 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04529 7950 7953 7794 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04528 8787 8674 7953 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04527 7948 7953 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04526 8787 7795 7952 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04525 7794 7871 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04524 7945 7948 7949 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04523 7792 7953 7945 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04522 8787 7947 7792 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04521 7947 7945 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04520 8787 7945 7947 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04519 8276 8368 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04518 8371 8369 8276 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04517 8787 8366 8371 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04516 8367 8371 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04515 4516 4718 4405 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04514 4405 4519 4516 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04513 8787 4706 4405 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04512 8064 8346 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04511 8063 8347 8064 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04510 2083 3960 2084 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04509 2084 2764 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04508 2573 3767 2083 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04507 6108 7353 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04506 6107 7592 6108 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04505 8787 6817 7691 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04504 7691 6818 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04503 8787 6900 7691 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04502 4668 4670 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04501 8787 4668 4672 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04500 4672 4676 4670 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04499 4670 4677 4671 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04498 8787 6232 4677 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04497 4676 4677 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04496 8787 4674 4675 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04495 4671 4669 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04494 4667 4676 4668 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04493 4666 4677 4667 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04492 8787 6283 4666 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04491 6283 4667 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04490 8787 4667 6283 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04489 2812 3106 2813 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04488 2813 3668 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04487 2920 3254 2812 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04486 2456 3960 2455 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04485 2455 2764 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04484 2798 2586 2456 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04483 7441 8246 7442 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04482 7442 8098 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04481 7574 8237 7441 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04480 8787 4342 4343 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04479 4343 4564 4344 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04478 4788 4344 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04477 3204 5013 3205 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04476 3205 6286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04475 3203 6021 3204 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04474 3275 4715 3203 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04473 3568 3678 3569 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04472 3569 3677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04471 3668 7718 3568 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04470 3474 3885 3473 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04469 3473 3471 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04468 3472 4999 3474 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04467 8211 8782 8210 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04466 8210 8209 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04465 8455 8780 8211 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04464 7653 7933 7652 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04463 7652 8132 7653 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04462 8787 7932 7652 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04461 7930 7653 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04460 7492 8121 7269 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04459 8787 8627 7270 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04458 7269 7270 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04457 4744 5643 4743 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04456 4743 5644 4744 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04455 8787 4754 4743 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04454 7832 8566 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04453 7884 8135 7832 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04452 6603 8490 6604 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04451 6604 7184 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04450 6602 6964 6603 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04449 6672 8240 6602 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04448 8787 4792 3227 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04447 3227 3493 3306 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04446 3305 3306 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04445 7651 8585 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04444 7650 8627 7651 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04443 5411 7880 5307 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04442 5307 6007 5411 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04441 8787 5851 5307 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04440 8787 5446 5447 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04439 5853 5447 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04438 8787 5447 5853 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04437 8787 5447 5853 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04436 5853 5447 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04435 8787 5853 5852 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04434 6272 5852 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04433 8787 5852 6272 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04432 8787 5852 6272 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04431 6272 5852 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04430 8787 5853 5854 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04429 7315 5854 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04428 8787 5854 7315 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04427 8787 5854 7315 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04426 7315 5854 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04425 8787 195 194 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04424 193 194 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04423 8787 194 193 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04422 8787 194 193 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04421 193 194 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04420 8787 193 191 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04419 5563 191 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04418 8787 191 5563 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04417 8787 191 5563 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04416 5563 191 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04415 8787 193 192 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04414 5471 192 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04413 8787 192 5471 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04412 8787 192 5471 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04411 5471 192 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04410 8787 1980 459 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04409 459 2159 610 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04408 609 610 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04407 2799 4230 2801 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04406 2801 2847 2800 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04405 8787 2798 2799 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04404 3058 2800 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04403 5704 5702 5705 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04402 5705 6132 5706 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04401 8787 5703 5704 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04400 5957 5706 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04399 1992 1566 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04398 8787 1564 1992 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04397 5435 5436 5315 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04396 5315 6246 5435 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04395 8787 7534 5315 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04394 5434 5435 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04393 5251 5255 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04392 8787 5251 5254 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04391 5254 5258 5255 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04390 5255 5259 5253 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04389 8787 6361 5259 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04388 5258 5259 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04387 8787 5256 5257 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04386 5253 5252 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04385 5250 5258 5251 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04384 5249 5259 5250 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04383 8787 5498 5249 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04382 5498 5250 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04381 8787 5250 5498 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04380 893 3898 894 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04379 894 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04378 892 5013 893 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04377 1382 1039 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04376 1039 891 892 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04375 6723 7118 6576 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04374 6576 7115 6723 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04373 8787 8372 6576 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04372 6816 6723 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04371 4221 4791 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04370 4573 4565 4221 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04369 3254 2538 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04368 8787 2949 2540 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04367 2417 2537 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04366 2538 2540 2417 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04365 2416 2949 2538 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04364 8787 4319 2416 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04363 3673 2141 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04362 8787 2949 2143 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04361 1950 2537 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04360 2141 2143 1950 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04359 1947 2949 2141 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04358 8787 2145 1947 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04357 43 2976 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04356 175 807 43 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04355 51 4346 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04354 181 2974 51 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04353 4864 7315 4863 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04352 4863 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04351 4978 4977 4864 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04350 8787 3414 1451 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04349 1454 2498 1448 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04348 1452 1716 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_04347 1448 1449 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04346 1451 1455 1450 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04345 1450 1716 1454 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04344 1454 1452 1453 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04343 1447 1454 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04342 8787 3414 1449 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_04341 1453 1722 1451 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04340 8787 3078 2660 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04339 2660 2936 2661 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04338 3654 2661 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04337 8787 3838 3565 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04336 3565 4693 3661 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04335 3660 3661 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04334 882 6040 881 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04333 881 4109 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04332 1552 6021 882 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04331 6527 6662 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04330 6526 6661 6527 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04329 5997 6272 5999 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04328 5999 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04327 6252 5998 5997 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04326 2658 2920 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04325 2659 3665 2658 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04324 8787 3257 2659 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04323 1170 5471 1169 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04322 1169 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04321 4529 4300 1170 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04320 6644 6736 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04319 8787 8430 6737 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04318 6583 7073 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04317 6736 6737 6583 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04316 6582 8430 6736 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04315 8787 6910 6582 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04314 7159 6933 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04313 8787 6934 6935 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04312 6932 7367 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04311 6933 6935 6932 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04310 6931 6934 6933 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04309 8787 7153 6931 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04308 6919 6922 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04307 8787 6934 6923 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04306 6924 7169 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04305 6922 6923 6924 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04304 6921 6934 6922 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04303 8787 6920 6921 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04302 3185 3395 3186 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04301 3186 3398 3250 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04300 8787 3411 3185 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04299 3389 3250 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04298 2081 5465 2082 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04297 2082 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04296 2080 5471 2081 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04295 2564 4300 2080 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04294 7394 7319 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04293 8787 8430 7322 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04292 7321 7320 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04291 7319 7322 7321 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04290 7318 8430 7319 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04289 8787 7323 7318 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04288 502 504 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04287 8787 988 506 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04286 421 4068 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04285 504 506 421 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04284 420 988 504 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04283 8787 721 420 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04282 8787 8227 8228 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04281 8228 8487 8229 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04280 8458 8229 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04279 6321 7735 6186 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04278 6186 6889 6321 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04277 8787 6466 6186 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04276 6320 6321 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04275 3267 6859 3196 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04274 3196 5408 3267 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04273 8787 6265 3196 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04272 3266 3267 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04271 7780 7857 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04270 7923 8063 7780 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04269 8787 7855 7923 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04268 8061 7923 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04267 4546 4548 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04266 8787 4546 4425 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04265 4425 4550 4548 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04264 4548 4552 4424 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04263 8787 6512 4552 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04262 4550 4552 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04261 8787 4426 4551 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04260 4424 4454 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04259 4545 4550 4546 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04258 4423 4552 4545 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04257 8787 4758 4423 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04256 4758 4545 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04255 8787 4545 4758 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04254 2750 3956 2751 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04253 2751 3898 2752 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04252 8787 2986 2750 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04251 2754 2752 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04250 7019 7358 7020 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04249 7020 7362 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04248 7018 7356 7019 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04247 7165 7166 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04246 7166 7017 7018 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04245 4125 4217 4006 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04244 4006 4126 4125 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04243 8787 4553 4006 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04242 4123 4125 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04241 3619 6718 3621 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04240 3621 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04239 3620 6717 3619 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04238 3763 3764 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04237 3764 3638 3620 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04236 1647 2161 1781 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04235 1781 2890 1647 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04234 8787 1779 1647 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04233 1647 2572 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04232 5194 6718 5193 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04231 5193 6285 5195 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04230 8787 5192 5194 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04229 7308 5195 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04228 7260 7261 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04227 8787 7260 7262 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04226 7262 7268 7261 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04225 7261 7267 7266 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04224 8787 8596 7267 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04223 7268 7267 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04222 8787 7263 7265 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04221 7266 7264 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04220 7258 7268 7260 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04219 7259 7267 7258 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04218 8787 7257 7259 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04217 7257 7258 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04216 8787 7258 7257 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04215 2584 1997 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04214 8787 1037 2584 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04213 8787 2188 3755 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04212 2188 2187 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04211 3755 2189 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04210 7132 7133 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04209 8787 7132 7004 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04208 7004 7139 7133 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04207 7133 7138 7006 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04206 8787 8728 7138 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04205 7139 7138 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04204 8787 7005 7137 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04203 7006 7046 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04202 7130 7139 7132 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04201 7003 7138 7130 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04200 8787 7140 7003 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04199 7140 7130 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04198 8787 7130 7140 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04197 3193 3678 3192 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04196 3192 3677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04195 3400 7142 3193 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04194 4538 5643 4421 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04193 4421 5644 4538 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04192 8787 5870 4421 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04191 8787 1980 1981 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04190 1981 3048 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04189 2769 1982 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04188 1981 2315 1982 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04187 1982 2890 1981 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04186 5200 5205 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04185 8787 5200 5201 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04184 5201 5207 5205 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04183 5205 5208 5206 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04182 8787 6512 5208 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04181 5207 5208 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04180 8787 5202 5204 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04179 5206 5203 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04178 5198 5207 5200 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04177 5199 5208 5198 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04176 8787 5872 5199 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04175 5872 5198 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04174 8787 5198 5872 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04173 1999 1602 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04172 8787 1596 1999 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04171 1999 1590 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04170 8787 1798 1999 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_04169 880 2764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04168 1363 4300 880 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04167 7815 8246 7814 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04166 7814 8236 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04165 7904 8237 7815 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04164 7773 7771 7774 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04163 7774 7912 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04162 7772 7770 7773 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04161 8232 8019 7772 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04160 1623 2277 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04159 1743 2937 1623 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04158 8787 1956 1743 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04157 1744 1743 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04156 3397 3395 3399 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04155 3399 3398 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04154 3396 3411 3397 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04153 2404 2942 2403 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04152 2403 3479 2510 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04151 8787 2940 2404 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04150 2509 2510 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04149 7692 7691 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04148 8768 7690 7692 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04147 6116 8490 6117 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04146 6117 8019 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04145 6115 8240 6116 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04144 7467 7592 7468 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04143 7468 7593 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04142 7466 8488 7467 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04141 7771 8240 7466 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04140 8787 4321 4323 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04139 4323 5557 4322 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04138 4320 4322 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04137 7482 7481 7412 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04136 7412 7480 7482 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04135 8787 8350 7412 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04134 7478 7482 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04133 2805 2804 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04132 2804 2802 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04131 8787 2803 2804 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04130 4385 4476 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04129 8787 4476 4478 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04128 4483 4475 4385 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04127 4384 4478 4483 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04126 8787 6720 4384 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04125 4475 6720 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04124 2038 2117 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04123 8787 2117 2118 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04122 4258 2115 2038 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04121 2037 2118 4258 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04120 8787 2128 2037 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04119 2115 2128 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04118 7531 7529 7426 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04117 7426 7528 7531 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04116 8787 8363 7426 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04115 7678 7531 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04114 8787 5044 3542 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04113 3542 3765 3543 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04112 3541 3543 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04111 3230 3944 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04110 3317 5046 3230 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04109 3229 3516 3317 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04108 8787 3314 3229 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04107 3229 3315 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04106 46 391 45 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04105 45 2976 178 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04104 8787 807 46 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04103 177 178 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04102 3856 6720 3855 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04101 3855 5408 3856 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04100 8787 6268 3855 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04099 3854 3856 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04098 3211 6282 3212 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04097 3212 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04096 3210 4300 3211 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04095 3291 3292 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04094 3292 3209 3210 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04093 84 86 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04092 8787 84 12 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04091 12 89 86 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04090 86 90 13 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04089 8787 1302 90 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04088 89 90 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04087 8787 14 88 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04086 13 83 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04085 82 89 84 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04084 11 90 82 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04083 8787 532 11 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04082 532 82 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04081 8787 82 532 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04080 2862 2945 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04079 3082 2944 2862 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04078 4842 4927 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04077 8787 4927 4926 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04076 4937 4924 4842 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04075 4841 4926 4937 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04074 8787 6433 4841 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04073 4924 6433 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04072 5267 5269 5266 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04071 5266 6115 5267 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04070 8787 5265 5266 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04069 1925 1931 1927 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04068 1927 1926 1925 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04067 8787 1923 1927 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04066 1924 1925 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04065 2396 5406 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04064 2499 2501 2396 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04063 2100 2588 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04062 2192 2376 2100 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04061 4156 4157 4023 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04060 4023 5702 4156 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04059 8787 4154 4023 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04058 4153 4156 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04057 6102 8764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04056 6109 6352 6102 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04055 6178 6290 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04054 6291 6316 6178 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04053 7972 7973 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04052 8787 7972 7801 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04051 7801 7971 7973 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04050 7973 7976 7803 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04049 8787 8674 7976 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04048 7971 7976 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04047 8787 7802 7975 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04046 7803 7891 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04045 7966 7971 7972 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04044 7800 7976 7966 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04043 8787 7969 7800 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04042 7969 7966 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04041 8787 7966 7969 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04040 5271 7347 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04039 5272 5270 5271 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04038 5757 8227 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04037 5914 6940 5757 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04036 7507 7509 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04035 8787 7507 7421 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04034 7421 7512 7509 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04033 7509 7513 7420 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04032 8787 8674 7513 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04031 7512 7513 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04030 8787 7422 7511 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04029 7420 7470 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04028 7506 7512 7507 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04027 7419 7513 7506 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04026 8787 7514 7419 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04025 7514 7506 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04024 8787 7506 7514 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04023 3974 4157 3975 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04022 3975 6966 3974 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04021 8787 3972 3975 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04020 3973 3974 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04019 608 607 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04018 8787 1019 607 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04017 607 492 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04016 8787 684 607 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04015 6151 7315 6150 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04014 6150 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04013 6422 6250 6151 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04012 3222 4109 3221 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04011 3221 6037 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04010 4533 3753 3222 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04009 328 330 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04008 8787 988 332 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04007 331 3709 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04006 330 332 331 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04005 329 988 330 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04004 8787 765 329 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04003 259 261 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04002 8787 988 262 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04001 260 3843 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04000 261 262 260 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03999 258 988 261 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03998 8787 274 258 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03997 291 293 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03996 8787 988 295 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03995 294 3849 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03994 293 295 294 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03993 292 988 293 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03992 8787 538 292 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03991 8787 6307 4901 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03990 5020 8427 4899 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03989 5018 5246 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03988 4899 5016 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03987 4901 5237 4900 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03986 4900 5246 5020 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03985 5020 5018 4902 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03984 5015 5020 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03983 8787 6307 5016 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03982 4902 5790 4901 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03981 3423 3678 3422 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03980 3422 3677 3421 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03979 8787 7718 3423 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03978 3666 3421 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03977 3224 5013 3223 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03976 3223 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03975 3493 5192 3224 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03974 1292 1293 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03973 8787 1525 1296 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03972 1221 4068 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03971 1293 1296 1221 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03970 1220 1525 1293 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03969 8787 1297 1220 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03968 4867 5557 4868 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03967 4868 5438 4983 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03966 8787 4988 4867 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03965 5169 4983 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03964 8787 3467 3468 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03963 4299 3468 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03962 8787 3468 4299 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03961 8787 3468 4299 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03960 4299 3468 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03959 8787 4299 4283 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03958 7273 4283 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03957 8787 4283 7273 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03956 8787 4283 7273 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03955 7273 4283 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03954 8787 3414 1230 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03953 1315 1309 1227 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03952 1313 1915 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03951 1227 1311 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03950 1230 1310 1228 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03949 1228 1915 1315 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03948 1315 1313 1229 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03947 1723 1315 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03946 8787 3414 1311 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03945 1229 1916 1230 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03944 2898 2788 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03943 8787 3000 2788 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03942 2788 2787 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03941 8787 3007 2788 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03940 6564 8135 7320 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03939 8787 8135 6700 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03938 6565 6864 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03937 7320 6700 6565 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03936 8787 6701 6564 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03935 8787 4299 4101 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03934 7880 4101 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03933 8787 4101 7880 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03932 8787 4101 7880 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03931 7880 4101 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03930 2975 4046 2839 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03929 2839 2974 2975 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03928 8787 4138 2839 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03927 2976 2975 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03926 6411 8065 7713 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03925 8787 8065 6413 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03924 6412 6852 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03923 7713 6413 6412 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03922 8787 6410 6411 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03921 4765 5465 4767 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03920 4767 5013 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03919 4766 6026 4765 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03918 5669 4764 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03917 4764 4763 4766 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03916 8787 4541 4542 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03915 5849 4542 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03914 8787 4542 5849 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03913 8787 4542 5849 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03912 5849 4542 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03911 8787 5849 5850 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03910 6254 5850 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03909 8787 5850 6254 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03908 8787 5850 6254 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03907 6254 5850 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03906 8787 5849 4991 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03905 6878 4991 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03904 8787 4991 6878 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03903 8787 4991 6878 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03902 6878 4991 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03901 3836 5785 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03900 8787 5785 3837 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03899 3835 3833 3836 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03898 3834 3837 3835 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03897 8787 3832 3834 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03896 3833 3832 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03895 1906 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03894 1905 1907 1906 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03893 1904 1914 1905 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03892 8787 2122 1904 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03891 1901 1905 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03890 8787 1902 1903 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03889 1903 2120 1905 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03888 1707 2511 1611 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03887 1611 1709 1707 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03886 8787 2936 1611 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03885 1706 1707 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03884 3664 3666 3566 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03883 3566 3685 3664 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03882 8787 3673 3566 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03881 3662 3664 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03880 7361 7358 7360 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03879 7360 7364 7359 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03878 8787 7356 7361 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03877 7357 7359 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03876 105 106 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03875 8787 105 20 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03874 20 111 106 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03873 106 112 22 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03872 8787 1516 112 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03871 111 112 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03870 8787 21 110 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03869 22 108 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03868 103 111 105 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03867 19 112 103 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03866 8787 555 19 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03865 555 103 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03864 8787 103 555 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03863 2913 3639 2809 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03862 2809 4469 2913 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03861 8787 2910 2809 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03860 2911 2913 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03859 1704 1886 1610 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03858 1610 1706 1704 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03857 8787 1710 1610 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03856 1882 1704 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03855 1543 1977 1544 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03854 1544 1978 1543 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03853 8787 1641 1544 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03852 1765 1543 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03851 250 253 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03850 8787 250 251 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03849 251 256 253 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03848 253 257 252 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03847 8787 1302 257 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03846 256 257 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03845 8787 254 255 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03844 252 249 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03843 248 256 250 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03842 247 257 248 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03841 8787 721 247 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03840 721 248 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03839 8787 248 721 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03838 3060 3058 3062 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03837 3062 3061 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03836 3059 3546 3060 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03835 3175 3174 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03834 3174 3057 3059 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03833 1690 2586 1691 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03832 1691 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03831 1689 4109 1690 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03830 1798 1799 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03829 1799 1688 1689 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03828 6889 4754 4428 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03827 4428 4557 6889 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03826 8787 4558 4428 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03825 3249 3247 3184 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03824 3184 3246 3249 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03823 8787 3646 3184 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03822 3641 3249 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03821 3637 3485 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_03820 8787 3484 3637 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_03819 3637 4330 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_03818 8787 4324 3637 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_03817 8787 3285 3126 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03816 3126 3291 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03815 8787 3288 3126 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03814 6729 7118 6578 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03813 6578 7115 6729 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03812 8787 7969 6578 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03811 6820 6729 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03810 8637 8643 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03809 8787 8637 8638 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03808 8638 8645 8643 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03807 8643 8647 8644 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03806 8787 8674 8647 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03805 8645 8647 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03804 8787 8640 8642 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03803 8644 8641 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03802 8635 8645 8637 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03801 8636 8647 8635 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03800 8787 8634 8636 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03799 8634 8635 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03798 8787 8635 8634 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03797 686 2764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03796 1641 3531 686 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03795 1261 2764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03794 1553 2586 1261 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03793 8238 8235 8239 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03792 8239 8236 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03791 8477 8237 8238 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03790 8308 8487 8307 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03789 8307 8486 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03788 8771 8485 8308 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03787 1489 1491 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03786 8787 1928 1493 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03785 1492 3254 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03784 1491 1493 1492 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03783 1490 1928 1491 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03782 8787 3673 1490 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03781 8787 7524 7957 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03780 7524 7522 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03779 7957 7523 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03778 8271 8625 8272 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03777 8272 8362 8360 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03776 8787 8623 8271 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03775 8630 8360 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03774 3206 3280 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03773 3281 4285 3206 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03772 4832 4835 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03771 8787 8764 4837 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03770 4836 6548 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03769 4835 4837 4836 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03768 4834 8764 4835 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03767 8787 4833 4834 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03766 2422 2732 2423 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03765 2423 2550 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03764 2421 2727 2422 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03763 2887 3885 2421 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03762 3771 3530 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03761 3530 3529 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03760 8787 3763 3530 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03759 1119 1114 1115 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03758 1115 1113 1119 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03757 8787 7877 1115 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03756 8335 8116 8118 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03755 8118 8343 8335 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03754 8787 8117 8118 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03753 2311 4532 2312 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03752 2312 3716 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03751 2309 2315 2311 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03750 2307 2310 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03749 2310 2308 2309 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03748 1678 1772 1677 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03747 1677 2160 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03746 1676 2559 1678 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03745 1771 1773 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03744 1773 1675 1676 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03743 6666 6768 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03742 6768 6665 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03741 8787 7749 6768 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03740 7769 8027 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03739 7767 8479 7769 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03738 7768 8490 7767 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03737 8787 8242 7768 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03736 7768 8026 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03735 1015 165 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03734 165 163 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03733 8787 2986 165 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03732 7060 7063 6980 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03731 6980 7243 7060 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03730 8787 7059 6980 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03729 8787 4108 3882 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03728 3882 4105 3883 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03727 3881 3883 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03726 8787 5013 3218 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03725 3218 4536 3299 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03724 3745 3299 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03723 6355 6356 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03722 8787 6355 6198 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03721 6198 6362 6356 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03720 6356 6363 6200 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03719 8787 6361 6363 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03718 6362 6363 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03717 8787 6199 6360 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03716 6200 6220 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03715 6353 6362 6355 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03714 6197 6363 6353 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03713 8787 6352 6197 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03712 6352 6353 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03711 8787 6353 6352 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03710 3940 5562 3939 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03709 3939 6717 3941 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03708 8787 6716 3940 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03707 3942 3941 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03706 2861 2949 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03705 3083 6925 2861 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03704 6955 7175 6956 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03703 6956 7169 6955 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03702 8787 8480 6956 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03701 5223 5228 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03700 8787 5223 5224 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03699 5224 5229 5228 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03698 5228 5232 5227 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03697 8787 6512 5232 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03696 5229 5232 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03695 8787 5225 5230 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03694 5227 5226 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03693 5221 5229 5223 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03692 5222 5232 5221 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03691 8787 5220 5222 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03690 5220 5221 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03689 8787 5221 5220 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03688 6894 7127 6895 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03687 6895 7126 6894 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03686 8787 8168 6895 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03685 6893 6894 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03684 7730 8764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03683 7732 8000 7730 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03682 2048 3678 2049 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03681 2049 3677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03680 2139 8427 2048 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03679 2811 2920 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03678 2918 3665 2811 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03677 8787 3257 2918 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03676 3065 2918 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03675 3945 4139 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03674 3969 3944 3945 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03673 3943 3960 3969 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03672 8787 7115 3943 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03671 3943 3942 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_03670 6215 8478 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03669 6377 8240 6215 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03668 313 315 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03667 8787 983 316 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03666 314 3680 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03665 315 316 314 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03664 312 983 315 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03663 8787 554 312 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03662 5755 8227 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03661 5911 7353 5755 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03660 8787 2707 2408 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03659 2408 2517 2519 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03658 2518 2519 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03657 8787 2501 2397 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03656 2397 5406 2502 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03655 2500 2502 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03654 4796 5562 4798 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03653 4798 5013 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03652 4797 6284 4796 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03651 4795 7905 4797 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03650 3587 3716 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03649 5844 3717 3587 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03648 4920 5280 4921 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03647 4921 6677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03646 4919 8478 4920 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03645 5059 6378 4919 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03644 3534 4109 3533 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03643 3533 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03642 3532 6717 3534 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03641 3547 3531 3532 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03640 920 922 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03639 8787 1525 924 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03638 714 3843 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03637 922 924 714 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03636 711 1525 922 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03635 8787 1092 711 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03634 7443 7741 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03633 7575 7573 7443 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03632 8446 8213 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03631 8212 8217 8213 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03630 8213 8215 8214 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03629 8214 8235 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03628 8787 8226 8212 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03627 8212 8220 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03626 7485 6433 6409 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03625 6409 6860 7485 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03624 8787 6408 6409 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03623 8787 3414 2390 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03622 2488 2499 2388 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03621 2486 2498 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03620 2388 2484 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03619 2390 2666 2389 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03618 2389 2498 2488 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03617 2488 2486 2391 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03616 2662 2488 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03615 8787 3414 2484 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03614 2391 2678 2390 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03613 728 730 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03612 8787 779 731 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03611 729 4068 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03610 730 731 729 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03609 727 779 730 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03608 8787 726 727 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03607 1521 1524 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03606 8787 1525 1527 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03605 1526 3709 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03604 1524 1527 1526 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03603 1523 1525 1524 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03602 8787 1522 1523 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03601 8262 8346 8263 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03600 8263 8349 8340 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03599 8787 8347 8262 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03598 8343 8340 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03597 6448 6446 6450 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03596 6450 6447 6449 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03595 8787 6637 6448 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03594 7288 6449 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03593 6599 8222 6600 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03592 6600 8483 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03591 6598 7394 6599 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03590 6770 8237 6598 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03589 777 782 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03588 8787 779 780 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03587 781 2718 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03586 782 780 781 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03585 778 779 782 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03584 8787 994 778 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03583 8787 4822 4825 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03582 4825 7181 4824 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03581 4823 4824 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03580 4741 4985 4740 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03579 4740 4987 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03578 4742 4984 4741 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03577 7529 4739 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03576 4739 4738 4742 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03575 8787 415 413 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03574 628 413 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03573 8787 413 628 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03572 8787 413 628 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03571 628 413 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03570 8787 628 629 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03569 4111 629 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03568 8787 629 4111 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03567 8787 629 4111 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03566 4111 629 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03565 8787 628 412 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03564 4536 412 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03563 8787 412 4536 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03562 8787 412 4536 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03561 4536 412 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03560 1341 1339 1242 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03559 1242 1338 1341 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03558 8787 2260 1242 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03557 2101 1341 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03556 4592 4593 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03555 8787 4592 4449 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03554 4449 4598 4593 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03553 4593 4597 4451 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03552 8787 6361 4597 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03551 4598 4597 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03550 8787 4450 4596 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03549 4451 4456 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03548 4590 4598 4592 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03547 4448 4597 4590 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03546 8787 4833 4448 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03545 4833 4590 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03544 8787 4590 4833 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03543 2879 3960 2880 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03542 2880 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03541 2878 3767 2879 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03540 3170 3003 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03539 3003 2877 2878 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03538 8787 8780 6944 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03537 6944 8235 6945 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03536 7169 6945 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03535 7718 7311 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03534 8168 7713 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03533 3289 2952 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03532 2871 6021 2952 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03531 2952 3531 2870 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03530 2870 3297 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03529 8787 3294 2871 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03528 2871 3295 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03527 4128 4127 4007 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03526 4007 6934 4128 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03525 8787 8430 4007 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03524 4126 4128 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03523 7723 7320 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03522 696 6717 698 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03521 698 3898 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03520 697 3531 696 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03519 1373 828 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03518 828 829 697 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03517 4387 4483 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03516 8787 4483 4484 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03515 4481 4480 4387 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03514 4386 4484 4481 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03513 8787 4479 4386 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03512 4480 4479 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03511 8387 8389 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03510 8787 8387 8278 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03509 8278 8392 8389 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03508 8389 8391 8280 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03507 8787 8674 8391 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03506 8392 8391 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03505 8787 8279 8390 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03504 8280 8310 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03503 8385 8392 8387 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03502 8277 8391 8385 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03501 8787 8383 8277 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03500 8383 8385 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03499 8787 8385 8383 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03498 3446 4502 3447 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03497 3447 5408 3446 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03496 8787 4096 3447 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03495 3445 3446 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03494 8403 8405 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03493 8787 8403 8282 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03492 8282 8408 8405 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03491 8405 8409 8284 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03490 8787 8728 8409 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03489 8408 8409 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03488 8787 8283 8407 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03487 8284 8311 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03486 8402 8408 8403 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03485 8281 8409 8402 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03484 8787 8399 8281 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03483 8399 8402 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03482 8787 8402 8399 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03481 1120 4968 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03480 2281 1119 1120 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03479 1456 1305 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03478 8787 1709 1307 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03477 1225 3254 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03476 1305 1307 1225 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03475 1224 1709 1305 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03474 8787 3673 1224 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03473 3208 3289 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03472 3290 5440 3208 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03471 1968 1966 1969 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03470 1969 2157 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03469 3484 1967 1968 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03468 8787 2770 2771 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03467 2770 2769 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03466 2771 2997 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03465 4723 4727 4725 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03464 8787 8065 4724 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03463 4725 4724 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03462 8670 8395 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03461 8787 8394 8397 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03460 8166 8716 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03459 8395 8397 8166 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03458 8162 8394 8395 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03457 8787 8661 8162 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03456 8373 8375 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03455 8787 8394 8377 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03454 8146 8665 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03453 8375 8377 8146 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03452 8144 8394 8375 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03451 8787 8372 8144 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03450 7669 7084 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03449 8787 8394 7086 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03448 6866 8617 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03447 7084 7086 6866 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03446 6865 8394 7084 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03445 8787 7660 6865 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03444 6205 8227 6204 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03443 6204 8487 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03442 6203 8030 6205 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03441 6368 8240 6203 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03440 8161 8164 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03439 8787 8394 8167 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03438 8165 8768 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03437 8164 8167 8165 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03436 8163 8394 8164 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03435 8787 8160 8163 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03434 6982 7065 6983 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03433 6983 7252 7064 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03432 8787 7066 6982 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03431 7243 7064 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03430 8787 1921 1922 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03429 1921 3266 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03428 1922 2101 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03427 1164 1553 1165 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03426 1165 4750 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03425 1163 4529 1164 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03424 1538 1162 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03423 1162 1161 1163 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03422 8787 6288 4388 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03421 4388 4487 4486 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03420 4485 4486 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03419 6846 6720 6418 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03418 6418 6860 6846 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03417 8787 6417 6418 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03416 7829 8325 7830 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03415 7830 8324 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03414 7828 8323 7829 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03413 8347 7920 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03412 7920 7827 7828 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03411 1881 2105 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03410 8787 2105 1878 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03409 2107 1877 1881 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03408 1880 1878 2107 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03407 8787 1879 1880 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03406 1877 1879 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03405 8787 959 747 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03404 747 5214 749 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03403 1114 749 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03402 8787 1505 1503 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03401 1503 5214 1504 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03400 2274 1504 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03399 7777 8222 7776 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03398 7776 8236 7775 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03397 8787 8247 7777 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03396 8486 7775 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03395 2963 3531 2744 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03394 2744 3767 2963 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03393 8787 3744 2744 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03392 8787 5142 4855 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03391 4855 4952 4950 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03390 4949 4950 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03389 1806 1809 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03388 8787 1806 1655 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03387 1655 1812 1809 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03386 1809 1811 1656 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03385 8787 2028 1811 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03384 1812 1811 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03383 8787 1692 1810 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03382 1656 1697 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03381 1805 1812 1806 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03380 1654 1811 1805 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03379 8787 5470 1654 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03378 5470 1805 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03377 8787 1805 5470 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03376 3177 4839 3176 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03375 3176 3178 3179 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03374 8787 3546 3177 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03373 3180 3179 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03372 7029 8098 7030 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03371 7030 8097 7176 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03370 8787 8247 7029 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03369 7175 7176 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03368 5125 5127 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03367 8787 5127 5126 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03366 5124 5122 5125 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03365 5123 5126 5124 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03364 8787 6843 5123 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03363 5122 6843 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03362 2707 2710 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03361 2710 2709 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03360 8787 2711 2710 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03359 477 613 478 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03358 478 616 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03357 476 614 477 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03356 5214 615 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03355 615 475 476 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03354 6207 8240 6208 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03353 6208 8478 6371 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03352 8787 8480 6207 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03351 6370 6371 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03350 1195 6040 1194 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03349 1194 4109 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03348 1192 6021 1195 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03347 1193 1191 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03346 1191 1190 1192 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03345 5262 7589 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03344 5261 5912 5262 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03343 8787 5260 5261 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03342 350 354 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03341 8787 350 353 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03340 353 358 354 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03339 354 359 352 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03338 8787 1367 359 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03337 358 359 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03336 8787 355 357 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03335 352 351 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03334 349 358 350 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03333 348 359 349 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03332 8787 767 348 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03331 767 349 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03330 8787 349 767 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03329 486 5562 485 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03328 485 3531 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03327 484 5471 486 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03326 625 626 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03325 626 483 484 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03324 5893 6339 5747 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03323 8787 8717 5894 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03322 5747 5894 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03321 5571 7404 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03320 5683 7353 5571 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03319 5753 7347 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03318 5908 5907 5753 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03317 3450 3455 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03316 8787 3450 3451 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03315 3451 3458 3455 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03314 3455 3459 3456 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03313 8787 3705 3459 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03312 3458 3459 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03311 8787 3453 3457 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03310 3456 3454 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03309 3448 3458 3450 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03308 3449 3459 3448 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03307 8787 4522 3449 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03306 4522 3448 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03305 8787 3448 4522 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03304 2386 5150 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03303 3066 2481 2386 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03302 8787 1586 1795 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03301 1795 1777 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03300 8787 1995 1795 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03299 4236 6670 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03298 4237 5280 4236 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03297 8289 8451 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03296 8444 8443 8289 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03295 799 5562 798 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03294 798 3490 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03293 1159 1009 799 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03292 8787 1496 1495 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03291 1495 1498 1494 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03290 1937 1494 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03289 8787 5790 3143 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03288 3143 3141 3142 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03287 3485 3142 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03286 3536 5044 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03285 3535 4143 3536 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03284 3615 6286 3614 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03283 3614 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03282 3613 6717 3615 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03281 3761 6026 3613 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03280 3618 5013 3617 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03279 3617 6286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03278 3616 6026 3618 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03277 3762 4139 3616 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03276 4417 6718 4416 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03275 4416 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03274 4986 5192 4417 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03273 3709 3711 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03272 8787 4075 3713 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03271 3585 4526 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03270 3711 3713 3585 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03269 3584 4075 3711 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03268 8787 8412 3584 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03267 2284 2286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03266 8787 4530 2288 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03265 2287 8427 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03264 2286 2288 2287 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03263 2285 4530 2286 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03262 8787 5440 2285 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03261 356 346 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03260 8787 779 347 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03259 345 3709 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03258 346 347 345 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03257 344 779 346 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03256 8787 767 344 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03255 534 536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03254 8787 779 537 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03253 431 3843 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03252 536 537 431 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03251 430 779 536 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03250 8787 532 430 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03249 7363 7734 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03248 7362 7578 7363 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03247 3896 5465 3895 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03246 3895 3956 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03245 3894 6021 3896 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03244 4064 3893 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03243 3893 3892 3894 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03242 4073 4076 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03241 8787 4075 4077 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03240 3991 4935 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03239 4076 4077 3991 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03238 3990 4075 4076 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03237 8787 7142 3990 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03236 4413 4984 4414 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03235 4414 4985 4531 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03234 8787 4986 4413 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03233 6860 4531 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03232 1949 2139 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03231 1948 3275 1949 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03230 8787 1956 1948 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03229 1946 1948 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03228 8787 1280 1090 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03227 1090 5214 1091 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03226 2247 1091 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03225 3525 3528 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03224 3528 4152 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03223 8787 3763 3528 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03222 3528 3526 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03221 8787 3527 3528 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03220 3313 3315 3228 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03219 3228 3314 3313 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03218 8787 4563 3228 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03217 3310 3313 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03216 8787 6843 5589 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03215 5589 5587 5588 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03214 5586 5588 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03213 5548 5826 5549 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03212 8787 8065 5550 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03211 5549 5550 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03210 3274 2274 2266 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03209 2266 2273 3274 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03208 8787 7877 2266 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03207 8787 3717 3213 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03206 3213 3716 3293 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03205 3885 3293 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03204 6094 6298 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03203 8787 6298 6093 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03202 6092 6090 6094 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03201 6091 6093 6092 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03200 8787 6654 6091 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03199 6090 6654 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03198 7445 8450 7447 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03197 7447 8209 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03196 7446 8483 7445 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03195 7576 7577 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03194 7577 7444 7446 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03193 5241 7315 5243 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03192 8787 7315 5245 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03191 5242 6307 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03190 5243 5245 5242 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03189 8787 6312 5241 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03188 2246 2664 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03187 2245 3090 2246 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03186 8787 3257 2245 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03185 7491 7493 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03184 7416 7535 7493 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03183 7493 7650 7415 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03182 7415 7492 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03181 8787 7536 7416 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03180 7416 7533 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03179 3121 7127 3119 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03178 3119 7126 3121 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03177 8787 8427 3119 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03176 968 971 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03175 8787 968 857 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03174 857 972 971 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03173 971 974 856 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03172 8787 1516 974 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03171 972 974 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03170 8787 858 973 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03169 856 908 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03168 967 972 968 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03167 855 974 967 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03166 8787 1125 855 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03165 1125 967 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03164 8787 967 1125 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03163 2110 2107 2032 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03162 2032 3652 2110 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03161 8787 2108 2032 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03160 4469 2110 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03159 2419 2732 2420 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03158 2420 2550 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03157 2418 2727 2419 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03156 3120 2541 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03155 2541 2463 2418 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03154 582 584 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03153 8787 582 450 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03152 450 587 584 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03151 584 588 451 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03150 8787 1516 588 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03149 587 588 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03148 8787 470 585 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03147 451 490 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03146 581 587 582 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03145 449 588 581 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03144 8787 993 449 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03143 993 581 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03142 8787 581 993 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03141 1864 2272 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03140 2129 2133 1864 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03139 8556 8560 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03138 8787 8556 8558 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03137 8558 8564 8560 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03136 8560 8565 8559 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03135 8787 8596 8565 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03134 8564 8565 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03133 8787 8562 8563 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03132 8559 8557 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03131 8555 8564 8556 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03130 8554 8565 8555 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03129 8787 8553 8554 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03128 8553 8555 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03127 8787 8555 8553 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03126 6730 7127 6579 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03125 6579 7126 6730 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03124 8787 8417 6579 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03123 6819 6730 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03122 8589 8593 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03121 8787 8589 8591 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03120 8591 8597 8593 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03119 8593 8598 8592 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03118 8787 8596 8598 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03117 8597 8598 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03116 8787 8594 8595 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03115 8592 8590 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03114 8588 8597 8589 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03113 8587 8598 8588 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03112 8787 8586 8587 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03111 8586 8588 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03110 8787 8588 8586 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03109 1132 1127 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03108 1131 1128 1132 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03107 1130 1129 1131 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03106 8787 1124 1130 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03105 2273 1131 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03104 8787 1123 1126 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03103 1126 1125 1131 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03102 6677 8483 6606 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03101 6606 8222 6677 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03100 8787 8247 6606 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03099 7756 7907 7755 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03098 7755 8220 7756 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03097 8787 8455 7755 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03096 3735 3725 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03095 8787 8627 3727 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03094 3593 3750 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03093 3725 3727 3593 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03092 3592 8627 3725 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03091 8787 4305 3592 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03090 2515 2517 2406 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03089 2406 2707 2515 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03088 8787 8627 2406 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03087 8787 5220 2717 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03086 2717 2949 2716 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03085 2715 2716 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03084 8787 3673 3189 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03083 3189 3254 3255 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03082 3257 3255 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03081 366 4111 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03080 369 5563 366 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03079 3848 5390 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03078 4490 3846 3848 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03077 3863 3865 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03076 8787 8394 3868 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03075 3867 3866 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03074 3865 3868 3867 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03073 3864 8394 3865 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03072 8787 6005 3864 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03071 4683 4493 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03070 8787 8394 4494 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03069 4270 4490 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03068 4493 4494 4270 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03067 4269 8394 4493 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03066 8787 6250 4269 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03065 3452 3116 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03064 8787 8394 3118 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03063 3117 3281 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03062 3116 3118 3117 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03061 3115 8394 3116 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03060 8787 4522 3115 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03059 6885 6883 6884 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03058 6884 6887 6886 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03057 8787 6882 6885 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03056 7285 6886 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03055 796 3753 797 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03054 797 6718 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03053 4027 5563 796 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03052 1954 1757 1630 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03051 1630 1758 1954 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03050 8787 7877 1630 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03049 4337 4577 4336 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03048 4336 6040 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03047 4335 5562 4337 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03046 4338 8717 4335 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03045 3693 3442 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03044 8787 8394 3444 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03043 3443 3441 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03042 3442 3444 3443 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03041 3440 8394 3442 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03040 8787 4501 3440 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03039 2527 2280 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03038 8787 8394 2283 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03037 2282 2281 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03036 2280 2283 2282 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03035 2279 8394 2280 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03034 8787 4977 2279 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03033 3777 4157 3633 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03032 3633 5915 3777 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03031 8787 3775 3633 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03030 3776 3777 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03029 1586 1585 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03028 1585 1584 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03027 8787 1592 1585 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03026 5762 7184 5763 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03025 5763 6940 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03024 5761 6677 5762 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03023 6373 8490 5761 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03022 2011 6286 2010 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03021 2010 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03020 2009 3956 2011 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03019 2176 3964 2009 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03018 8787 2572 1991 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03017 1991 3048 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03016 2578 1990 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03015 1991 2161 1990 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03014 1990 2890 1991 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03013 7111 6859 6437 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03012 6437 6873 7111 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03011 8787 6721 6437 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03010 2322 2321 2323 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03009 2323 2743 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03008 2319 2318 2322 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03007 2320 2963 2319 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03006 1534 1766 1536 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03005 1536 1535 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03004 1533 1769 1534 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03003 1975 1768 1533 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03002 5445 5643 5317 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03001 5317 5644 5445 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03000 8787 6466 5317 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02999 8022 7908 7762 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02998 7762 7906 8022 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02997 8787 7761 7762 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02996 6688 6841 6559 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02995 6559 7246 6688 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02994 8787 6690 6559 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02993 8787 5805 5301 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02992 5301 5990 5389 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02991 5388 5389 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02990 4955 4960 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02989 4960 4957 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02988 8787 7880 4960 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02987 4960 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02986 8787 7877 4960 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02985 7842 8235 7841 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02984 7841 8097 8021 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02983 8787 8215 7842 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02982 8487 8021 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02981 6264 7713 6158 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02980 6158 6276 6264 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02979 8787 6879 6158 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02978 6262 6264 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02977 8787 2760 1638 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02976 1638 1772 1767 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02975 1766 1767 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02974 1658 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02973 1702 1890 1658 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02972 1657 1706 1702 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02971 8787 3655 1657 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02970 1657 1710 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02969 379 2974 381 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02968 381 805 380 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02967 8787 4350 379 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02966 378 380 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02965 4962 4963 4857 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02964 4857 6246 4962 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02963 8787 7491 4857 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02962 4961 4962 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02961 5052 5053 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02960 8787 5052 4916 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02959 4916 5057 5053 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02958 5053 5058 4918 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02957 8787 6361 5058 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02956 5057 5058 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02955 8787 4917 5056 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02954 4918 4923 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02953 5050 5057 5052 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02952 4915 5058 5050 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02951 8787 5270 4915 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02950 5270 5050 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02949 8787 5050 5270 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02948 7294 7307 7293 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02947 7293 7308 7294 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02946 8787 8168 7293 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02945 4066 5112 3987 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02944 3987 4247 4066 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02943 8787 4064 3987 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02942 4065 4066 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02941 1597 3898 1598 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02940 1598 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02939 1595 6282 1597 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02938 1596 1594 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02937 1594 1593 1595 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02936 4150 6373 4021 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02935 4021 4157 4150 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02934 8787 4147 4021 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02933 4148 4150 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02932 4208 4210 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02931 8787 4208 4209 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02930 4209 4255 4210 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02929 4210 4256 4253 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02928 8787 6232 4256 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02927 4255 4256 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02926 8787 4251 4254 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02925 4253 4252 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02924 4250 4255 4208 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02923 4207 4256 4250 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02922 8787 4943 4207 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02921 4943 4250 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02920 8787 4250 4943 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02919 6081 6082 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02918 8787 6081 6083 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02917 6083 6088 6082 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02916 6082 6089 6086 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02915 8787 6512 6089 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02914 6088 6089 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02913 8787 6084 6087 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02912 6086 6085 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02911 6080 6088 6081 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02910 6079 6089 6080 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02909 8787 6324 6079 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02908 6324 6080 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02907 8787 6080 6324 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02906 5185 6279 5184 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02905 5184 5408 5185 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02904 8787 6275 5184 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02903 5183 5185 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02902 3721 3897 3590 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02901 3590 7115 3721 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02900 8787 6027 3590 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02899 788 3678 787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02898 787 1013 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02897 786 1147 788 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02896 1150 3678 1148 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02895 1148 1151 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02894 1149 1147 1150 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02893 7843 8022 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02892 8475 8023 7843 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02891 8296 8457 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02890 8459 8458 8296 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02889 8304 8477 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02888 8770 8478 8304 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02887 8787 1496 1223 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02886 1223 1456 1299 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02885 1712 1299 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02884 8787 2936 2387 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02883 2387 2922 2483 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02882 2482 2483 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02881 8787 4107 4108 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02880 4107 6878 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02879 4108 5643 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02878 3056 3175 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02877 3055 3772 3056 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02876 6299 5873 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02875 8787 6920 5875 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02874 5670 5872 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02873 5873 5875 5670 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02872 5667 6920 5873 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02871 8787 5870 5667 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02870 7037 7595 7038 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02869 7038 7182 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02868 7181 7589 7037 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02867 8094 8764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02866 8443 8433 8094 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02865 6039 6718 6038 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02864 6038 6037 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02863 6036 6716 6039 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02862 6455 6311 6036 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02861 2424 3753 2425 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02860 2425 6286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02859 2732 2566 2424 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02858 2574 2890 2443 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02857 2443 2572 2574 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02856 8787 2573 2443 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02855 2576 2574 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02854 3622 3946 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02853 3765 4140 3622 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02852 8787 3950 3765 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02851 4079 2247 2036 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02850 2036 2248 4079 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02849 8787 7877 2036 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02848 6014 6717 6015 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02847 6015 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02846 6013 6021 6014 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02845 6432 7660 6013 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02844 517 519 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02843 8787 983 521 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02842 426 4068 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02841 519 521 426 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02840 425 983 519 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02839 8787 720 425 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02838 8787 3414 2240 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02837 2242 2235 2236 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02836 2239 2499 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02835 2236 2237 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02834 2240 2245 2238 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02833 2238 2499 2242 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02832 2242 2239 2241 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02831 2639 2242 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02830 8787 3414 2237 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02829 2241 3090 2240 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02828 6018 6286 6020 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02827 6020 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02826 6019 6021 6018 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02825 6713 6290 6019 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02824 543 545 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02823 8787 983 547 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02822 436 3849 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02821 545 547 436 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02820 435 983 545 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02819 8787 542 435 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02818 4695 6433 4694 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02817 4694 5408 4695 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02816 8787 4965 4694 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02815 4693 4695 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02814 8787 5445 5308 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02813 5308 5619 5413 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02812 5412 5413 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02811 8787 5415 4397 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02810 4397 4499 4500 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02809 4527 4500 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02808 8787 2570 2085 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02807 2085 2170 2169 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02806 2172 2169 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02805 8787 5818 5715 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02804 5715 5985 5804 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02803 5803 5804 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02802 3146 5563 3145 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02801 3145 3753 3147 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02800 8787 5470 3146 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02799 3144 3147 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02798 8787 8247 7369 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02797 7369 8098 7368 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02796 7367 7368 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02795 5129 5466 5128 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02794 5128 5790 5131 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02793 8787 5415 5129 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02792 5127 5131 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02791 8314 8553 8047 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02790 8787 8627 8048 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02789 8047 8048 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02788 3553 3170 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02787 8787 3171 3553 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02786 8427 8185 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02785 8412 8175 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02784 6591 7165 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02783 6659 6947 6591 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02782 8787 6761 6659 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02781 8787 5864 5665 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02780 5665 7115 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02779 5660 5664 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02778 5665 5877 5664 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02777 5664 5662 5665 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02776 8787 1364 4292 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02775 4292 1362 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02774 8787 1358 4292 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02773 4223 4225 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02772 8787 4223 4224 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02771 4224 4355 4225 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02770 4225 4356 4352 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02769 8787 6361 4356 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02768 4355 4356 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02767 8787 4353 4354 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02766 4352 4351 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02765 4349 4355 4223 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02764 4222 4356 4349 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02763 8787 4350 4222 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02762 4350 4349 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02761 8787 4349 4350 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02760 8787 181 41 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02759 41 374 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02758 1123 171 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02757 41 177 171 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02756 171 179 41 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02755 7323 7987 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02754 7556 7558 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02753 8787 7556 7436 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02752 7436 7561 7558 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02751 7558 7563 7435 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02750 8787 8728 7563 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02749 7561 7563 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02748 8787 7437 7562 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02747 7435 7471 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02746 7555 7561 7556 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02745 7434 7563 7555 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02744 8787 7553 7434 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02743 7553 7555 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02742 8787 7555 7553 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02741 3202 4088 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02740 3441 3274 3202 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02739 8787 4533 4309 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02738 4309 4532 4310 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02737 6276 4310 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02736 2831 4533 2832 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02735 2832 4027 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02734 2949 3300 2831 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02733 4314 5644 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02732 4313 4318 4314 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02731 8787 5643 4313 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02730 6129 8478 6130 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02729 6130 6677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02728 6128 6378 6129 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02727 8787 6878 2079 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02726 2079 3048 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02725 2178 2167 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02724 2079 3716 2167 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02723 2167 2890 2079 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02722 8787 395 396 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02721 395 2986 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02720 396 1567 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02719 3934 6037 3933 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02718 3933 4132 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02717 3932 4109 3934 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02716 3931 6284 3932 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02715 8787 617 815 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02714 617 1567 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02713 815 2986 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02712 5035 5038 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02711 8787 8764 5040 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02710 4910 7382 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02709 5038 5040 4910 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02708 4909 8764 5038 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02707 8787 5036 4909 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02706 3152 3494 3151 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02705 3151 3716 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02704 3153 3493 3152 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02703 3150 4532 3153 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02702 2730 2727 2733 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02701 2733 2732 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02700 2731 3885 2730 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02699 5408 2729 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02698 2729 2728 2731 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02697 3886 4040 3887 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02696 3887 3885 3886 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02695 8787 4313 3887 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02694 3884 3886 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02693 8020 7720 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02692 8787 8430 7721 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02691 7719 7718 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02690 7720 7721 7719 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02689 7717 8430 7720 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02688 8787 7716 7717 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02687 8787 3753 3599 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02686 3599 5192 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02685 7307 3743 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02684 3599 3745 3743 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02683 3743 3744 3599 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02682 1621 1738 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02681 8787 1738 1735 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02680 2117 1734 1621 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02679 1620 1735 2117 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02678 8787 1923 1620 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02677 1734 1923 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02676 3674 3676 3571 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02675 3571 3672 3674 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02674 8787 3673 3571 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02673 3671 3674 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02672 8787 3547 3549 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02671 3549 5059 3548 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02670 3546 3548 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02669 4383 4929 4382 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02668 4382 4473 4474 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02667 8787 5415 4383 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02666 4476 4474 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02665 8787 5415 5140 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02664 5140 5139 5141 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02663 5137 5141 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02662 2363 2364 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02661 8787 2363 2365 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02660 2365 2370 2364 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02659 2364 2371 2369 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02658 8787 3329 2371 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02657 2370 2371 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02656 8787 2366 2368 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02655 2369 2367 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02654 2362 2370 2363 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02653 2361 2371 2362 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02652 8787 2566 2361 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02651 2566 2362 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02650 8787 2362 2566 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02649 3899 6282 3901 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02648 3901 3898 3900 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02647 8787 4577 3899 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02646 3897 3900 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02645 8787 2749 2968 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02644 2968 2958 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02643 8787 2748 2968 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02642 8787 8351 8618 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02641 8351 8605 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02640 8618 8350 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02639 2523 2524 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02638 8787 2523 2410 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02637 2410 2530 2524 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02636 2524 2531 2412 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02635 8787 3705 2531 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02634 2530 2531 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02633 8787 2411 2529 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02632 2412 2526 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02631 2521 2530 2523 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02630 2409 2531 2521 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02629 8787 4977 2409 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02628 4977 2521 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02627 8787 2521 4977 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02626 1570 1574 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02625 8787 1570 1571 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02624 1571 1576 1574 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02623 1574 1578 1575 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02622 8787 2028 1578 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02621 1576 1578 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02620 8787 1572 1577 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02619 1575 1573 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02618 1568 1576 1570 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02617 1569 1578 1568 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02616 8787 1567 1569 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02615 1567 1568 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02614 8787 1568 1567 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02613 1973 2325 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_02612 8787 2555 1973 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_02611 1973 1976 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_02610 8787 2320 1973 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_02609 3980 4157 3981 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02608 3981 5703 3980 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02607 8787 3978 3981 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02606 3979 3980 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02605 803 1552 801 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02604 801 800 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02603 802 1980 803 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02602 4680 4682 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02601 8787 4680 4681 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02600 4681 4688 4682 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02599 4682 4689 4686 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02598 8787 6232 4689 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02597 4688 4689 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02596 8787 4684 4687 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02595 4686 4685 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02594 4679 4688 4680 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02593 4678 4689 4679 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02592 8787 6250 4678 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02591 6250 4679 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02590 8787 4679 6250 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02589 5159 8329 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02588 5160 5158 5159 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02587 8787 5843 5157 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02586 5157 5851 5160 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02585 8787 6708 5156 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02584 5156 5844 5160 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02583 8787 2533 2940 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02582 2533 2532 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02581 2940 2535 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02580 3508 3512 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02579 3509 6092 3508 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02578 811 5465 812 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02577 812 3753 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02576 1980 5471 811 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02575 7534 7538 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02574 7427 7535 7538 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02573 7538 7884 7428 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02572 7428 7887 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02571 8787 7536 7427 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02570 7427 7533 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02569 681 2734 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02568 988 1123 681 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02567 8787 3414 2385 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02566 2478 3066 2382 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02565 2475 2499 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02564 2382 2473 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02563 2385 2476 2383 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02562 2383 2499 2478 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02561 2478 2475 2384 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02560 2645 2478 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02559 8787 3414 2473 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02558 2384 2923 2385 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02557 8134 8359 8133 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02556 8133 8132 8134 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02555 8787 8131 8133 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02554 8356 8134 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02553 2304 4530 2306 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02552 2306 2305 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02551 3285 2334 2304 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02550 5734 6043 5733 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02549 5733 6037 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02548 5732 6716 5734 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02547 6032 5851 5732 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02546 1609 1702 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02545 8787 1702 1698 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02544 2103 1699 1609 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02543 1608 1698 2103 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02542 8787 1710 1608 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02541 1699 1710 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02540 4827 5280 4829 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02539 4829 6677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02538 4828 8478 4827 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02537 4826 8480 4828 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02536 3963 6040 3962 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02535 3962 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02534 3961 3964 3963 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02533 3972 5562 3961 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02532 3849 3851 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02531 8787 4075 3853 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02530 3852 4947 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02529 3851 3853 3852 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02528 3850 4075 3851 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02527 8787 8168 3850 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02526 8787 6307 4905 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02525 5030 8202 4903 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02524 5025 5043 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02523 4903 5026 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02522 4905 5270 4904 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02521 4904 5043 5030 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02520 5030 5025 4906 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02519 5023 5030 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02518 8787 6307 5026 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02517 4906 6288 4905 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02516 3843 3844 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02515 8787 4075 3847 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02514 3845 4481 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02513 3844 3847 3845 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02512 3842 4075 3844 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02511 8787 7326 3842 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02510 2718 2720 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02509 8787 4530 2722 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02508 2721 7723 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02507 2720 2722 2721 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02506 2719 4530 2720 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02505 8787 6027 2719 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02504 3560 3648 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02503 8787 3648 3649 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02502 3822 3645 3560 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02501 3559 3649 3822 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02500 8787 3646 3559 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02499 3645 3646 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02498 7106 7307 7000 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02497 7000 7308 7106 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02496 8787 7142 7000 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02495 2897 2774 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02494 8787 2772 2774 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02493 2774 2773 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02492 8787 3163 2774 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02491 3009 3008 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02490 3008 3544 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02489 8787 3538 3008 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02488 3008 2898 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02487 8787 3525 3008 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02486 6990 8135 7073 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02485 8787 8135 7075 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02484 6991 7257 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02483 7073 7075 6991 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02482 8787 7071 6990 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02481 5173 5175 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02480 5175 5174 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02479 8787 7880 5175 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02478 5175 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02477 8787 7877 5175 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02476 8787 5161 4859 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02475 4859 5153 4969 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02474 4968 4969 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02473 8787 1567 1182 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02472 1182 2986 1183 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02471 2586 1183 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02470 8787 7473 7476 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02469 7473 7472 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02468 7476 8350 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02467 5152 6843 5151 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02466 5151 5408 5152 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02465 8787 6259 5151 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02464 5150 5152 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02463 4560 4754 4429 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02462 4429 4557 4560 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02461 8787 4558 4429 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02460 8010 4560 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02459 8787 4999 2834 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02458 2834 2960 2959 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02457 2962 2959 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02456 3128 3290 3127 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02455 3127 3723 3129 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02454 8787 3126 3128 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02453 3125 3129 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02452 7458 8450 7459 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02451 7459 8781 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02450 7457 8483 7458 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02449 7582 7581 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02448 7581 7456 7457 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02447 8410 8677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02446 6910 7553 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02445 2449 2784 2450 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02444 2450 3960 2581 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02443 8787 3767 2449 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02442 2781 2581 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02441 1077 1080 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02440 8787 1077 1081 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02439 1081 1084 1080 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02438 1080 1085 1079 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02437 8787 1302 1085 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02436 1084 1085 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02435 8787 1082 1083 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02434 1079 1078 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02433 1076 1084 1077 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02432 1075 1085 1076 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02431 8787 1297 1075 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02430 1297 1076 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02429 8787 1076 1297 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02428 4061 4059 3985 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02427 3985 4062 4061 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02426 8787 8627 3985 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02425 5048 5284 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02424 4046 4583 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02423 8472 8461 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02422 1664 1738 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02421 1910 1737 1664 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02420 3191 3258 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02419 3259 3670 3191 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02418 8787 3257 3259 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02417 3415 3259 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02416 6798 6799 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02415 8787 6798 6800 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02414 6800 6801 6799 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02413 6799 6838 6837 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02412 8787 8596 6838 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02411 6801 6838 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02410 8787 6834 6836 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02409 6837 6835 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02408 6833 6801 6798 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02407 6797 6838 6833 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02406 8787 7472 6797 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02405 7472 6833 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02404 8787 6833 7472 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02403 1240 1489 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02402 1479 1496 1240 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02401 4931 5130 4845 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02400 4845 5586 4931 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02399 8787 5119 4845 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02398 4934 4931 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02397 1253 1363 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02396 1364 4792 1253 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02395 1160 1159 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02394 1362 1768 1160 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02393 8058 8060 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02392 8787 8058 8059 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02391 8059 8062 8060 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02390 8060 8113 8112 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02389 8787 8596 8113 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02388 8062 8113 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02387 8787 8114 8115 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02386 8112 8111 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02385 8109 8062 8058 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02384 8057 8113 8109 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02383 8787 8110 8057 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02382 8110 8109 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02381 8787 8109 8110 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02380 8787 7674 7675 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02379 7674 7947 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02378 7675 8065 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02377 1671 1765 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02376 2884 1766 1671 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02375 794 1016 456 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02374 456 7536 794 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02373 8787 6077 456 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02372 2817 3102 2816 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02371 2816 3092 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02370 2815 3082 2817 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02369 2922 3083 2815 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02368 6133 7185 6131 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02367 6131 6677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02366 6132 6378 6133 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02365 8097 7312 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02364 8787 8430 7314 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02363 7313 7311 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02362 7312 7314 7313 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02361 7310 8430 7312 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02360 8787 7547 7310 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02359 8216 8450 8219 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02358 8219 8781 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02357 8218 8483 8216 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02356 8217 8215 8218 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02355 6612 6713 6613 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02354 6613 6715 6712 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02353 8787 6714 6612 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02352 7283 6712 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02351 4018 6029 4019 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02350 4019 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02349 4017 4577 4018 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02348 4147 5013 4017 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02347 8236 7712 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02346 8787 8430 7715 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02345 7714 7713 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02344 7712 7715 7714 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02343 7711 8430 7712 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02342 8787 7895 7711 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02341 3433 6859 3434 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02340 3434 5408 3433 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02339 8787 6265 3434 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02338 1649 3490 1650 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02337 1650 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02336 1648 3531 1649 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02335 2174 5465 1648 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02334 8787 8433 4769 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02333 4769 5011 4770 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02332 4768 4770 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02331 8787 7404 7044 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02330 7044 8487 7186 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02329 7588 7186 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02328 8787 6672 6551 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02327 6551 6553 6550 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02326 6549 6550 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02325 1670 4530 1669 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02324 1669 2305 1764 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02323 8787 2334 1670 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02322 1763 1764 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02321 8787 4139 2840 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02320 2840 3160 2984 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02319 2983 2984 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02318 6538 6644 6539 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02317 6539 8483 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02316 6536 8246 6538 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02315 6537 6535 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02314 6535 6534 6536 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02313 1588 2586 1587 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02312 1587 2764 1589 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02311 8787 4139 1588 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02310 1590 1589 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02309 4895 5471 4894 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02308 4894 5465 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02307 4893 6021 4895 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02306 5011 5012 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02305 5012 4892 4893 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02304 8002 8003 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02303 8787 8002 7811 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02302 7811 8001 8003 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02301 8003 8007 7813 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02300 8787 8728 8007 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02299 8001 8007 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02298 8787 7812 8005 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02297 7813 7902 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02296 7998 8001 8002 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02295 7810 8007 7998 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02294 8787 8000 7810 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02293 8000 7998 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02292 8787 7998 8000 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02291 1727 2511 1617 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02290 1617 1862 1727 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02289 8787 2936 1617 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02288 1902 1727 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02287 4334 4333 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02286 4333 4219 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02285 8787 4795 4333 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02284 769 767 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02283 770 1128 769 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02282 768 1129 770 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02281 8787 764 768 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02280 1758 770 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02279 8787 1123 766 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02278 766 765 770 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02277 5638 5851 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_02276 8787 6311 5638 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_02275 5638 6283 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_02274 8787 5440 5638 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_02273 2301 1973 1974 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02272 1974 1972 2301 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02271 8787 2151 1974 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02270 5379 5381 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02269 8787 5379 5300 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02268 5300 5378 5381 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02267 5381 5385 5299 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02266 8787 6232 5385 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02265 5378 5385 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02264 8787 5342 5384 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02263 5299 5359 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02262 5377 5378 5379 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02261 5298 5385 5377 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02260 8787 6290 5298 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02259 6290 5377 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02258 8787 5377 6290 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02257 8787 5371 3986 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02256 3986 4065 4063 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02255 4062 4063 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02254 7469 8487 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02253 7595 7913 7469 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02252 8787 7594 7595 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02251 4436 7315 4435 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02250 4435 5244 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02249 4564 4563 4436 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02248 2874 3494 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02247 2958 3300 2874 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02246 866 2734 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02245 1525 5214 866 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02244 3977 4157 3976 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02243 3976 5703 3977 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02242 8787 3978 3976 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02241 8293 8483 8292 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02240 8292 8450 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02239 8454 8780 8293 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02238 7819 8019 7818 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02237 7818 8487 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02236 8744 8018 7819 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02235 8787 5856 5658 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02234 5861 6062 5650 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02233 5859 7315 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02232 5650 5857 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02231 5658 6294 5652 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02230 5652 7315 5861 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02229 5861 5859 5653 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02228 6052 5861 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02227 8787 5856 5857 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02226 5653 7718 5658 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02225 874 3753 873 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02224 873 6285 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02223 1535 1203 874 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02222 2327 3956 2329 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02221 2329 3767 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02220 2328 2961 2327 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02219 5339 6940 5340 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02218 5340 7592 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02217 5338 6677 5339 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02216 5702 8490 5338 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02215 5697 7592 5699 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02214 5699 7353 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02213 5698 6677 5697 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02212 5703 8490 5698 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02211 2746 2747 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02210 8787 3144 2747 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02209 2747 4768 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02208 8787 2745 2747 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02207 1618 2508 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02206 1732 3269 1618 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02205 8787 1956 1732 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02204 2787 2345 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02203 8787 2343 2345 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02202 2345 2344 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02201 8787 3156 2345 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02200 6041 6040 6044 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02199 6044 6043 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02198 6042 6716 6041 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02197 6719 8661 6042 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02196 8787 6940 5748 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02195 5748 8030 5896 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02194 5895 5896 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02193 8787 418 419 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02192 1046 419 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02191 8787 419 1046 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02190 8787 419 1046 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02189 1046 419 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02188 8787 1046 1043 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02187 3898 1043 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02186 8787 1043 3898 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02185 8787 1043 3898 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02184 3898 1043 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02183 8787 1046 1047 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02182 4109 1047 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02181 8787 1047 4109 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02180 8787 1047 4109 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02179 4109 1047 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02178 8787 1092 1094 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02177 1094 5214 1093 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02176 1462 1093 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02175 8787 2974 393 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02174 393 4346 394 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02173 614 394 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02172 7401 8488 7403 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02171 7403 8027 7402 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02170 8787 8240 7401 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02169 7400 7402 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02168 5881 5882 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02167 8787 5881 5738 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02166 5738 5886 5882 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02165 5882 5887 5740 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02164 8787 6512 5887 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02163 5886 5887 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02162 8787 5739 5885 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02161 5740 5777 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02160 5879 5886 5881 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02159 5737 5887 5879 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02158 8787 6072 5737 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02157 6072 5879 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02156 8787 5879 6072 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02155 8787 4148 2355 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02154 2355 2354 2356 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02153 2359 2356 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02152 5560 5563 5564 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02151 5564 5562 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02150 5561 6284 5560 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02149 8019 5682 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02148 5682 5559 5561 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02147 1446 1702 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02146 1883 1447 1446 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02145 4031 6717 4030 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02144 4030 4109 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02143 4029 4577 4031 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02142 5643 4110 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02141 4110 4028 4029 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02140 2868 4529 2869 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02139 2869 4750 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02138 2867 6878 2868 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02137 3471 2948 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02136 2948 2866 2867 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02135 6908 7140 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02134 7895 8399 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02133 2961 5470 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02132 8734 8735 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02131 8787 8734 8736 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02130 8736 8742 8735 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02129 8735 8743 8737 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02128 8787 8758 8743 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02127 8742 8743 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02126 8787 8738 8740 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02125 8737 8739 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02124 8733 8742 8734 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02123 8732 8743 8733 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02122 8787 8731 8732 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02121 8731 8733 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02120 8787 8733 8731 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02119 1457 1456 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02118 1455 1496 1457 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02117 1682 2173 1683 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02116 1683 1794 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02115 1681 1795 1682 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02114 3061 1796 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02113 1796 1680 1681 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02112 195 2566 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02111 8787 1390 195 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02110 185 1567 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02109 8787 2986 185 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02108 5996 6251 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02107 5143 5998 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02106 1863 2277 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02105 1928 2937 1863 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02104 2555 2558 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02103 2558 2556 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02102 8787 3150 2558 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02101 4976 6288 4862 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02100 4862 6860 4976 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02099 8787 4974 4862 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02098 4973 4976 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02097 6459 7315 6460 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02096 6460 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02095 6458 8661 6459 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02094 8679 8683 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02093 8787 8679 8682 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02092 8682 8687 8683 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02091 8683 8689 8681 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02090 8787 8728 8689 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02089 8687 8689 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02088 8787 8685 8686 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02087 8681 8680 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02086 8678 8687 8679 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02085 8676 8689 8678 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02084 8787 8677 8676 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02083 8677 8678 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02082 8787 8678 8677 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02081 1668 5183 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02080 1755 1951 1668 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02079 3141 2544 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02078 2426 4300 2544 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02077 2544 3295 2427 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02076 2427 3964 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02075 8787 2542 2426 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02074 2426 3133 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02073 4971 7880 4861 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02072 4861 6007 4971 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02071 8787 5440 4861 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02070 5460 4994 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02069 8787 4997 4996 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02068 4879 7142 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02067 4994 4996 4879 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02066 4878 4997 4994 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02065 8787 6271 4878 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02064 1944 2139 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02063 1945 3275 1944 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02062 8787 1956 1945 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02061 3080 3083 3081 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02060 3081 3082 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02059 3079 3400 3080 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02058 3078 3429 3079 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02057 6567 7315 6568 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02056 6568 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02055 6715 7514 6567 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02054 7817 8450 7816 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02053 7816 8781 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02052 8220 8237 7817 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02051 1679 2784 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02050 2572 3964 1679 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02049 6303 6306 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02048 8787 6307 6308 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02047 6183 7326 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02046 6306 6308 6183 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02045 6182 6307 6306 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02044 8787 6309 6182 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02043 8787 5166 5164 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02042 5164 5171 5165 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02041 7066 5165 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02040 3097 3678 3096 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02039 3096 3677 3098 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02038 8787 8168 3097 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02037 3095 3098 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02036 4015 5563 4014 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02035 4014 5465 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02034 4013 6716 4015 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02033 4138 4833 4013 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02032 6415 6691 6414 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02031 8787 8065 6416 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02030 6414 6416 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02029 8344 8348 8264 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02028 8264 8343 8344 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02027 8787 8350 8264 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02026 8603 8344 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02025 3104 5013 3105 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02024 3105 6286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02023 3103 6021 3104 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02022 3102 7472 3103 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02021 8787 188 190 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02020 188 1390 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02019 190 2566 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02018 8787 8770 8773 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02017 8773 8771 8772 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02016 8769 8772 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02015 5710 5789 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02014 8787 5789 5792 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02013 5974 5788 5710 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02012 5709 5792 5974 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02011 8787 5790 5709 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02010 5788 5790 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02009 3603 3750 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02008 8787 3750 3751 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02007 3749 3747 3603 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02006 3602 3751 3749 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02005 8787 5790 3602 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02004 3747 5790 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02003 4090 4091 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02002 4091 4289 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02001 8787 7880 4091 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02000 4091 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01999 8787 7877 4091 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01998 6594 7367 6595 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01997 6595 8030 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01996 6593 6964 6594 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01995 6661 8240 6593 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01994 4706 4715 4707 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01993 8787 8350 4708 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01992 4707 4708 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01991 8787 4529 3465 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01990 3465 4750 3466 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01989 3463 3466 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01988 8787 4533 3907 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01987 3907 4027 3906 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01986 5010 3906 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01985 8787 5173 4865 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01984 4865 5179 4980 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01983 4979 4980 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01982 7495 7497 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01981 7417 7535 7497 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01980 7497 7648 7418 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01979 7418 7655 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01978 8787 7536 7417 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01977 7417 7533 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01976 4267 4488 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01975 8787 4488 4266 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01974 4279 4265 4267 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01973 4264 4266 4279 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01972 8787 6288 4264 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01971 4265 6288 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01970 2679 2931 2680 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01969 2680 2934 2679 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01968 8787 3673 2680 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01967 2678 2679 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01966 5731 8363 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01965 5848 5845 5731 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01964 8787 5843 5729 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01963 5729 6290 5848 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01962 8787 8572 5730 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01961 5730 5844 5848 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01960 8787 2586 2448 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01959 2448 2764 2580 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01958 3165 2580 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01957 8436 8437 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01956 8787 8436 8286 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01955 8286 8441 8437 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01954 8437 8442 8288 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01953 8787 8728 8442 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01952 8441 8442 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01951 8787 8287 8440 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01950 8288 8312 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01949 8434 8441 8436 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01948 8285 8442 8434 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01947 8787 8433 8285 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01946 8433 8434 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01945 8787 8434 8433 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01944 509 512 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01943 8787 509 423 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01942 423 515 512 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01941 512 516 424 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01940 8787 1302 516 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01939 515 516 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01938 8787 467 514 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01937 424 487 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01936 510 515 509 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01935 422 516 510 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01934 8787 925 422 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01933 925 510 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01932 8787 510 925 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01931 4646 5790 4648 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01930 8787 8350 4647 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01929 4648 4647 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01928 8626 8625 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01927 8624 8623 8626 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01926 3846 2251 2253 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01925 2253 2252 3846 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01924 8787 7877 2253 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01923 3689 3691 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01922 8787 3689 3577 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01921 3577 3695 3691 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01920 3691 3696 3578 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01919 8787 3705 3696 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01918 3695 3696 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01917 8787 3579 3694 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01916 3578 3634 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01915 3688 3695 3689 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01914 3576 3696 3688 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01913 8787 4501 3576 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01912 4501 3688 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01911 8787 3688 4501 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01910 2681 2927 2683 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01909 2683 2933 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01908 2682 3254 2681 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01907 7587 8235 7463 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01906 7463 8246 7587 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01905 8787 8247 7463 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01904 7761 7587 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01903 2822 3678 2821 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01902 2821 3677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01901 2933 7723 2822 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01900 3700 3703 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01899 8787 3700 3581 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01898 3581 3706 3703 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01897 3703 3707 3583 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01896 8787 3705 3707 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01895 3706 3707 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01894 8787 3582 3704 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01893 3583 3635 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01892 3698 3706 3700 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01891 3580 3707 3698 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01890 8787 6005 3580 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01889 6005 3698 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01888 8787 3698 6005 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01887 8787 3414 3408 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01886 3410 3637 3404 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01885 3407 5580 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_01884 3404 3403 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01883 3408 3405 3406 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01882 3406 5580 3410 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01881 3410 3407 3409 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01880 3832 3410 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01879 8787 3414 3403 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_01878 3409 3670 3408 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01877 5268 7353 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01876 5269 7184 5268 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01875 2066 4109 2065 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01874 2065 6037 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01873 2318 6284 2066 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01872 343 2734 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01871 779 1128 343 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01870 6952 7593 6951 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01869 6951 7391 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01868 6950 8030 6952 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01867 8787 6878 6156 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01866 6156 6257 6258 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01865 6858 6258 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01864 8787 3414 3071 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01863 3070 5580 3064 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01862 3067 3066 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_01861 3064 3063 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01860 3071 3065 3068 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01859 3068 3066 3070 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01858 3070 3067 3069 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01857 3644 3070 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01856 8787 3414 3063 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_01855 3069 3662 3071 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01854 7353 8020 7022 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01853 7022 8235 7353 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01852 8787 8237 7022 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01851 8320 8323 8252 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01850 8252 8326 8320 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01849 8787 8627 8252 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01848 8570 8320 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01847 8257 8325 8256 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01846 8256 8324 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01845 8255 8323 8257 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01844 8327 8326 8255 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01843 6441 6438 6440 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01842 6440 6635 6442 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01841 8787 6439 6441 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01840 7099 6442 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01839 6047 6282 6046 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01838 6046 6286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01837 6045 6284 6047 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01836 6287 7969 6045 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01835 8787 815 816 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01834 1173 816 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01833 8787 816 1173 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01832 8787 816 1173 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01831 1173 816 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01830 8787 1173 1174 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01829 3767 1174 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01828 8787 1174 3767 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01827 8787 1174 3767 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01826 3767 1174 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01825 8787 1173 1023 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01824 3753 1023 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01823 8787 1023 3753 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01822 8787 1023 3753 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01821 3753 1023 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01820 8787 1173 1024 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01819 4577 1024 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01818 8787 1024 4577 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01817 8787 1024 4577 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01816 4577 1024 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01815 2378 2672 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01814 8787 2672 2468 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01813 3639 2466 2378 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01812 2377 2468 3639 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01811 8787 2662 2377 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01810 2466 2662 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01809 5196 5643 5197 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01808 5197 5644 5196 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01807 8787 5872 5197 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01806 8787 2559 2340 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01805 2340 2890 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01804 2579 2341 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01803 2340 2760 2341 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01802 2341 3048 2340 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01801 8787 190 187 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01800 621 187 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01799 8787 187 621 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01798 8787 187 621 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01797 621 187 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01796 8787 621 400 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01795 3490 400 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01794 8787 400 3490 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01793 8787 400 3490 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01792 3490 400 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01791 8787 621 622 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01790 5013 622 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01789 8787 622 5013 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01788 8787 622 5013 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01787 5013 622 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01786 8787 621 620 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01785 3956 620 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01784 8787 620 3956 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01783 8787 620 3956 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01782 3956 620 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01781 8787 396 182 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01780 398 182 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01779 8787 182 398 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01778 8787 182 398 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01777 398 182 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01776 8787 398 183 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01775 5192 183 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01774 8787 183 5192 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01773 8787 183 5192 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01772 5192 183 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01771 8787 398 397 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01770 3964 397 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01769 8787 397 3964 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01768 8787 397 3964 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01767 3964 397 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01766 8787 398 399 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01765 3531 399 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01764 8787 399 3531 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01763 8787 399 3531 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01762 3531 399 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01761 8137 8361 8136 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01760 8136 8630 8137 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01759 8787 8135 8136 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01758 8368 8137 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01757 4285 4284 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01756 4284 5428 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01755 8787 7880 4284 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01754 4284 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01753 8787 7877 4284 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01752 7451 8235 7452 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01751 7452 8020 7580 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01750 8787 8237 7451 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01749 7593 7580 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01748 8787 6765 6592 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01747 6592 7171 6764 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01746 6946 6764 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01745 5218 5363 5217 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01744 5217 5214 5218 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01743 8787 5215 5217 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01742 8787 3964 1651 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01741 1651 2784 1800 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01740 2017 1800 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01739 8324 5428 5313 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01738 5313 8132 8324 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01737 8787 5426 5313 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01736 1508 1509 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01735 8787 1508 1510 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01734 1510 1517 1509 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01733 1509 1518 1515 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01732 8787 1516 1518 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01731 1517 1518 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01730 8787 1511 1514 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01729 1515 1512 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01728 1506 1517 1508 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01727 1507 1518 1506 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01726 8787 1505 1507 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01725 1505 1506 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01724 8787 1506 1505 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01723 376 2974 375 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01722 375 805 377 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01721 8787 4358 376 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01720 374 377 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01719 8787 3956 2833 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01718 2833 4109 2957 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01717 3137 2957 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01716 8787 8215 6969 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01715 6969 8222 6971 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01714 6970 6971 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01713 8787 2315 2078 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01712 2078 3048 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01711 2570 2164 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01710 2078 2305 2164 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01709 2164 2890 2078 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01708 6818 6279 6168 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01707 6168 6873 6818 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01706 8787 6462 6168 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01705 1900 1898 1899 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01704 1899 1911 1900 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01703 8787 1901 1899 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01702 2105 1900 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01701 3665 3666 3567 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01700 3567 3685 3665 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01699 8787 3673 3567 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01698 5612 4977 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01697 6006 6005 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01696 7739 8209 7740 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01695 7740 7735 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01694 7737 8782 7739 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01693 7734 7738 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01692 7738 7736 7737 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01691 4794 5023 4793 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01690 4793 5031 4794 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01689 8787 4792 4793 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01688 4791 4794 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01687 8787 6316 5484 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01686 5484 5907 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01685 8787 5565 5484 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01684 1002 1004 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01683 8787 1002 863 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01682 863 1005 1004 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01681 1004 1007 865 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01680 8787 1516 1007 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01679 1005 1007 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01678 8787 864 1006 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01677 865 909 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01676 1001 1005 1002 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01675 862 1007 1001 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01674 8787 1140 862 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01673 1140 1001 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01672 8787 1001 1140 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01671 1659 2255 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01670 1709 2127 1659 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01669 897 6286 898 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01668 898 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01667 896 3964 897 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01666 1592 1040 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01665 1040 895 896 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01664 8128 8605 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01663 7521 8363 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01662 4963 4501 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01661 8787 2320 1972 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01660 1972 1975 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01659 8787 2551 1972 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01658 1226 3854 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01657 1716 1308 1226 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01656 6227 5783 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01655 8787 6934 5786 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01654 5581 5785 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01653 5783 5786 5581 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01652 5579 6934 5783 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01651 8787 6223 5579 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01650 4447 7347 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01649 4822 4580 4447 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01648 3598 3745 4985 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01647 4985 3744 3598 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01646 8787 3739 3598 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01645 3598 3753 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01644 7052 7053 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01643 8787 7052 6977 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01642 6977 7058 7053 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01641 7053 7057 6979 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01640 8787 8596 7057 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01639 7058 7057 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01638 8787 6978 7056 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01637 6979 7045 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01636 7050 7058 7052 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01635 6976 7057 7050 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01634 8787 7049 6976 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01633 7049 7050 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01632 8787 7050 7049 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01631 2039 2119 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01630 2120 2509 2039 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01629 6309 6313 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01628 8787 6312 6315 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01627 6185 6311 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01626 6313 6315 6185 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01625 6184 6312 6313 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01624 8787 6489 6184 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01623 6170 7315 6169 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01622 6169 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01621 6281 7969 6170 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01620 5701 8478 5700 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01619 5700 6677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01618 5917 8480 5701 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01617 4789 4787 4790 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01616 4790 4788 4789 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01615 8787 5015 4790 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01614 5496 5499 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01613 8787 7347 5503 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01612 5333 6526 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01611 5499 5503 5333 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01610 5332 7347 5499 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01609 8787 5498 5332 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01608 6655 6757 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01607 8787 8764 6759 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01606 6590 6760 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01605 6757 6759 6590 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01604 6589 8764 6757 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01603 8787 6758 6589 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01602 5324 5465 5325 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01601 5325 6073 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01600 5323 5471 5324 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01599 5666 6021 5323 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01598 5833 5427 5312 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01597 5312 7066 5833 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01596 8787 5548 5312 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01595 4838 5280 4840 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01594 4840 6674 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01593 4839 6378 4838 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01592 7750 8450 7751 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01591 7751 8235 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01590 7748 8223 7750 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01589 7749 8780 7748 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01588 6874 6872 6875 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01587 6875 6873 6874 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01586 8787 6879 6875 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01585 6076 6077 6075 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01584 8787 6077 6078 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01583 6074 6319 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01582 6075 6078 6074 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01581 8787 6307 6076 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01580 7063 7252 6981 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01579 6981 7246 7063 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01578 8787 8350 6981 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01577 7848 8483 7849 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01576 7849 8236 8031 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01575 8787 8247 7848 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01574 8029 8031 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01573 5633 8202 5632 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01572 5632 6276 5633 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01571 8787 6287 5632 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01570 5631 5633 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01569 2930 2931 2820 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01568 2820 2934 2930 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01567 8787 3673 2820 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01566 6481 6485 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01565 8787 6481 6482 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01564 6482 6487 6485 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01563 6485 6490 6486 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01562 8787 6512 6490 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01561 6487 6490 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01560 8787 6483 6488 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01559 6486 6484 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01558 6479 6487 6481 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01557 6480 6490 6479 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01556 8787 6739 6480 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01555 6739 6479 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01554 8787 6479 6739 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01553 2093 2180 2094 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01552 2094 2179 2181 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01551 8787 2178 2093 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01550 3178 2181 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01549 8787 3049 3527 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01548 3527 3305 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01547 8787 3307 3527 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01546 5490 5493 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01545 8787 5490 5331 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01544 5331 5489 5493 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01543 5493 5495 5330 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01542 8787 6361 5495 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01541 5489 5495 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01540 8787 5353 5494 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01539 5330 5366 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01538 5488 5489 5490 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01537 5329 5495 5488 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01536 8787 5565 5329 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01535 5565 5488 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01534 8787 5488 5565 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01533 7068 6872 6563 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01532 6563 6860 7068 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01531 8787 6699 6563 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01530 4051 4053 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01529 8787 4051 3983 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01528 3983 4050 4053 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01527 4053 4058 3984 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01526 8787 4057 4058 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01525 4050 4058 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01524 8787 4024 4056 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01523 3984 4033 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01522 4049 4050 4051 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01521 3982 4058 4049 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01520 8787 6027 3982 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01519 6027 4049 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01518 8787 4049 6027 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01517 6292 6071 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01516 6071 6070 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01515 8787 6352 6071 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01514 8787 1496 1241 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01513 1241 1489 1334 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01512 1333 1334 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01511 3482 3483 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01510 3483 4324 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01509 8787 3485 3483 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01508 3483 3484 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01507 8787 4330 3483 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01506 8747 8746 8748 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01505 8748 8744 8747 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01504 8787 8745 8748 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01503 6294 6292 6179 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01502 6179 6293 6294 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01501 8787 6291 6179 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01500 7926 8346 7781 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01499 7781 8347 7926 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01498 8787 8065 7781 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01497 7857 7926 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01496 2380 3102 2381 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01495 2381 3092 2472 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01494 8787 3657 2380 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01493 2471 2472 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01492 6135 8030 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01491 6134 8240 6135 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01490 1644 4577 1645 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01489 1645 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01488 2334 5013 1644 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01487 5745 7349 5746 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01486 5746 5891 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01485 5892 8478 5745 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01484 5736 6312 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01483 5877 6307 5736 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01482 8787 7115 5877 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01481 6454 6455 6456 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01480 6456 6458 6457 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01479 8787 6453 6454 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01478 7300 6457 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01477 464 5562 465 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01476 465 3531 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01475 2159 5471 464 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01474 6172 6282 6173 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01473 6173 6286 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01472 6171 6284 6172 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01471 6462 8160 6171 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01470 1037 624 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01469 8787 498 624 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01468 624 499 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01467 8787 625 624 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01466 3467 2950 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01465 2950 2887 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01464 8787 7127 2950 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01463 2950 2884 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01462 8787 7126 2950 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01461 8787 4090 3995 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01460 3995 4703 4089 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01459 4088 4089 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01458 8787 1793 1600 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01457 1600 1599 1601 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01456 2183 1601 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01455 800 611 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01454 611 2566 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01453 8787 5470 611 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01452 611 1203 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01451 8787 1390 611 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01450 7409 7592 7408 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01449 7408 7593 7410 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01448 8787 8490 7409 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01447 7594 7410 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01446 8787 2159 1985 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01445 1985 3048 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01444 2563 1986 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01443 1985 3717 1986 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01442 1986 2890 1985 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01441 8787 8240 8241 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01440 8241 8488 8243 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01439 8479 8243 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01438 7351 8098 7350 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01437 7350 8020 7352 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01436 8787 8780 7351 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01435 7349 7352 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01434 7778 7852 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01433 7915 8327 7778 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01432 8787 7850 7915 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01431 8055 7915 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01430 5003 5005 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01429 8787 5003 4890 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01428 4890 5007 5005 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01427 5005 5009 4889 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01426 8787 6512 5009 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01425 5007 5009 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01424 8787 4891 5008 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01423 4889 4922 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01422 5002 5007 5003 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01421 4888 5009 5002 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01420 8787 5466 4888 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01419 5466 5002 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01418 8787 5002 5466 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01417 8787 4579 4581 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01416 4830 4581 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01415 8787 4581 4830 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01414 8787 4581 4830 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01413 4830 4581 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01412 8787 4830 4582 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01411 7347 4582 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01410 8787 4582 7347 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01409 8787 4582 7347 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01408 7347 4582 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01407 8787 4830 4831 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01406 8764 4831 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01405 8787 4831 8764 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01404 8787 4831 8764 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01403 8764 4831 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01402 7658 8329 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01401 5428 8103 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01400 4319 7329 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01399 8346 7933 7787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01398 7787 8132 8346 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01397 8787 7932 7787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01396 8751 8752 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01395 8787 8751 8753 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01394 8753 8759 8752 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01393 8752 8760 8757 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01392 8787 8758 8760 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01391 8759 8760 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01390 8787 8754 8756 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01389 8757 8755 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01388 8750 8759 8751 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01387 8749 8760 8750 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01386 8787 8761 8749 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01385 8761 8750 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01384 8787 8750 8761 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01383 2647 2672 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01382 2910 2662 2647 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01381 4957 8553 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01380 3860 7472 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01379 1545 2986 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01378 1978 1567 1545 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01377 6877 7118 6876 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01376 6876 7115 6877 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01375 8787 7514 6876 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01374 7092 6877 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01373 8787 1323 1235 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01372 1235 3110 1324 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01371 1325 1324 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01370 2064 2784 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01369 7535 4577 2064 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01368 8095 8764 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01367 8745 8731 8095 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01366 1861 2508 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01365 1862 3269 1861 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01364 441 560 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01363 556 1128 441 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01362 440 1129 556 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01361 8787 554 440 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01360 1113 556 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01359 8787 1123 439 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01358 439 555 556 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01357 2890 8350 1563 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01356 8787 3158 1565 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01355 1563 1565 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01354 8787 6254 6155 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01353 6155 6255 6256 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01352 6417 6256 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01351 8787 3414 1940 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01350 1942 1952 1936 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01349 1939 2138 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_01348 1936 1935 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01347 1940 1937 1938 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01346 1938 2138 1942 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01345 1942 1939 1941 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01344 2268 1942 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01343 8787 3414 1935 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_01342 1941 1946 1940 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_01341 3873 3874 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01340 6975 3872 3873 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01339 5645 5643 5646 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01338 5646 5644 5645 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01337 8787 6060 5646 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01336 7450 8020 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01335 7579 8247 7450 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01334 7454 8019 7455 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01333 7455 7593 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01332 7453 8490 7454 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01331 7731 8240 7453 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01330 8235 7143 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01329 8787 8430 7145 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01328 6909 7142 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01327 7143 7145 6909 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01326 6907 8430 7143 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01325 8787 7140 6907 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01324 8787 6878 4746 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01323 4746 4758 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01322 4990 4745 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01321 4746 4748 4745 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01320 4745 6077 4746 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01319 4296 4302 4298 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01318 4298 4523 4297 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01317 8787 4295 4296 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01316 5176 4297 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01315 2415 3716 2414 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01314 2414 4750 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01313 2413 6878 2415 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01312 2535 3717 2413 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01311 3157 4984 3156 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01310 3156 3154 3157 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01309 8787 3155 3157 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01308 3157 4988 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01307 7275 7276 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01306 7276 7277 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01305 8787 7880 7276 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01304 7276 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01303 8787 7499 7276 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01302 8787 5033 4908 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01301 4908 7347 5034 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01300 5260 5034 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01299 1013 3531 870 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01298 870 3753 1013 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01297 8787 1154 870 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01296 8787 181 42 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01295 42 374 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01294 1129 173 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01293 42 175 173 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01292 173 378 42 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01291 8787 5989 5991 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01290 5991 6245 5992 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01289 5990 5992 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01288 8787 7184 7028 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01287 7028 7593 7174 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01286 7227 7174 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01285 8787 7315 6206 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01284 6206 6541 6369 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01283 6374 6369 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01282 8787 786 784 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01281 784 793 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01280 2302 785 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01279 784 1149 785 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01278 785 783 784 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_01277 6696 6693 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01276 8787 6696 6562 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01275 6562 6695 6693 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01274 6693 6698 6561 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01273 8787 8596 6698 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01272 6695 6698 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01271 8787 6609 6697 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01270 6561 6626 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01269 6692 6695 6696 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01268 6560 6698 6692 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01267 8787 6691 6560 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01266 6691 6692 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01265 8787 6692 6691 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01264 139 142 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01263 8787 139 32 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01262 32 143 142 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01261 142 145 34 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01260 8787 1516 145 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01259 143 145 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01258 8787 33 144 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01257 34 140 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01256 137 143 139 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01255 31 145 137 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01254 8787 764 31 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01253 764 137 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01252 8787 137 764 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01251 836 8350 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01250 8787 3158 836 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01249 5136 5790 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01248 8787 5790 5138 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01247 5139 5135 5136 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01246 5134 5138 5139 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01245 8787 5466 5134 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01244 5135 5466 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01243 7640 8572 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01242 7639 7643 7640 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01241 8787 7641 7639 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01240 93 97 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01239 8787 93 16 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01238 16 99 97 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01237 97 101 17 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01236 8787 1302 101 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01235 99 101 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01234 8787 18 100 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01233 17 95 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01232 94 99 93 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01231 15 101 94 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01230 8787 542 15 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01229 542 94 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01228 8787 94 542 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01227 3772 3771 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01226 8787 3773 3772 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01225 3772 4152 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01224 8787 3977 3772 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01223 3265 2505 2398 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01222 2398 2504 3265 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01221 8787 7877 2398 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01220 8787 7116 7541 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01219 7541 7111 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01218 8787 7112 7541 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01217 5419 5420 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01216 8787 5419 5310 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01215 5310 5418 5420 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01214 5420 5424 5311 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01213 8787 5835 5424 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01212 5418 5424 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01211 8787 5344 5422 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01210 5311 5361 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01209 5416 5418 5419 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01208 5309 5424 5416 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01207 8787 5415 5309 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01206 5415 5416 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01205 8787 5416 5415 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01204 3187 3400 3188 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01203 3188 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01202 3398 3429 3187 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01201 3601 3767 3600 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01200 3600 6282 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01199 4999 5562 3601 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01198 4419 4536 4420 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01197 4420 4539 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01196 4418 6040 4419 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01195 4720 6021 4418 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01194 5383 5114 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01193 8787 6934 5115 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01192 5113 5112 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01191 5114 5115 5113 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01190 5111 6934 5114 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01189 8787 6290 5111 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01188 6521 7171 6520 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01187 6520 7170 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01186 6760 6765 6521 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01185 4911 5048 4912 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01184 4912 5043 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01183 5041 5042 4911 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01182 3314 1015 871 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01181 871 1016 3314 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01180 8787 2151 871 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01179 3497 3494 3496 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01178 3496 3498 3495 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01177 8787 3493 3497 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01176 4321 3495 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01175 7798 8135 8175 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01174 8787 8135 7961 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01173 7799 8383 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01172 8175 7961 7799 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01171 8787 8566 7798 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01170 8787 4538 4287 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01169 4287 4712 4288 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01168 4286 4288 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01167 4142 4137 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01166 8787 5036 4137 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01165 4137 5790 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01164 8787 8731 4137 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01163 3388 3271 3099 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01162 3099 3262 3388 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01161 8787 3261 3099 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01160 8787 807 44 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01159 44 2976 176 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01158 382 176 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01157 7782 8135 8202 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01156 8787 8135 7927 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01155 7783 7937 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01154 8202 7927 7783 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01153 8787 7928 7782 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01152 7386 8246 7385 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01151 7385 8098 7387 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01150 8787 8237 7386 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01149 8227 7387 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01148 7374 8236 7376 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01147 7376 8020 7375 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01146 8787 8247 7374 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01145 7373 7375 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01144 526 528 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01143 8787 526 428 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01142 428 530 528 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01141 528 531 429 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01140 8787 1302 531 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01139 530 531 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01138 8787 468 529 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01137 429 488 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01136 524 530 526 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01135 427 531 524 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01134 8787 726 427 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01133 726 524 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01132 8787 524 726 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01131 899 4300 900 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01130 900 2764 1041 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01129 8787 4139 899 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01128 1202 1041 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01127 1467 1729 1468 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01126 1468 1902 1467 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01125 8787 1723 1468 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01124 1898 1467 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01123 4040 7228 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01122 5162 6708 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01121 3604 3767 3605 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01120 3605 4109 3752 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01119 8787 3956 3604 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01118 3912 3752 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01117 8117 8329 8066 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01116 8787 8065 8067 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01115 8066 8067 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01114 8085 8087 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01113 8787 8085 8086 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01112 8086 8088 8087 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01111 8087 8150 8148 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01110 8787 8674 8150 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01109 8088 8150 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01108 8787 8151 8152 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01107 8148 8147 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01106 8145 8088 8085 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01105 8084 8150 8145 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01104 8787 8372 8084 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01103 8372 8145 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01102 8787 8145 8372 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01101 952 955 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01100 8787 952 852 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01099 852 956 955 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01098 955 958 854 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01097 8787 1516 958 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01096 956 958 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01095 8787 853 957 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01094 854 907 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01093 951 956 952 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01092 851 958 951 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01091 8787 959 851 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01090 959 951 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01089 8787 951 959 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01088 4289 4715 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01087 7905 8761 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01086 5042 5270 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01085 3610 3936 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01084 3759 3931 3610 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01083 4263 4498 4262 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01082 4262 4485 4263 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01081 8787 4944 4262 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01080 4479 4263 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01079 1793 1381 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01078 8787 1382 1793 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01077 1793 1590 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01076 8787 1798 1793 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01075 474 6718 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01074 1016 5563 474 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01073 5829 5831 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01072 8787 5829 5722 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01071 5722 5836 5831 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01070 5831 5837 5721 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01069 8787 5835 5837 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01068 5836 5837 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01067 8787 5723 5834 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01066 5721 5775 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01065 5828 5836 5829 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01064 5720 5837 5828 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01063 8787 5826 5720 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01062 5826 5828 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01061 8787 5828 5826 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01060 2764 5470 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01059 8787 1203 2764 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01058 2764 1390 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01057 8787 2566 2764 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_01056 8785 8781 8783 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01055 8783 8782 8785 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01054 8787 8780 8783 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01053 5347 5469 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01052 5888 6072 5347 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01051 6617 6950 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01050 6660 6766 6617 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01049 8069 8327 7784 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01048 7784 7930 8069 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01047 8787 7929 7784 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01046 3430 3956 3432 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01045 3432 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01044 3431 4300 3430 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01043 3429 8553 3431 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01042 7735 6733 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01041 8787 8430 6734 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01040 6581 6735 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01039 6733 6734 6581 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01038 6580 8430 6733 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01037 8787 6908 6580 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01036 7991 7725 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01035 8787 8423 7726 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01034 7724 7723 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01033 7725 7726 7724 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01032 7722 8423 7725 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01031 8787 7987 7722 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01030 7707 7549 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01029 8787 8423 7551 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01028 7433 7718 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01027 7549 7551 7433 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01026 7432 8423 7549 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01025 8787 7716 7432 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01024 8787 5246 5248 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01023 5248 5484 5247 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01022 5244 5247 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01021 4408 7315 4409 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01020 4409 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01019 4523 4522 4408 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01018 3190 3258 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01017 3405 3670 3190 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01016 8787 3257 3405 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01015 3624 3960 3625 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01014 3625 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01013 3623 3964 3624 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01012 3775 5471 3623 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01011 8696 8418 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01010 8787 8423 8420 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01009 8190 8417 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01008 8418 8420 8190 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01007 8188 8423 8418 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01006 8787 8690 8188 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01005 2061 2153 2062 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01004 2062 2155 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01003 2060 2307 2061 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01002 3677 2154 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01001 2154 2059 2060 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01000 7331 7333 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00999 8787 7347 7334 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00998 7332 7575 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00997 7333 7334 7332 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00996 7330 7347 7333 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00995 8787 7329 7330 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00994 2057 2305 2058 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00993 2058 6878 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00992 2056 4530 2057 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00991 3678 2152 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00990 2152 2055 2056 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00989 3821 3822 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00988 8787 3822 3823 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00987 5112 3819 3821 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00986 3820 3823 5112 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00985 8787 3826 3820 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00984 3819 3826 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00983 1100 1463 1099 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00982 1099 1462 1100 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00981 8787 2723 1099 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00980 3840 1462 1464 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00979 1464 1463 3840 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00978 8787 7877 1464 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00977 5805 5809 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00976 5809 5810 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00975 8787 7880 5809 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00974 5809 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00973 8787 7877 5809 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00972 7076 7079 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00971 6993 7535 7079 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00970 7079 7077 6992 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00969 6992 7081 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00968 8787 7536 6993 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00967 6993 7533 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00966 7016 7358 7015 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00965 7015 7362 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00964 7014 7167 7016 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00963 7573 7356 7014 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00962 8482 8776 8305 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00961 8305 8479 8482 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00960 8787 8480 8305 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00959 6841 7065 6842 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00958 6842 7066 6841 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00957 8787 8065 6842 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00956 8787 1140 1133 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00955 1133 5214 1134 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00954 1339 1134 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00953 8787 5280 4022 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00952 4022 5508 4151 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00951 4152 4151 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00950 8348 7879 7425 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00949 7425 8132 8348 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00948 8787 7532 7425 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00947 8787 5563 39 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00946 39 4536 159 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00945 602 159 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00944 7390 8483 7389 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00943 7389 8098 7388 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00942 8787 8237 7390 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00941 7391 7388 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00940 7242 7245 7241 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00939 7241 7480 7242 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00938 8787 7240 7241 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00937 2137 2274 1943 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00936 1943 2273 2137 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00935 8787 2260 1943 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00934 1108 1114 1109 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00933 1109 1113 1108 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00932 8787 2260 1109 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00931 1476 1108 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00930 5771 5922 5772 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00929 5772 6134 5921 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00928 8787 6136 5771 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00927 5920 5921 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00926 2022 2021 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00925 8787 2022 1875 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00924 1875 2026 2021 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00923 2021 2029 2024 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00922 8787 2028 2029 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00921 2026 2029 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00920 8787 2025 2027 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00919 2024 2023 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00918 2020 2026 2022 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00917 1874 2029 2020 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00916 8787 2189 1874 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00915 2189 2020 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00914 8787 2020 2189 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00913 3643 3641 3557 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00912 3557 3826 3643 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00911 8787 3827 3557 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00910 3814 3643 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00909 776 994 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00908 1135 775 776 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00907 8787 1123 773 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00906 773 993 1135 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00905 8787 992 774 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00904 774 1129 1135 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00903 278 532 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00902 279 1128 278 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00901 277 1129 279 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00900 8787 276 277 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00899 1463 279 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00898 8787 1123 275 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00897 275 274 279 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00896 5900 5903 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00895 8787 5900 5750 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00894 5750 5905 5903 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00893 5903 5906 5752 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00892 8787 6361 5906 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00891 5905 5906 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00890 8787 5751 5904 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00889 5752 5778 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00888 5898 5905 5900 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00887 5749 5906 5898 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00886 8787 6316 5749 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00885 6316 5898 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00884 8787 5898 6316 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00883 885 3960 886 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00882 886 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00881 884 5013 885 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00880 1034 1035 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00879 1035 883 884 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00878 8787 7120 7693 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00877 7693 7121 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00876 8787 7124 7693 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00875 6225 6229 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00874 8787 6225 6140 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00873 6140 6230 6229 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00872 6229 6233 6142 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00871 8787 6232 6233 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00870 6230 6233 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00869 8787 6141 6231 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00868 6142 6217 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00867 6226 6230 6225 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00866 6139 6233 6226 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00865 8787 6223 6139 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00864 6223 6226 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00863 8787 6226 6223 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00862 3564 3657 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00861 5785 3658 3564 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00860 3563 3654 5785 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00859 8787 3832 3563 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00858 3563 3655 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00857 2691 2942 2692 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00856 2692 3479 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00855 3655 2940 2691 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00854 2829 3471 2830 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00853 2830 3478 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00852 2947 3885 2829 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00851 4145 4157 4020 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00850 4020 6672 4145 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00849 8787 4144 4020 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00848 4143 4145 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00847 6899 7118 6898 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00846 6898 7115 6899 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00845 8787 8661 6898 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00844 7120 6899 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00843 7465 8488 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00842 7589 7759 7465 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00841 7464 8479 7589 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00840 8787 7588 7464 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00839 7464 8027 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00838 5708 5958 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00837 8787 5958 5780 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00836 8787 6223 5707 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00835 5781 5779 5708 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00834 5707 5780 5781 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00833 5789 5781 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00832 8787 5781 5789 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00831 5779 6223 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00830 4651 4652 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00829 8787 4651 4653 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00828 4653 4658 4652 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00827 4652 4659 4656 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00826 8787 6232 4659 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00825 4658 4659 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00824 8787 4654 4657 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00823 4656 4655 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00822 4650 4658 4651 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00821 4649 4659 4650 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00820 8787 5851 4649 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00819 5851 4650 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00818 8787 4650 5851 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00817 2087 2171 2086 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00816 2086 2178 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00815 2776 2170 2087 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00814 7429 7541 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00813 8688 7540 7429 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00812 7461 8235 7460 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00811 7460 8097 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00810 7757 8215 7461 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00809 4660 4664 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00808 8787 6934 4665 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00807 4663 4662 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00806 4664 4665 4663 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00805 4661 6934 4664 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00804 8787 5851 4661 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00803 8787 6432 4858 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00802 4858 4966 4967 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00801 4965 4967 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00800 8787 5870 4325 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00799 4325 4328 4326 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00798 4324 4326 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00797 8394 2301 2303 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00796 2303 2302 8394 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00795 8787 8065 2303 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00794 8787 4978 4721 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00793 4721 4720 4722 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00792 4974 4722 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00791 7641 6843 6845 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00790 6845 6860 7641 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00789 8787 6844 6845 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00788 7249 7251 7248 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00787 7248 7481 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00786 7247 7252 7249 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00785 7637 7246 7247 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00784 3046 5013 3045 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00783 3045 6029 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00782 3044 6021 3046 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00781 3100 3101 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00780 3101 3043 3044 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00779 1965 7536 1964 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00778 1964 7533 1965 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00777 8787 2334 1964 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00776 1967 1965 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00775 6610 6701 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00774 6632 8135 6610 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00773 3160 3159 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00772 3159 3050 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00771 8787 8731 3159 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00770 3048 1774 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00769 1774 1695 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00768 8787 3158 1774 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00767 6525 6673 6524 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00766 6524 6954 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00765 6765 8490 6525 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00764 8787 8778 8245 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00763 8245 8248 8244 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00762 8242 8244 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00761 6986 7252 6987 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00760 6987 7251 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00759 6985 7065 6986 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00758 7480 7067 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00757 7067 6984 6985 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00756 8254 8323 8253 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00755 8253 8325 8322 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00754 8787 8326 8254 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00753 8321 8322 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00752 6615 6726 6614 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00751 6614 6728 6725 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00750 8787 6727 6615 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00749 7542 6725 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00748 6989 7071 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00747 7077 8135 6989 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00746 5281 8490 5282 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00745 5282 6677 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00744 5278 5280 5281 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00743 5279 6378 5278 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00742 7888 7959 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00741 7959 7879 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00740 8787 7880 7959 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00739 7959 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00738 8787 7877 7959 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00737 8787 6946 6949 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00736 6949 7381 6948 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00735 6947 6948 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00734 5432 7307 5314 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00733 5314 7308 5432 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00732 8787 8427 5314 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00731 8787 2315 2313 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00730 2313 6878 2314 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00729 2727 2314 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00728 8787 3776 3554 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00727 3554 3553 3555 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00726 3552 3555 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00725 8787 5920 5337 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00724 5337 6118 5511 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00723 5510 5511 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00722 6962 8222 6963 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00721 6963 8246 6962 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00720 8787 8780 6963 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00719 6961 6962 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00718 7649 7928 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00717 7648 8135 7649 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00716 8787 5411 5154 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00715 5154 5611 5155 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00714 5153 5155 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00713 2924 3095 2818 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00712 2818 3100 2924 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00711 8787 3673 2818 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00710 2923 2924 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00709 7035 8235 7034 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00708 7034 8097 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00707 7033 8246 7035 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00706 7178 7179 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00705 7179 7032 7033 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00704 2726 3885 2725 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00703 2725 3471 2724 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00702 8787 4999 2726 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00701 2723 2724 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00700 2460 2981 2461 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00699 2461 3012 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00698 2459 3335 2460 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00697 2588 2590 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00696 2590 2465 2459 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00695 3523 4109 3522 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00694 3522 6037 3524 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00693 8787 3753 3523 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00692 3944 3524 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00691 5477 5478 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00690 8787 5477 5327 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00689 5327 5476 5478 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00688 5478 5482 5328 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00687 8787 6512 5482 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00686 5476 5482 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00685 8787 5352 5481 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00684 5328 5364 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00683 5474 5476 5477 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00682 5326 5482 5474 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00681 8787 5676 5326 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00680 5676 5474 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00679 8787 5474 5676 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00678 6121 6543 6124 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00677 6124 6123 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00676 6122 6372 6121 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00675 6118 6120 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00674 6120 6119 6122 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00673 2357 2584 2358 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00672 2358 2359 2360 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00671 8787 3324 2357 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00670 2592 2360 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00669 2185 1591 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00668 8787 1592 2185 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00667 6288 5851 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00666 6859 6027 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00665 4928 5790 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00664 2646 2644 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00663 2906 2645 2646 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00662 4502 5440 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00661 4929 5466 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00660 2875 2962 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00659 3307 2963 2875 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00658 2440 2570 2439 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00657 2439 2569 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00656 2775 2756 2440 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00655 7104 7127 6999 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00654 6999 7126 7104 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00653 8787 7718 6999 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00652 7102 7104 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00651 4880 4999 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00650 4997 6077 4880 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00649 4748 4747 4749 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00648 4749 4755 4748 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00647 8787 5188 4749 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00646 6002 6272 6001 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00645 6001 6889 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00644 6255 6000 6002 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00643 8787 1308 1102 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00642 1102 3854 1101 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00641 1309 1101 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00640 5556 5890 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00639 5555 5554 5556 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00638 869 1011 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00637 1147 1009 869 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00636 868 2542 1147 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00635 8787 3531 868 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00634 868 3753 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00633 8787 3102 2650 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00632 2650 3092 2649 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00631 2648 2649 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00630 2067 6285 2068 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00629 2068 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00628 2315 3767 2067 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00627 5346 5469 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00626 5554 5466 5346 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00625 8787 6878 6154 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00624 6154 6252 6253 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00623 6408 6253 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00622 8787 3414 1238 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00621 1332 1325 1236 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00620 1327 1755 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_00619 1236 1328 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00618 1238 1333 1237 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00617 1237 1755 1332 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00616 1332 1327 1239 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00615 1923 1332 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00614 8787 3414 1328 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_00613 1239 1744 1238 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00612 3090 3095 3091 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00611 3091 3100 3090 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00610 8787 3673 3091 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00609 1541 1538 1540 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00608 1540 4795 1542 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00607 8787 1539 1541 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00606 1537 1542 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00605 2966 2755 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00604 2755 2753 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00603 8787 2754 2755 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00602 8450 8187 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00601 8787 8430 8189 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00600 8186 8185 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00599 8187 8189 8186 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00598 8184 8430 8187 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00597 8787 8191 8184 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00596 6633 6864 6611 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00595 8787 8135 6705 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00594 6611 6705 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00593 6323 6325 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00592 8787 7347 6328 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00591 6188 7164 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00590 6325 6328 6188 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00589 6187 7347 6325 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00588 8787 6324 6187 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00587 2669 2682 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00586 2670 2930 2669 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00585 8787 3257 2670 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00584 2856 3956 2857 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00583 2857 6043 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00582 2855 6284 2856 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00581 2934 2935 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00580 2935 2854 2855 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00579 8483 8193 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00578 8787 8430 8197 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00577 8195 8417 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00576 8193 8197 8195 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00575 8192 8430 8193 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00574 8787 8690 8192 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00573 6420 6852 6419 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00572 8787 8135 6421 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00571 6419 6421 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00570 8302 8475 8303 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00569 8303 8769 8476 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00568 8787 8482 8302 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00567 8474 8476 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00566 3387 3832 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00565 3390 3828 3387 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00564 3386 3827 3390 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00563 8787 3825 3386 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00562 3386 3826 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00561 8787 4139 4016 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00560 4016 4142 4141 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00559 4140 4141 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00558 4553 3158 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00557 5231 6758 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00556 8625 8128 7673 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00555 7673 8132 8625 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00554 8787 8127 7673 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00553 386 382 387 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00552 387 388 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00551 384 614 386 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00550 1128 385 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00549 385 383 384 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00548 8445 8717 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00547 5365 5565 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00546 4759 4758 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00545 8787 3324 2454 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00544 2454 2584 2585 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00543 2589 2585 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00542 8787 3717 2758 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_00541 2758 3048 8787 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_00540 2756 2757 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00539 2758 4530 2757 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_00538 2757 2890 2758 8787 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_00537 6861 6859 6862 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00536 6862 6860 6861 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00535 8787 6858 6862 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00534 6812 6814 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00533 8787 6812 6813 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00532 6813 6815 6814 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00531 6814 6869 6868 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00530 8787 8674 6869 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00529 6815 6869 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00528 8787 6870 6871 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00527 6868 6867 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00526 6863 6815 6812 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00525 6811 6869 6863 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00524 8787 6864 6811 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00523 6864 6863 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00522 8787 6863 6864 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00521 3954 6029 3955 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00520 3955 5046 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00519 3953 5471 3954 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00518 3950 3952 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00517 3952 3951 3953 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00516 4135 5790 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00515 8787 8731 4135 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00514 1152 7536 1153 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00513 1153 7533 1152 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00512 8787 2161 1153 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00511 1151 1152 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00510 68 71 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00509 8787 68 6 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00508 6 73 71 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00507 71 74 8 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00506 8787 1302 74 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00505 73 74 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00504 8787 7 72 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00503 8 69 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00502 67 73 68 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00501 5 74 67 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00500 8787 276 5 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00499 276 67 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00498 8787 67 276 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00497 8361 7681 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00496 7681 7679 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00495 8787 7680 7681 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00494 8787 6820 7545 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00493 7545 6821 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00492 8787 6819 7545 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00491 7413 8553 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00490 7636 7643 7413 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00489 8787 7485 7636 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00488 6050 6055 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00487 8787 6050 6051 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00486 6051 6057 6055 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00485 6055 6059 6056 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00484 8787 6512 6059 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00483 6057 6059 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00482 8787 6053 6058 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00481 6056 6054 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00480 6048 6057 6050 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00479 6049 6059 6048 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00478 8787 6062 6049 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00477 6062 6048 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00476 8787 6048 6062 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00475 5452 5455 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00474 8787 5452 5319 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00473 5319 5453 5455 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00472 5455 5456 5320 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00471 8787 6512 5456 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00470 5453 5456 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00469 8787 5345 5457 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00468 5320 5362 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00467 5450 5453 5452 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00466 5318 5456 5450 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00465 8787 6060 5318 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00464 6060 5450 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00463 8787 5450 6060 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00462 2243 2664 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00461 2244 3090 2243 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00460 8787 3257 2244 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00459 2476 2244 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00458 3089 3429 3088 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00457 3088 3400 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00456 3258 3254 3089 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00455 4415 4532 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00454 4534 4533 4415 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00453 8787 6735 4534 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00452 4966 4534 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00451 7694 7693 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00450 8716 7888 7694 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00449 1498 1500 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00448 8787 2263 1502 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00447 1501 3254 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00446 1500 1502 1501 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00445 1499 2263 1500 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00444 8787 3673 1499 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00443 1889 2127 1888 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00442 1888 2255 1887 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00441 8787 3657 1889 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00440 1886 1887 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00439 8787 7291 7290 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00438 7290 7288 7289 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00437 8127 7289 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00436 2766 3960 2765 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00435 2765 2764 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00434 2763 3964 2766 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00433 6428 6431 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00432 6429 7535 6431 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00431 6431 6632 6430 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00430 6430 6633 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00429 8787 7536 6429 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00428 6429 7533 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00427 7820 8235 7821 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00426 7821 8020 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00425 7906 8237 7820 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00424 8787 5637 5640 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00423 5640 5638 5639 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00422 5662 5639 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00421 6213 8240 6214 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00420 6214 8478 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00419 6376 8480 6213 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00418 7572 7574 7440 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00417 7440 7731 7572 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00416 8787 7570 7440 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00415 7823 8483 7822 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00414 7822 8236 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00413 7907 8247 7823 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00412 7760 7757 7759 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00411 7759 7907 7760 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00410 8787 7758 7760 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00409 7760 7906 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00408 4872 4985 4873 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00407 4873 4987 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00406 4871 4984 4872 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00405 5438 4986 4871 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00404 2031 2105 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00403 8787 2105 2106 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00402 5978 2102 2031 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00401 2030 2106 5978 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00400 8787 2103 2030 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00399 2102 2103 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00398 2780 6718 2779 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00397 2779 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00396 2778 3956 2780 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00395 3006 6284 2778 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00394 3905 6873 3904 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00393 3904 3903 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00392 3902 5010 3905 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00391 7881 4999 3902 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00390 7747 8236 7745 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00389 7745 8020 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00388 7746 8247 7747 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00387 8787 3278 1096 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00386 1095 1096 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00385 8787 1096 1095 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00384 8787 1096 1095 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00383 1095 1096 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00382 8787 3278 1301 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00381 1300 1301 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00380 8787 1301 1300 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00379 8787 1301 1300 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00378 1300 1301 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00377 8787 3278 1303 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00376 1302 1303 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00375 8787 1303 1302 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00374 8787 1303 1302 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00373 1302 1303 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00372 3958 4109 3959 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00371 3959 3960 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00370 3957 4577 3958 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00369 4144 3956 3957 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00368 5161 5163 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00367 5163 5162 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00366 8787 7273 5163 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00365 5163 7881 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00364 8787 7877 5163 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00363 8787 8010 8009 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00362 8207 8009 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00361 8787 8009 8207 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00360 8787 8009 8207 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00359 8207 8009 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00358 8787 8207 8206 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00357 8215 8206 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00356 8787 8206 8215 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00355 8787 8206 8215 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00354 8215 8206 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00353 8787 8207 8013 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00352 8237 8013 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00351 8787 8013 8237 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00350 8787 8013 8237 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00349 8237 8013 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00348 8787 8207 8014 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00347 8247 8014 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00346 8787 8014 8247 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00345 8787 8014 8247 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00344 8247 8014 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00343 8787 8207 8208 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00342 8780 8208 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00341 8787 8208 8780 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00340 8787 8208 8780 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00339 8780 8208 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00338 1896 1897 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00337 8787 1897 1894 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00336 4662 1893 1896 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00335 1895 1894 4662 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00334 8787 1911 1895 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00333 1893 1911 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00332 3324 3325 3236 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00331 3236 6365 3324 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00330 8787 3333 3236 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00329 4392 5466 4391 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00328 4391 4943 4489 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00327 8787 5415 4392 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00326 4488 4489 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00325 8787 198 197 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00324 416 197 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00323 8787 197 416 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00322 8787 197 416 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00321 416 197 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00320 8787 416 411 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00319 5465 411 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00318 8787 411 5465 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00317 8787 411 5465 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00316 5465 411 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00315 8787 416 417 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00314 5562 417 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00313 8787 417 5562 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00312 8787 417 5562 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00311 5562 417 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00310 8787 3278 1122 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00309 1121 1122 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00308 8787 1122 1121 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00307 8787 1122 1121 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00306 1121 1122 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00305 8787 3278 1336 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00304 1335 1336 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00303 8787 1336 1335 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00302 8787 1336 1335 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00301 1335 1336 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00300 8787 3278 1337 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00299 1516 1337 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00298 8787 1337 1516 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00297 8787 1337 1516 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00296 1516 1337 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00295 8787 3278 3077 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00294 3076 3077 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00293 8787 3077 3076 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00292 8787 3077 3076 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00291 3076 3077 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00290 8787 3278 3252 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00289 3251 3252 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00288 8787 3252 3251 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00287 8787 3252 3251 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00286 3251 3252 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00285 8787 3278 3253 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00284 4057 3253 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00283 8787 3253 4057 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00282 8787 3253 4057 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00281 4057 3253 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00280 8787 3278 3114 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00279 3113 3114 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00278 8787 3114 3113 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00277 8787 3114 3113 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00276 3113 3114 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00275 1097 1462 1098 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00274 1098 1463 1097 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00273 8787 2260 1098 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00272 2121 1097 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00271 2019 4139 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00270 2795 2017 2019 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00269 2018 3960 2795 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00268 8787 2015 2018 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00267 2018 2016 8787 8787 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00266 2706 5440 2705 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00265 8787 8627 2708 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00264 2705 2708 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00263 3878 3875 3877 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00262 3877 3880 3876 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00261 8787 3881 3878 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00260 3874 3876 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00259 2436 2769 2435 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00258 2435 2564 2565 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00257 8787 2563 2436 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00256 2972 2565 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00255 4876 5010 4877 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00254 4877 6873 4992 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00253 8787 4999 4876 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00252 6246 4992 8787 8787 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00251 8787 3278 3277 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00250 3276 3277 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00249 8787 3277 3276 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00248 8787 3277 3276 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00247 3276 3277 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00246 8787 3278 3279 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00245 3705 3279 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00244 8787 3279 3705 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00243 8787 3279 3705 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00242 3705 3279 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00241 8787 3330 1167 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00240 1166 1167 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00239 8787 1167 1166 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00238 8787 1167 1166 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00237 1166 1167 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00236 8787 3330 1366 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00235 1365 1366 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00234 8787 1366 1365 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00233 8787 1366 1365 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00232 1365 1366 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00231 8787 3330 1368 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00230 1367 1368 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00229 8787 1368 1367 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00228 8787 1368 1367 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00227 1367 1368 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00226 8787 3330 1200 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00225 1199 1200 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00224 8787 1200 1199 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00223 8787 1200 1199 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00222 1199 1200 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00221 8787 3330 1387 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00220 1386 1387 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00219 8787 1387 1386 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00218 8787 1387 1386 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00217 1386 1387 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00216 8787 3330 1388 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00215 2028 1388 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00214 8787 1388 2028 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00213 8787 1388 2028 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00212 2028 1388 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00211 592 594 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00210 8787 592 453 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00209 453 597 594 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00208 594 598 454 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00207 8787 1367 598 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00206 597 598 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00205 8787 471 596 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00204 454 491 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00203 591 597 592 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00202 452 598 591 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00201 8787 994 452 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00200 994 591 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00199 8787 591 994 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00198 1259 4109 1260 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00197 1260 6037 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00196 1258 4577 1259 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00195 1564 1370 8787 8787 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00194 1370 1275 1258 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00193 4847 4937 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00192 8787 4937 4938 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00191 4935 4933 4847 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00190 4846 4938 4935 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00189 8787 4934 4846 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00188 4933 4934 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00187 8787 3338 2596 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00186 2596 3015 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00185 8787 2593 2596 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00184 2179 1602 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00183 8787 1596 2179 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00182 8787 6072 6073 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00181 6073 6352 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00180 8787 6316 6073 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00179 8787 3330 3149 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00178 3148 3149 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00177 8787 3149 3148 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00176 8787 3149 3148 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00175 3148 3149 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00174 8787 3330 3303 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00173 3302 3303 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00172 8787 3303 3302 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00171 8787 3303 3302 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00170 3302 3303 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00169 8787 3330 3304 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00168 4121 3304 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00167 8787 3304 4121 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00166 8787 3304 4121 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00165 4121 3304 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00164 8787 3330 3173 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00163 3172 3173 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00162 8787 3173 3172 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00161 8787 3173 3172 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00160 3172 3173 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00159 8787 3330 3328 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00158 3327 3328 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00157 8787 3328 3327 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00156 8787 3328 3327 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00155 3327 3328 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00154 8787 3330 3331 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00153 3329 3331 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00152 8787 3331 3329 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00151 8787 3331 3329 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00150 3329 3331 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00149 8664 8669 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00148 8787 8664 8668 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00147 8668 8672 8669 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00146 8669 8675 8667 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00145 8787 8674 8675 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00144 8672 8675 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00143 8787 8671 8673 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00142 8667 8666 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00141 8663 8672 8664 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00140 8662 8675 8663 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00139 8787 8661 8662 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00138 8661 8663 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00137 8787 8663 8661 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00136 7021 8030 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00135 7167 7353 7021 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00134 6827 8030 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00133 7358 6940 6827 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00132 4342 5036 4012 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00131 4012 6077 4342 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00130 8787 6307 4012 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00129 8787 7684 5387 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00128 5386 5387 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00127 8787 5387 5386 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00126 8787 5387 5386 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00125 5386 5387 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00124 1956 1961 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00123 8787 2949 1963 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00122 1960 1959 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00121 1961 1963 1960 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00120 1957 2949 1961 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00119 8787 6324 1957 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00118 2783 2782 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_00117 8787 2787 2783 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_00116 2783 3001 8787 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_00115 8787 2781 2783 8787 sg13_lv_nmos L=0.13U W=0.84U AS=0.2016P AD=0.2016P PS=2.17U PD=2.17U 
Mtr_00114 1249 6285 1250 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00113 1250 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00112 3717 3964 1249 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00111 3226 6040 3225 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00110 3225 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00109 4530 3964 3226 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00108 6201 8487 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00107 6364 8227 6201 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00106 4437 5031 8787 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00105 4565 4754 4437 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00104 7305 7307 7306 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00103 7306 7308 7305 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00102 8787 8417 7306 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00101 8787 7684 5591 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00100 5590 5591 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00099 8787 5591 5590 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00098 8787 5591 5590 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00097 5590 5591 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00096 8787 7684 5592 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00095 6232 5592 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00094 8787 5592 6232 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00093 8787 5592 6232 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00092 6232 5592 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00091 8787 7684 5431 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00090 5430 5431 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00089 8787 5431 5430 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00088 8787 5431 5430 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00087 5430 5431 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00086 8787 7684 5629 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00085 5628 5629 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00084 8787 5629 5628 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00083 8787 5629 5628 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00082 5628 5629 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00081 7664 7667 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00080 8787 7664 7665 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00079 7665 7671 7667 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00078 7667 7672 7666 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00077 8787 8674 7672 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00076 7671 7672 8787 8787 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00075 8787 7668 7670 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00074 7666 7663 8787 8787 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00073 7662 7671 7664 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00072 7661 7672 7662 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00071 8787 7660 7661 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00070 7660 7662 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00069 8787 7662 7660 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00068 8787 3414 1615 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00067 1718 1922 1612 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00066 1715 1716 8787 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_00065 1612 1711 8787 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00064 1615 1712 1613 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00063 1613 1716 1718 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00062 1718 1715 1614 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00061 1710 1718 8787 8787 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00060 8787 3414 1711 8787 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_00059 1614 1717 1615 8787 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00058 8787 7684 5630 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00057 5835 5630 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00056 8787 5630 5835 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00055 8787 5630 5835 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00054 5835 5630 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00053 8787 7684 7489 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00052 7488 7489 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00051 8787 7489 7488 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00050 8787 7489 7488 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00049 7488 7489 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00048 8787 7684 7646 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00047 7645 7646 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00046 8787 7646 7645 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00045 8787 7646 7645 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00044 7645 7646 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00043 8787 7684 7647 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00042 8596 7647 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00041 8787 7647 8596 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00040 8787 7647 8596 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00039 8596 7647 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00038 2668 2682 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00037 2667 2930 2668 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00036 8787 3257 2667 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00035 2666 2667 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00034 8787 6878 6435 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00033 6435 6711 6436 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00032 6714 6436 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00031 1634 5013 1635 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00030 1635 4536 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00029 3716 4300 1634 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00028 8222 7147 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00027 8787 8430 7149 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00026 6913 7326 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00025 7147 7149 6913 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00024 6912 8430 7147 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00023 8787 7553 6912 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00022 3927 3756 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00021 8787 4747 3758 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00020 3609 3755 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00019 3756 3758 3609 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00018 3608 4747 3756 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00017 8787 4792 3608 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00016 6648 6738 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00015 8787 6934 6740 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00014 6585 7151 8787 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00013 6738 6740 6585 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00012 6584 6934 6738 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00011 8787 6739 6584 8787 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00010 8028 8486 7825 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00009 7825 8029 8028 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00008 8787 8030 7825 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00007 7913 8028 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00006 8787 3717 2316 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00005 2316 2315 2317 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00004 2321 2317 8787 8787 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00003 7065 5162 4860 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00002 4860 5169 7065 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00001 8787 4973 4860 8787 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
.ends arlet6502_cts_r_transistors_ihp

