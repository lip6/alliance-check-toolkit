* nand4_x0
* nand4_x0
.subckt nand4_x0 vdd vss nq i0 i1 i2 i3
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net0 i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos _net1 i2 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi3_nmos _net2 i3 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi3_pmos nq i3 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nand4_x0
