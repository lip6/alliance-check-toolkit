-- no model for nor2_x0
