* fill_w2
* fill_w2
.subckt fill_w2 vdd vss

.ends fill_w2
