* Spice description of ts_x4
* Spice driver version -1161363685
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:42

* INTERF cmd i q vdd vss 


.subckt ts_x4 4 3 8 1 7 
* NET 1 = vdd
* NET 3 = i
* NET 4 = cmd
* NET 5 = 4
* NET 7 = vss
* NET 8 = q
Mtr_00012 8 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 1 2 8 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 5 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00009 1 4 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00008 2 5 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 2 3 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 6 3 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00005 8 6 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 7 6 8 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 5 4 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 7 5 6 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 2 4 6 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C8 1 7 3.35605e-15
C7 2 7 2.84697e-15
C6 3 7 1.73025e-15
C5 4 7 3.52478e-15
C4 5 7 1.82426e-15
C3 6 7 2.37576e-15
C2 7 7 2.94905e-15
C1 8 7 2.15173e-15
.ends ts_x4

