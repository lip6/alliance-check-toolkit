* Spice description of nmx2_x1
* Spice driver version -964804837
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:57

* INTERF cmd i0 i1 nq vdd vss 


.subckt nmx2_x1 9 8 4 6 3 10 
* NET 3 = vdd
* NET 4 = i1
* NET 6 = nq
* NET 8 = i0
* NET 9 = cmd
* NET 10 = vss
* NET 11 = q
Mtr_00010 3 4 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 6 9 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 2 8 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 3 9 11 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 1 11 6 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 10 4 5 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 6 11 7 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 7 8 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 10 9 11 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 5 9 6 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C9 3 10 1.95945e-15
C8 4 10 2.38696e-15
C6 6 10 1.79621e-15
C4 8 10 1.63898e-15
C3 9 10 2.11531e-15
C2 10 10 1.95945e-15
C1 11 10 3.2315e-15
.ends nmx2_x1

