-- no model for tie_poly_w2
