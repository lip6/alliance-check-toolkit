* RCClampResistor
.subckt RCClampResistor pin1 pin2

.ends RCClampResistor
