/*                                                                      */
/*  Avertec Release v3.4p5 (64 bits on Linux 5.10.0-0.bpo.9-amd64)      */
/*  [AVT_only] host: fsdev                                              */
/*  [AVT_only] arch: x86_64                                             */
/*  [AVT_only] path: /opt/tasyag-3.4p5/bin/avt_shell                    */
/*  argv:                                                               */
/*                                                                      */
/*  User: verhaegs                                                      */
/*  Generation date Thu Feb 10 13:11:38 2022                            */
/*                                                                      */
/*  Verilog data flow description generated from `one_x1`               */
/*                                                                      */


`timescale 1 ps/1 ps

module one_x1 (one);

  output one;
  assign one = 1;

endmodule
