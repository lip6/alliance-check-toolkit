* Spice description of a4_x2
* Spice driver version 718499611
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:31

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt a4_x2 7 8 4 3 2 1 11 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i3
* NET 4 = i2
* NET 7 = i0
* NET 8 = i1
* NET 11 = vss
Mtr_00010 2 6 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 1 3 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00008 6 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00007 6 7 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00006 1 8 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00005 2 6 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.12U AS=0.5088P AD=0.5088P PS=4.73U PD=4.73U 
Mtr_00004 6 3 5 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00003 5 4 10 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00002 9 7 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00001 10 8 9 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
C11 1 11 2.84014e-15
C10 2 11 2.15173e-15
C9 3 11 1.42163e-15
C8 4 11 1.72566e-15
C6 6 11 2.12904e-15
C5 7 11 1.40338e-15
C4 8 11 1.70741e-15
C1 11 11 2.20267e-15
.ends a4_x2

