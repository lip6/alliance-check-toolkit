.model tp pmos(level=3 kp=40u gamma=0.5 phi=0.36 ld=0.1u tox=20n nsub=4e+16 vmax=2e+5 cj=1.23e-4)
.model tn nmos(level=3 kp=80u gamma=0.4 phi=0.37 ld=0.1u tox=20n nsub=2e+16 vmax=2e+5 cj=3.85e-4)
