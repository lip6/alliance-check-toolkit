* Spice description of oa2a22_x4
* Spice driver version -393371877
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:28

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt oa2a22_x4 8 9 5 4 3 2 11 
* NET 2 = vdd
* NET 3 = q
* NET 4 = i3
* NET 5 = i2
* NET 8 = i0
* NET 9 = i1
* NET 11 = vss
Mtr_00012 1 4 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.78U AS=0.4272P AD=0.4272P PS=4.05U PD=4.05U 
Mtr_00011 3 6 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 2 6 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 6 8 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.78U AS=0.4272P AD=0.4272P PS=4.05U PD=4.05U 
Mtr_00008 2 5 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.78U AS=0.4272P AD=0.4272P PS=4.05U PD=4.05U 
Mtr_00007 1 9 6 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.78U AS=0.4272P AD=0.4272P PS=4.05U PD=4.05U 
Mtr_00006 3 6 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 11 6 3 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 10 8 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00003 11 4 7 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 7 5 6 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 6 9 10 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C11 1 11 9.1453e-16
C10 2 11 3.91506e-15
C9 3 11 2.15173e-15
C8 4 11 1.95384e-15
C7 5 11 1.92646e-15
C6 6 11 3.13739e-15
C4 8 11 1.86257e-15
C3 9 11 1.86257e-15
C1 11 11 3.32564e-15
.ends oa2a22_x4

