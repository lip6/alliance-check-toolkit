* Spice description of inv_x4
* Spice driver version -1910976741
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:42

* INTERF i nq vdd vss 


.subckt inv_x4 2 4 1 3 
* NET 1 = vdd
* NET 2 = i
* NET 3 = vss
* NET 4 = nq
Mtr_00004 4 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00003 1 2 4 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00002 3 2 4 3 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 4 2 3 3 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C4 1 3 1.89615e-15
C3 2 3 2.75301e-15
C2 3 3 1.48915e-15
C1 4 3 2.15173e-15
.ends inv_x4

