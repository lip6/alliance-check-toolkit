-- no model for and4_x1
