* DP8TColumnBlock_128R64B4M8W
* DP8TCell
.subckt DP8TCell vdd vss wl1 wl2 bl1 bl1_n bl2 bl2_n
Mpu1 vdd bit_n bit vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpu2 vdd bit bit_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpd1 vss bit_n bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpd2 vss bit bit_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg1 bl1 wl1 bit vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg1n bl1_n wl1 bit_n vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg2 bl2 wl2 bit vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg2n bl2_n wl2 bit_n vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
.ends DP8TCell
* DP8TArray_2X1
.subckt DP8TArray_2X1 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 vdd vss wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
Xinst1x0 vdd vss wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
.ends DP8TArray_2X1
* DP8TArray_2X2
.subckt DP8TArray_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TArray_2X1
Xinst0x1 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X1
.ends DP8TArray_2X2
* DP8TArray_4X2
.subckt DP8TArray_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
.ends DP8TArray_4X2
* DP8TArray_4X4
.subckt DP8TArray_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X2
.ends DP8TArray_4X4
* DP8TArray_8X4
.subckt DP8TArray_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X4
.ends DP8TArray_8X4
* DP8TArray_8X8
.subckt DP8TArray_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X4
.ends DP8TArray_8X8
* DP8TArray_16X8
.subckt DP8TArray_16X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X8
.ends DP8TArray_16X8
* DP8TArray_16X16
.subckt DP8TArray_16X16 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_16X8
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X8
.ends DP8TArray_16X16
* DP8TArray_32X16
.subckt DP8TArray_32X16 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X16
Xinst1x0 vss vdd wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X16
.ends DP8TArray_32X16
* nand2_x0
.subckt nand2_x0 vdd vss nq i0 i1
Mn0 vss i0 int0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp0 vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn1 int0 i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp1 nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends nand2_x0
* buf_x2
.subckt buf_x2 vdd vss i q
Mn1 ni i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn2_0 vss ni q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn2_1 q ni vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mp1 ni i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp2_0 vdd ni q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp2_1 q ni vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
.ends buf_x2
* inv_x0
.subckt inv_x0 vdd vss i nq
Mn vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends inv_x0
* nor2_x0
.subckt nor2_x0 vdd vss nq i0 i1
Mn0 vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp0 vdd i0 int0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn1 nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp1 int0 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
.ends nor2_x0
* sff1_x4
.subckt sff1_x4 vdd ck vss i q
Mp_ck nckr ck vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_ck nckr ck vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ckr_1 _net1 ckr sff_m vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_ckr_2 y ckr sff_s vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_ckr_1 sff_m ckr _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ckr_2 sff_s ckr _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i u i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i u i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_2 sff_m nckr _net5 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_3 y nckr sff_s vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_1 vdd nckr ckr vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nckr_1 vss nckr ckr vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nckr_3 sff_s nckr _net6 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nckr_2 _net2 nckr sff_m vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_q_1 _net6 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_q_1 _net0 q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_sffm_1 vss sff_m y vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_sffm_1 vdd sff_m y vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_sffs_1 vdd sff_s q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_sffs_1 vss sff_s q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mn_sffs_2 q sff_s vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_sffs_2 q sff_s vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_u vss u _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_u vdd u _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_y_1 _net4 y vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_y_1 _net5 y vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends sff1_x4
* tie
.subckt tie vdd vss

.ends tie
* nsnrlatch_x1
.subckt nsnrlatch_x1 vss nq q vdd nrst nset
Mn_nq_1 _net1 nq vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_nq_1 q nq vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nrst_1 nq nrst vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nrst_1 _net0 nrst nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_nset_1 vdd nset q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nset_1 q nset _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_q_1 vdd q nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_q_1 vss q _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
.ends nsnrlatch_x1
* DP8TArray_32X32
.subckt DP8TArray_32X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_32X16
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X16
.ends DP8TArray_32X32
* DP8TColMux_4C_bl2
.subckt DP8TColMux_4C_bl2 bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl muxbl_n
Mpgbl0 bl[0] mux[0] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln0 muxbl_n mux[0] bl_n[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl1 bl[1] mux[1] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln1 muxbl_n mux[1] bl_n[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl2 bl[2] mux[2] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln2 muxbl_n mux[2] bl_n[2] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl3 bl[3] mux[3] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln3 muxbl_n mux[3] bl_n[3] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
.ends DP8TColMux_4C_bl2
* DP8TPrecharge_bl2
.subckt DP8TPrecharge_bl2 vdd bl bl_n precharge_n
Mpc1 vdd precharge_n bl vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc2 bl precharge_n bl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc3 bl_n precharge_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
.ends DP8TPrecharge_bl2
* DP8TClockWE
.subckt DP8TClockWE vss vdd clkup clklow we we_en we_n
Xclkbuf vdd vss clkup clklow buf_x2
Xweff vdd clklow vss we we_latched sff1_x4
Xwenand vdd vss we_n we_en we_latched nand2_x0
.ends DP8TClockWE
* DP8TWriteDriver_4M2B
.subckt DP8TWriteDriver_4M2B vss vdd clk we_n bl[0] bl_n[0] d[0] bl[1] bl_n[1] d[1]
Xff[0] vdd clk vss d[0] d_latched[0] sff1_x4
Xff[1] vdd clk vss d[1] d_latched[1] sff1_x4
Xnora[0] vdd vss bl_drive[0] d_latched[0] we_n nor2_x0
Xnora[1] vdd vss bl_drive[1] d_latched[1] we_n nor2_x0
Xinv[0] vdd vss d_latched[0] d_n[0] inv_x0
Xinv[1] vdd vss d_latched[1] d_n[1] inv_x0
Xnorb[0] vdd vss bln_drive[0] d_n[0] we_n nor2_x0
Xnorb[1] vdd vss bln_drive[1] d_n[1] we_n nor2_x0
Mblpd[0] vss bl_drive[0] bl[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblpd[1] vss bl_drive[1] bl[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblnpd[0] bl_n[0] bln_drive[0] vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblnpd[1] bl_n[1] bln_drive[1] vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
.ends DP8TWriteDriver_4M2B
* DP8TSenseAmp_4M
.subckt DP8TSenseAmp_4M vss vdd bl bl_n q
Xlatch vss nq q vdd bl bl_n nsnrlatch_x1
Xtie vdd vss tie
.ends DP8TSenseAmp_4M
* DP8TColMux_4C_bl1
.subckt DP8TColMux_4C_bl1 bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl muxbl_n
Mpgbl0 bl[0] mux[0] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln0 muxbl_n mux[0] bl_n[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl1 bl[1] mux[1] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln1 muxbl_n mux[1] bl_n[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl2 bl[2] mux[2] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln2 muxbl_n mux[2] bl_n[2] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl3 bl[3] mux[3] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln3 muxbl_n mux[3] bl_n[3] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
.ends DP8TColMux_4C_bl1
* DP8TPrecharge_bl1
.subckt DP8TPrecharge_bl1 vdd bl bl_n precharge_n
Mpc1 vdd precharge_n bl vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc2 bl precharge_n bl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc3 bl_n precharge_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
.ends DP8TPrecharge_bl1
* DP8TArray_64X32
.subckt DP8TArray_64X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X32
Xinst1x0 vss vdd wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X32
.ends DP8TArray_64X32
* DP8TColumnPeriphery_8B4M_bl2
.subckt DP8TColumnPeriphery_8B4M_bl2 vss vdd clk precharge_n we we_en q[0] d[0] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] q[1] d[1] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] q[2] d[2] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] q[3] d[3] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] q[4] d[4] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] q[5] d[5] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] q[6] d[6] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] q[7] d[7] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] mux[0] mux[1] mux[2] mux[3]
Xprecharge[0] vdd bl[0] bl_n[0] precharge_n DP8TPrecharge_bl2
Xprecharge[1] vdd bl[1] bl_n[1] precharge_n DP8TPrecharge_bl2
Xprecharge[2] vdd bl[2] bl_n[2] precharge_n DP8TPrecharge_bl2
Xprecharge[3] vdd bl[3] bl_n[3] precharge_n DP8TPrecharge_bl2
Xprecharge[4] vdd bl[4] bl_n[4] precharge_n DP8TPrecharge_bl2
Xprecharge[5] vdd bl[5] bl_n[5] precharge_n DP8TPrecharge_bl2
Xprecharge[6] vdd bl[6] bl_n[6] precharge_n DP8TPrecharge_bl2
Xprecharge[7] vdd bl[7] bl_n[7] precharge_n DP8TPrecharge_bl2
Xprecharge[8] vdd bl[8] bl_n[8] precharge_n DP8TPrecharge_bl2
Xprecharge[9] vdd bl[9] bl_n[9] precharge_n DP8TPrecharge_bl2
Xprecharge[10] vdd bl[10] bl_n[10] precharge_n DP8TPrecharge_bl2
Xprecharge[11] vdd bl[11] bl_n[11] precharge_n DP8TPrecharge_bl2
Xprecharge[12] vdd bl[12] bl_n[12] precharge_n DP8TPrecharge_bl2
Xprecharge[13] vdd bl[13] bl_n[13] precharge_n DP8TPrecharge_bl2
Xprecharge[14] vdd bl[14] bl_n[14] precharge_n DP8TPrecharge_bl2
Xprecharge[15] vdd bl[15] bl_n[15] precharge_n DP8TPrecharge_bl2
Xprecharge[16] vdd bl[16] bl_n[16] precharge_n DP8TPrecharge_bl2
Xprecharge[17] vdd bl[17] bl_n[17] precharge_n DP8TPrecharge_bl2
Xprecharge[18] vdd bl[18] bl_n[18] precharge_n DP8TPrecharge_bl2
Xprecharge[19] vdd bl[19] bl_n[19] precharge_n DP8TPrecharge_bl2
Xprecharge[20] vdd bl[20] bl_n[20] precharge_n DP8TPrecharge_bl2
Xprecharge[21] vdd bl[21] bl_n[21] precharge_n DP8TPrecharge_bl2
Xprecharge[22] vdd bl[22] bl_n[22] precharge_n DP8TPrecharge_bl2
Xprecharge[23] vdd bl[23] bl_n[23] precharge_n DP8TPrecharge_bl2
Xprecharge[24] vdd bl[24] bl_n[24] precharge_n DP8TPrecharge_bl2
Xprecharge[25] vdd bl[25] bl_n[25] precharge_n DP8TPrecharge_bl2
Xprecharge[26] vdd bl[26] bl_n[26] precharge_n DP8TPrecharge_bl2
Xprecharge[27] vdd bl[27] bl_n[27] precharge_n DP8TPrecharge_bl2
Xprecharge[28] vdd bl[28] bl_n[28] precharge_n DP8TPrecharge_bl2
Xprecharge[29] vdd bl[29] bl_n[29] precharge_n DP8TPrecharge_bl2
Xprecharge[30] vdd bl[30] bl_n[30] precharge_n DP8TPrecharge_bl2
Xprecharge[31] vdd bl[31] bl_n[31] precharge_n DP8TPrecharge_bl2
Xcolmux[0] bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl[0] muxbl_n[0] DP8TColMux_4C_bl2
Xcolmux[1] bl[4] bl_n[4] mux[0] bl[5] bl_n[5] mux[1] bl[6] bl_n[6] mux[2] bl[7] bl_n[7] mux[3] vss muxbl[1] muxbl_n[1] DP8TColMux_4C_bl2
Xcolmux[2] bl[8] bl_n[8] mux[0] bl[9] bl_n[9] mux[1] bl[10] bl_n[10] mux[2] bl[11] bl_n[11] mux[3] vss muxbl[2] muxbl_n[2] DP8TColMux_4C_bl2
Xcolmux[3] bl[12] bl_n[12] mux[0] bl[13] bl_n[13] mux[1] bl[14] bl_n[14] mux[2] bl[15] bl_n[15] mux[3] vss muxbl[3] muxbl_n[3] DP8TColMux_4C_bl2
Xcolmux[4] bl[16] bl_n[16] mux[0] bl[17] bl_n[17] mux[1] bl[18] bl_n[18] mux[2] bl[19] bl_n[19] mux[3] vss muxbl[4] muxbl_n[4] DP8TColMux_4C_bl2
Xcolmux[5] bl[20] bl_n[20] mux[0] bl[21] bl_n[21] mux[1] bl[22] bl_n[22] mux[2] bl[23] bl_n[23] mux[3] vss muxbl[5] muxbl_n[5] DP8TColMux_4C_bl2
Xcolmux[6] bl[24] bl_n[24] mux[0] bl[25] bl_n[25] mux[1] bl[26] bl_n[26] mux[2] bl[27] bl_n[27] mux[3] vss muxbl[6] muxbl_n[6] DP8TColMux_4C_bl2
Xcolmux[7] bl[28] bl_n[28] mux[0] bl[29] bl_n[29] mux[1] bl[30] bl_n[30] mux[2] bl[31] bl_n[31] mux[3] vss muxbl[7] muxbl_n[7] DP8TColMux_4C_bl2
Xsenseamp[0] vss vdd muxbl[0] muxbl_n[0] q[0] DP8TSenseAmp_4M
Xsenseamp[1] vss vdd muxbl[1] muxbl_n[1] q[1] DP8TSenseAmp_4M
Xsenseamp[2] vss vdd muxbl[2] muxbl_n[2] q[2] DP8TSenseAmp_4M
Xsenseamp[3] vss vdd muxbl[3] muxbl_n[3] q[3] DP8TSenseAmp_4M
Xsenseamp[4] vss vdd muxbl[4] muxbl_n[4] q[4] DP8TSenseAmp_4M
Xsenseamp[5] vss vdd muxbl[5] muxbl_n[5] q[5] DP8TSenseAmp_4M
Xsenseamp[6] vss vdd muxbl[6] muxbl_n[6] q[6] DP8TSenseAmp_4M
Xsenseamp[7] vss vdd muxbl[7] muxbl_n[7] q[7] DP8TSenseAmp_4M
Xwritedrive[0] vss vdd intclk we_n muxbl[0] muxbl_n[0] d[0] muxbl[1] muxbl_n[1] d[1] DP8TWriteDriver_4M2B
Xwritedrive[1] vss vdd intclk we_n muxbl[2] muxbl_n[2] d[2] muxbl[3] muxbl_n[3] d[3] DP8TWriteDriver_4M2B
Xwritedrive[2] vss vdd intclk we_n muxbl[4] muxbl_n[4] d[4] muxbl[5] muxbl_n[5] d[5] DP8TWriteDriver_4M2B
Xwritedrive[3] vss vdd intclk we_n muxbl[6] muxbl_n[6] d[6] muxbl[7] muxbl_n[7] d[7] DP8TWriteDriver_4M2B
Xclkwe vss vdd clk intclk we we_en we_n DP8TClockWE
.ends DP8TColumnPeriphery_8B4M_bl2
* DP8TColumnPeriphery_8B4M_bl1
.subckt DP8TColumnPeriphery_8B4M_bl1 vss vdd clk precharge_n we we_en q[0] d[0] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] q[1] d[1] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] q[2] d[2] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] q[3] d[3] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] q[4] d[4] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] q[5] d[5] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] q[6] d[6] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] q[7] d[7] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] mux[0] mux[1] mux[2] mux[3]
Xprecharge[0] vdd bl[0] bl_n[0] precharge_n DP8TPrecharge_bl1
Xprecharge[1] vdd bl[1] bl_n[1] precharge_n DP8TPrecharge_bl1
Xprecharge[2] vdd bl[2] bl_n[2] precharge_n DP8TPrecharge_bl1
Xprecharge[3] vdd bl[3] bl_n[3] precharge_n DP8TPrecharge_bl1
Xprecharge[4] vdd bl[4] bl_n[4] precharge_n DP8TPrecharge_bl1
Xprecharge[5] vdd bl[5] bl_n[5] precharge_n DP8TPrecharge_bl1
Xprecharge[6] vdd bl[6] bl_n[6] precharge_n DP8TPrecharge_bl1
Xprecharge[7] vdd bl[7] bl_n[7] precharge_n DP8TPrecharge_bl1
Xprecharge[8] vdd bl[8] bl_n[8] precharge_n DP8TPrecharge_bl1
Xprecharge[9] vdd bl[9] bl_n[9] precharge_n DP8TPrecharge_bl1
Xprecharge[10] vdd bl[10] bl_n[10] precharge_n DP8TPrecharge_bl1
Xprecharge[11] vdd bl[11] bl_n[11] precharge_n DP8TPrecharge_bl1
Xprecharge[12] vdd bl[12] bl_n[12] precharge_n DP8TPrecharge_bl1
Xprecharge[13] vdd bl[13] bl_n[13] precharge_n DP8TPrecharge_bl1
Xprecharge[14] vdd bl[14] bl_n[14] precharge_n DP8TPrecharge_bl1
Xprecharge[15] vdd bl[15] bl_n[15] precharge_n DP8TPrecharge_bl1
Xprecharge[16] vdd bl[16] bl_n[16] precharge_n DP8TPrecharge_bl1
Xprecharge[17] vdd bl[17] bl_n[17] precharge_n DP8TPrecharge_bl1
Xprecharge[18] vdd bl[18] bl_n[18] precharge_n DP8TPrecharge_bl1
Xprecharge[19] vdd bl[19] bl_n[19] precharge_n DP8TPrecharge_bl1
Xprecharge[20] vdd bl[20] bl_n[20] precharge_n DP8TPrecharge_bl1
Xprecharge[21] vdd bl[21] bl_n[21] precharge_n DP8TPrecharge_bl1
Xprecharge[22] vdd bl[22] bl_n[22] precharge_n DP8TPrecharge_bl1
Xprecharge[23] vdd bl[23] bl_n[23] precharge_n DP8TPrecharge_bl1
Xprecharge[24] vdd bl[24] bl_n[24] precharge_n DP8TPrecharge_bl1
Xprecharge[25] vdd bl[25] bl_n[25] precharge_n DP8TPrecharge_bl1
Xprecharge[26] vdd bl[26] bl_n[26] precharge_n DP8TPrecharge_bl1
Xprecharge[27] vdd bl[27] bl_n[27] precharge_n DP8TPrecharge_bl1
Xprecharge[28] vdd bl[28] bl_n[28] precharge_n DP8TPrecharge_bl1
Xprecharge[29] vdd bl[29] bl_n[29] precharge_n DP8TPrecharge_bl1
Xprecharge[30] vdd bl[30] bl_n[30] precharge_n DP8TPrecharge_bl1
Xprecharge[31] vdd bl[31] bl_n[31] precharge_n DP8TPrecharge_bl1
Xcolmux[0] bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl[0] muxbl_n[0] DP8TColMux_4C_bl1
Xcolmux[1] bl[4] bl_n[4] mux[0] bl[5] bl_n[5] mux[1] bl[6] bl_n[6] mux[2] bl[7] bl_n[7] mux[3] vss muxbl[1] muxbl_n[1] DP8TColMux_4C_bl1
Xcolmux[2] bl[8] bl_n[8] mux[0] bl[9] bl_n[9] mux[1] bl[10] bl_n[10] mux[2] bl[11] bl_n[11] mux[3] vss muxbl[2] muxbl_n[2] DP8TColMux_4C_bl1
Xcolmux[3] bl[12] bl_n[12] mux[0] bl[13] bl_n[13] mux[1] bl[14] bl_n[14] mux[2] bl[15] bl_n[15] mux[3] vss muxbl[3] muxbl_n[3] DP8TColMux_4C_bl1
Xcolmux[4] bl[16] bl_n[16] mux[0] bl[17] bl_n[17] mux[1] bl[18] bl_n[18] mux[2] bl[19] bl_n[19] mux[3] vss muxbl[4] muxbl_n[4] DP8TColMux_4C_bl1
Xcolmux[5] bl[20] bl_n[20] mux[0] bl[21] bl_n[21] mux[1] bl[22] bl_n[22] mux[2] bl[23] bl_n[23] mux[3] vss muxbl[5] muxbl_n[5] DP8TColMux_4C_bl1
Xcolmux[6] bl[24] bl_n[24] mux[0] bl[25] bl_n[25] mux[1] bl[26] bl_n[26] mux[2] bl[27] bl_n[27] mux[3] vss muxbl[6] muxbl_n[6] DP8TColMux_4C_bl1
Xcolmux[7] bl[28] bl_n[28] mux[0] bl[29] bl_n[29] mux[1] bl[30] bl_n[30] mux[2] bl[31] bl_n[31] mux[3] vss muxbl[7] muxbl_n[7] DP8TColMux_4C_bl1
Xsenseamp[0] vss vdd muxbl[0] muxbl_n[0] q[0] DP8TSenseAmp_4M
Xsenseamp[1] vss vdd muxbl[1] muxbl_n[1] q[1] DP8TSenseAmp_4M
Xsenseamp[2] vss vdd muxbl[2] muxbl_n[2] q[2] DP8TSenseAmp_4M
Xsenseamp[3] vss vdd muxbl[3] muxbl_n[3] q[3] DP8TSenseAmp_4M
Xsenseamp[4] vss vdd muxbl[4] muxbl_n[4] q[4] DP8TSenseAmp_4M
Xsenseamp[5] vss vdd muxbl[5] muxbl_n[5] q[5] DP8TSenseAmp_4M
Xsenseamp[6] vss vdd muxbl[6] muxbl_n[6] q[6] DP8TSenseAmp_4M
Xsenseamp[7] vss vdd muxbl[7] muxbl_n[7] q[7] DP8TSenseAmp_4M
Xwritedrive[0] vss vdd intclk we_n muxbl[0] muxbl_n[0] d[0] muxbl[1] muxbl_n[1] d[1] DP8TWriteDriver_4M2B
Xwritedrive[1] vss vdd intclk we_n muxbl[2] muxbl_n[2] d[2] muxbl[3] muxbl_n[3] d[3] DP8TWriteDriver_4M2B
Xwritedrive[2] vss vdd intclk we_n muxbl[4] muxbl_n[4] d[4] muxbl[5] muxbl_n[5] d[5] DP8TWriteDriver_4M2B
Xwritedrive[3] vss vdd intclk we_n muxbl[6] muxbl_n[6] d[6] muxbl[7] muxbl_n[7] d[7] DP8TWriteDriver_4M2B
Xclkwe vss vdd clk intclk we we_en we_n DP8TClockWE
.ends DP8TColumnPeriphery_8B4M_bl1
* DP8TArray_128X32
.subckt DP8TArray_128X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_64X32
Xinst1x0 vss vdd wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_64X32
.ends DP8TArray_128X32
* DP8TColumn_128R8B4M
.subckt DP8TColumn_128R8B4M vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1 clk1 we_en1 precharge1_n we2 clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3]
Xarray vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_128X32
Xperiph1 vss vdd clk1 precharge1_n we1 we_en1 q1[0] d1[0] bl1[0] bl1_n[0] bl1[1] bl1_n[1] bl1[2] bl1_n[2] bl1[3] bl1_n[3] q1[1] d1[1] bl1[4] bl1_n[4] bl1[5] bl1_n[5] bl1[6] bl1_n[6] bl1[7] bl1_n[7] q1[2] d1[2] bl1[8] bl1_n[8] bl1[9] bl1_n[9] bl1[10] bl1_n[10] bl1[11] bl1_n[11] q1[3] d1[3] bl1[12] bl1_n[12] bl1[13] bl1_n[13] bl1[14] bl1_n[14] bl1[15] bl1_n[15] q1[4] d1[4] bl1[16] bl1_n[16] bl1[17] bl1_n[17] bl1[18] bl1_n[18] bl1[19] bl1_n[19] q1[5] d1[5] bl1[20] bl1_n[20] bl1[21] bl1_n[21] bl1[22] bl1_n[22] bl1[23] bl1_n[23] q1[6] d1[6] bl1[24] bl1_n[24] bl1[25] bl1_n[25] bl1[26] bl1_n[26] bl1[27] bl1_n[27] q1[7] d1[7] bl1[28] bl1_n[28] bl1[29] bl1_n[29] bl1[30] bl1_n[30] bl1[31] bl1_n[31] mux1[0] mux1[1] mux1[2] mux1[3] DP8TColumnPeriphery_8B4M_bl1
Xperiph2 vss vdd clk2 precharge2_n we2 we_en2 q2[0] d2[0] bl2[0] bl2_n[0] bl2[1] bl2_n[1] bl2[2] bl2_n[2] bl2[3] bl2_n[3] q2[1] d2[1] bl2[4] bl2_n[4] bl2[5] bl2_n[5] bl2[6] bl2_n[6] bl2[7] bl2_n[7] q2[2] d2[2] bl2[8] bl2_n[8] bl2[9] bl2_n[9] bl2[10] bl2_n[10] bl2[11] bl2_n[11] q2[3] d2[3] bl2[12] bl2_n[12] bl2[13] bl2_n[13] bl2[14] bl2_n[14] bl2[15] bl2_n[15] q2[4] d2[4] bl2[16] bl2_n[16] bl2[17] bl2_n[17] bl2[18] bl2_n[18] bl2[19] bl2_n[19] q2[5] d2[5] bl2[20] bl2_n[20] bl2[21] bl2_n[21] bl2[22] bl2_n[22] bl2[23] bl2_n[23] q2[6] d2[6] bl2[24] bl2_n[24] bl2[25] bl2_n[25] bl2[26] bl2_n[26] bl2[27] bl2_n[27] q2[7] d2[7] bl2[28] bl2_n[28] bl2[29] bl2_n[29] bl2[30] bl2_n[30] bl2[31] bl2_n[31] mux2[0] mux2[1] mux2[2] mux2[3] DP8TColumnPeriphery_8B4M_bl2
.ends DP8TColumn_128R8B4M
* DP8TColumnBlock_128R64B4M8W
.subckt DP8TColumnBlock_128R64B4M8W vss vdd clk1 clk2 precharge1_n precharge2_n we_en1 we_en2 wl1[0] wl1[1] wl1[2] wl1[3] wl1[4] wl1[5] wl1[6] wl1[7] wl1[8] wl1[9] wl1[10] wl1[11] wl1[12] wl1[13] wl1[14] wl1[15] wl1[16] wl1[17] wl1[18] wl1[19] wl1[20] wl1[21] wl1[22] wl1[23] wl1[24] wl1[25] wl1[26] wl1[27] wl1[28] wl1[29] wl1[30] wl1[31] wl1[32] wl1[33] wl1[34] wl1[35] wl1[36] wl1[37] wl1[38] wl1[39] wl1[40] wl1[41] wl1[42] wl1[43] wl1[44] wl1[45] wl1[46] wl1[47] wl1[48] wl1[49] wl1[50] wl1[51] wl1[52] wl1[53] wl1[54] wl1[55] wl1[56] wl1[57] wl1[58] wl1[59] wl1[60] wl1[61] wl1[62] wl1[63] wl1[64] wl1[65] wl1[66] wl1[67] wl1[68] wl1[69] wl1[70] wl1[71] wl1[72] wl1[73] wl1[74] wl1[75] wl1[76] wl1[77] wl1[78] wl1[79] wl1[80] wl1[81] wl1[82] wl1[83] wl1[84] wl1[85] wl1[86] wl1[87] wl1[88] wl1[89] wl1[90] wl1[91] wl1[92] wl1[93] wl1[94] wl1[95] wl1[96] wl1[97] wl1[98] wl1[99] wl1[100] wl1[101] wl1[102] wl1[103] wl1[104] wl1[105] wl1[106] wl1[107] wl1[108] wl1[109] wl1[110] wl1[111] wl1[112] wl1[113] wl1[114] wl1[115] wl1[116] wl1[117] wl1[118] wl1[119] wl1[120] wl1[121] wl1[122] wl1[123] wl1[124] wl1[125] wl1[126] wl1[127] wl2[0] wl2[1] wl2[2] wl2[3] wl2[4] wl2[5] wl2[6] wl2[7] wl2[8] wl2[9] wl2[10] wl2[11] wl2[12] wl2[13] wl2[14] wl2[15] wl2[16] wl2[17] wl2[18] wl2[19] wl2[20] wl2[21] wl2[22] wl2[23] wl2[24] wl2[25] wl2[26] wl2[27] wl2[28] wl2[29] wl2[30] wl2[31] wl2[32] wl2[33] wl2[34] wl2[35] wl2[36] wl2[37] wl2[38] wl2[39] wl2[40] wl2[41] wl2[42] wl2[43] wl2[44] wl2[45] wl2[46] wl2[47] wl2[48] wl2[49] wl2[50] wl2[51] wl2[52] wl2[53] wl2[54] wl2[55] wl2[56] wl2[57] wl2[58] wl2[59] wl2[60] wl2[61] wl2[62] wl2[63] wl2[64] wl2[65] wl2[66] wl2[67] wl2[68] wl2[69] wl2[70] wl2[71] wl2[72] wl2[73] wl2[74] wl2[75] wl2[76] wl2[77] wl2[78] wl2[79] wl2[80] wl2[81] wl2[82] wl2[83] wl2[84] wl2[85] wl2[86] wl2[87] wl2[88] wl2[89] wl2[90] wl2[91] wl2[92] wl2[93] wl2[94] wl2[95] wl2[96] wl2[97] wl2[98] wl2[99] wl2[100] wl2[101] wl2[102] wl2[103] wl2[104] wl2[105] wl2[106] wl2[107] wl2[108] wl2[109] wl2[110] wl2[111] wl2[112] wl2[113] wl2[114] wl2[115] wl2[116] wl2[117] wl2[118] wl2[119] wl2[120] wl2[121] wl2[122] wl2[123] wl2[124] wl2[125] wl2[126] wl2[127] mux1[0] mux1[1] mux1[2] mux1[3] mux2[0] mux2[1] mux2[2] mux2[3] we1[0] we2[0] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1[1] we2[1] q1[8] q2[8] d1[8] d2[8] q1[9] q2[9] d1[9] d2[9] q1[10] q2[10] d1[10] d2[10] q1[11] q2[11] d1[11] d2[11] q1[12] q2[12] d1[12] d2[12] q1[13] q2[13] d1[13] d2[13] q1[14] q2[14] d1[14] d2[14] q1[15] q2[15] d1[15] d2[15] we1[2] we2[2] q1[16] q2[16] d1[16] d2[16] q1[17] q2[17] d1[17] d2[17] q1[18] q2[18] d1[18] d2[18] q1[19] q2[19] d1[19] d2[19] q1[20] q2[20] d1[20] d2[20] q1[21] q2[21] d1[21] d2[21] q1[22] q2[22] d1[22] d2[22] q1[23] q2[23] d1[23] d2[23] we1[3] we2[3] q1[24] q2[24] d1[24] d2[24] q1[25] q2[25] d1[25] d2[25] q1[26] q2[26] d1[26] d2[26] q1[27] q2[27] d1[27] d2[27] q1[28] q2[28] d1[28] d2[28] q1[29] q2[29] d1[29] d2[29] q1[30] q2[30] d1[30] d2[30] q1[31] q2[31] d1[31] d2[31] we1[4] we2[4] q1[32] q2[32] d1[32] d2[32] q1[33] q2[33] d1[33] d2[33] q1[34] q2[34] d1[34] d2[34] q1[35] q2[35] d1[35] d2[35] q1[36] q2[36] d1[36] d2[36] q1[37] q2[37] d1[37] d2[37] q1[38] q2[38] d1[38] d2[38] q1[39] q2[39] d1[39] d2[39] we1[5] we2[5] q1[40] q2[40] d1[40] d2[40] q1[41] q2[41] d1[41] d2[41] q1[42] q2[42] d1[42] d2[42] q1[43] q2[43] d1[43] d2[43] q1[44] q2[44] d1[44] d2[44] q1[45] q2[45] d1[45] d2[45] q1[46] q2[46] d1[46] d2[46] q1[47] q2[47] d1[47] d2[47] we1[6] we2[6] q1[48] q2[48] d1[48] d2[48] q1[49] q2[49] d1[49] d2[49] q1[50] q2[50] d1[50] d2[50] q1[51] q2[51] d1[51] d2[51] q1[52] q2[52] d1[52] d2[52] q1[53] q2[53] d1[53] d2[53] q1[54] q2[54] d1[54] d2[54] q1[55] q2[55] d1[55] d2[55] we1[7] we2[7] q1[56] q2[56] d1[56] d2[56] q1[57] q2[57] d1[57] d2[57] q1[58] q2[58] d1[58] d2[58] q1[59] q2[59] d1[59] d2[59] q1[60] q2[60] d1[60] d2[60] q1[61] q2[61] d1[61] d2[61] q1[62] q2[62] d1[62] d2[62] q1[63] q2[63] d1[63] d2[63]
Xcolumn[0] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1[0] clk1 we_en1 precharge1_n we2[0] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[1] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[8] q2[8] d1[8] d2[8] q1[9] q2[9] d1[9] d2[9] q1[10] q2[10] d1[10] d2[10] q1[11] q2[11] d1[11] d2[11] q1[12] q2[12] d1[12] d2[12] q1[13] q2[13] d1[13] d2[13] q1[14] q2[14] d1[14] d2[14] q1[15] q2[15] d1[15] d2[15] we1[1] clk1 we_en1 precharge1_n we2[1] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[2] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[16] q2[16] d1[16] d2[16] q1[17] q2[17] d1[17] d2[17] q1[18] q2[18] d1[18] d2[18] q1[19] q2[19] d1[19] d2[19] q1[20] q2[20] d1[20] d2[20] q1[21] q2[21] d1[21] d2[21] q1[22] q2[22] d1[22] d2[22] q1[23] q2[23] d1[23] d2[23] we1[2] clk1 we_en1 precharge1_n we2[2] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[3] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[24] q2[24] d1[24] d2[24] q1[25] q2[25] d1[25] d2[25] q1[26] q2[26] d1[26] d2[26] q1[27] q2[27] d1[27] d2[27] q1[28] q2[28] d1[28] d2[28] q1[29] q2[29] d1[29] d2[29] q1[30] q2[30] d1[30] d2[30] q1[31] q2[31] d1[31] d2[31] we1[3] clk1 we_en1 precharge1_n we2[3] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[4] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[32] q2[32] d1[32] d2[32] q1[33] q2[33] d1[33] d2[33] q1[34] q2[34] d1[34] d2[34] q1[35] q2[35] d1[35] d2[35] q1[36] q2[36] d1[36] d2[36] q1[37] q2[37] d1[37] d2[37] q1[38] q2[38] d1[38] d2[38] q1[39] q2[39] d1[39] d2[39] we1[4] clk1 we_en1 precharge1_n we2[4] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[5] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[40] q2[40] d1[40] d2[40] q1[41] q2[41] d1[41] d2[41] q1[42] q2[42] d1[42] d2[42] q1[43] q2[43] d1[43] d2[43] q1[44] q2[44] d1[44] d2[44] q1[45] q2[45] d1[45] d2[45] q1[46] q2[46] d1[46] d2[46] q1[47] q2[47] d1[47] d2[47] we1[5] clk1 we_en1 precharge1_n we2[5] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[6] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[48] q2[48] d1[48] d2[48] q1[49] q2[49] d1[49] d2[49] q1[50] q2[50] d1[50] d2[50] q1[51] q2[51] d1[51] d2[51] q1[52] q2[52] d1[52] d2[52] q1[53] q2[53] d1[53] d2[53] q1[54] q2[54] d1[54] d2[54] q1[55] q2[55] d1[55] d2[55] we1[6] clk1 we_en1 precharge1_n we2[6] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[7] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[56] q2[56] d1[56] d2[56] q1[57] q2[57] d1[57] d2[57] q1[58] q2[58] d1[58] d2[58] q1[59] q2[59] d1[59] d2[59] q1[60] q2[60] d1[60] d2[60] q1[61] q2[61] d1[61] d2[61] q1[62] q2[62] d1[62] d2[62] q1[63] q2[63] d1[63] d2[63] we1[7] clk1 we_en1 precharge1_n we2[7] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
.ends DP8TColumnBlock_128R64B4M8W
