* BulkConn_2000WNoUp
.subckt BulkConn_2000WNoUp vdd vss iovdd iovss

.ends BulkConn_2000WNoUp
