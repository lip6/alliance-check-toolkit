* GuardRing_P17368W3836HFF
.subckt GuardRing_P17368W3836HFF conn

.ends GuardRing_P17368W3836HFF
