* NPN_05v5_W1u00L2u00
* NPN_05v5_W1u00L2u00
.subckt NPN_05v5_W1u00L2u00 collector base emitter
Xnpn collector base emitter sky130_fd_pr__npn_05v5_W1p00L2p00
.ends NPN_05v5_W1u00L2u00
