*
* top_inv_x2.spi
* ngspice simulation
* 

*****************

.TEMP 25

******************
* BSIM4 transistor model parameters for ngspice
*.lib /users/soft/analogdesign/scalable/techno/sky130_models_20220217/C4M.Sky130_all_lib.spice logic_tt 

*******************************
*Simulation conditions

Vground evss 0 0
Vsupply evdd 0 DC 1.8
*gfoncd evdd 0 evdd 0 1.0e-15

******************
* circuit model
* include circuit netlist
.INCLUDE inv_x2.spi
*****************

*****************
* Circuit Instantiation
*.subckt inv_x2 vdd vss i nq

Xc evdd evss in out inv_x2

.end

