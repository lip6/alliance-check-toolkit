* Spice description of buf_x4
* Spice driver version -529400037
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:39

* INTERF i q vdd vss 


.subckt buf_x4 3 2 1 4 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i
* NET 4 = vss
Mtr_00006 1 5 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.23U AS=0.7752P AD=0.7752P PS=6.94U PD=6.94U 
Mtr_00005 2 5 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.23U AS=0.7752P AD=0.7752P PS=6.94U PD=6.94U 
Mtr_00004 1 3 5 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00003 4 5 2 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00002 2 5 4 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00001 4 3 5 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C5 1 4 2.14102e-15
C4 2 4 2.15173e-15
C3 3 4 2.45696e-15
C2 4 4 1.73402e-15
C1 5 4 1.89409e-15
.ends buf_x4

