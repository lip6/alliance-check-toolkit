-- no model for fill_w2
