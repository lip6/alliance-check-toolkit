* Spice description of arlet6502_cts_r
* Spice driver version -777225304
* Date ( dd/mm/yyyy hh:mm:ss ):  7/06/2024 at  1:11:39

* INTERF a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] a[9] a[10] a[11] a[12] 
* INTERF a[13] a[14] a[15] clk di[0] di[1] di[2] di[3] di[4] di[5] di[6] 
* INTERF di[7] do[0] do[1] do[2] do[3] do[4] do[5] do[6] do[7] irq nmi rdy 
* INTERF reset vdd vss we 


.subckt arlet6502_cts_r 3012 2081 2717 2024 2073 2003 4524 4240 3263 11039 11012 10977 10951 10917 10877 10847 5554 10901 10789 10620 9505 9316 8840 8064 6465 3425 2416 2427 1815 10081 8816 8017 6793 5811 2373 5611 5199 11024 11074 1877 
* NET 119 = subckt_1739_sff1_x4.sff_s
* NET 121 = subckt_1739_sff1_x4.y
* NET 123 = subckt_1739_sff1_x4.sff_m
* NET 124 = subckt_1739_sff1_x4.u
* NET 125 = subckt_1739_sff1_x4.ckr
* NET 126 = subckt_1739_sff1_x4.nckr
* NET 127 = subckt_1622_sff1_x4.sff_s
* NET 129 = subckt_1622_sff1_x4.y
* NET 130 = subckt_1622_sff1_x4.sff_m
* NET 133 = subckt_1622_sff1_x4.u
* NET 134 = subckt_1622_sff1_x4.ckr
* NET 135 = subckt_1622_sff1_x4.nckr
* NET 137 = subckt_1623_sff1_x4.sff_s
* NET 139 = subckt_1623_sff1_x4.y
* NET 141 = subckt_1623_sff1_x4.sff_m
* NET 142 = subckt_1623_sff1_x4.u
* NET 143 = subckt_1623_sff1_x4.ckr
* NET 144 = subckt_1623_sff1_x4.nckr
* NET 145 = abc_11867_auto_rtlil_cc_2608_muxgate_11616
* NET 150 = subckt_1637_sff1_x4.sff_s
* NET 153 = subckt_1637_sff1_x4.y
* NET 154 = subckt_1637_sff1_x4.sff_m
* NET 155 = subckt_1637_sff1_x4.u
* NET 157 = subckt_1637_sff1_x4.ckr
* NET 158 = subckt_1637_sff1_x4.nckr
* NET 160 = subckt_1650_sff1_x4.sff_s
* NET 162 = subckt_1650_sff1_x4.y
* NET 164 = subckt_1650_sff1_x4.sff_m
* NET 165 = subckt_1650_sff1_x4.u
* NET 166 = subckt_1650_sff1_x4.ckr
* NET 167 = subckt_1650_sff1_x4.nckr
* NET 169 = subckt_1632_sff1_x4.sff_s
* NET 170 = subckt_1632_sff1_x4.y
* NET 173 = subckt_1632_sff1_x4.sff_m
* NET 174 = subckt_1632_sff1_x4.u
* NET 175 = subckt_1632_sff1_x4.ckr
* NET 176 = subckt_1632_sff1_x4.nckr
* NET 177 = subckt_1647_sff1_x4.sff_s
* NET 179 = subckt_1647_sff1_x4.y
* NET 180 = subckt_1647_sff1_x4.sff_m
* NET 183 = subckt_1647_sff1_x4.u
* NET 184 = subckt_1647_sff1_x4.ckr
* NET 185 = subckt_1647_sff1_x4.nckr
* NET 187 = subckt_1617_sff1_x4.sff_s
* NET 188 = subckt_1617_sff1_x4.y
* NET 190 = subckt_1617_sff1_x4.sff_m
* NET 192 = subckt_1617_sff1_x4.u
* NET 193 = subckt_1617_sff1_x4.ckr
* NET 194 = subckt_1617_sff1_x4.nckr
* NET 195 = abc_11867_auto_rtlil_cc_2608_muxgate_11604
* NET 200 = subckt_1631_sff1_x4.sff_s
* NET 202 = subckt_1631_sff1_x4.y
* NET 203 = subckt_1631_sff1_x4.sff_m
* NET 206 = subckt_1631_sff1_x4.u
* NET 207 = subckt_1631_sff1_x4.ckr
* NET 208 = subckt_1631_sff1_x4.nckr
* NET 213 = abc_11867_new_n872
* NET 215 = abc_11867_new_n871
* NET 217 = abc_11867_new_n877
* NET 219 = abc_11867_new_n860
* NET 220 = abc_11867_new_n878
* NET 223 = subckt_1655_sff1_x4.sff_s
* NET 224 = subckt_1655_sff1_x4.y
* NET 227 = subckt_1655_sff1_x4.sff_m
* NET 228 = subckt_1655_sff1_x4.u
* NET 229 = subckt_1655_sff1_x4.ckr
* NET 230 = subckt_1655_sff1_x4.nckr
* NET 231 = abc_11867_auto_rtlil_cc_2608_muxgate_11670
* NET 238 = abc_11867_new_n608
* NET 241 = abc_11867_new_n1175
* NET 244 = mos6502_nmi_1
* NET 246 = subckt_1656_sff1_x4.sff_s
* NET 247 = subckt_1656_sff1_x4.y
* NET 250 = subckt_1656_sff1_x4.sff_m
* NET 251 = subckt_1656_sff1_x4.u
* NET 252 = subckt_1656_sff1_x4.ckr
* NET 253 = subckt_1656_sff1_x4.nckr
* NET 311 = subckt_1653_sff1_x4.sff_s
* NET 312 = subckt_1653_sff1_x4.y
* NET 316 = subckt_1653_sff1_x4.sff_m
* NET 317 = subckt_1653_sff1_x4.ckr
* NET 318 = subckt_1653_sff1_x4.u
* NET 319 = subckt_1653_sff1_x4.nckr
* NET 320 = abc_11867_auto_rtlil_cc_2608_muxgate_11664
* NET 329 = abc_11867_auto_rtlil_cc_2608_muxgate_11614
* NET 338 = mos6502_axys_2_6
* NET 341 = mos6502_axys_3_6
* NET 347 = abc_11867_auto_rtlil_cc_2608_muxgate_11632
* NET 348 = mos6502_axys_0_6
* NET 358 = subckt_1648_sff1_x4.sff_s
* NET 360 = subckt_1648_sff1_x4.y
* NET 364 = subckt_1648_sff1_x4.sff_m
* NET 365 = subckt_1648_sff1_x4.u
* NET 366 = subckt_1648_sff1_x4.ckr
* NET 367 = subckt_1648_sff1_x4.nckr
* NET 368 = abc_11867_auto_rtlil_cc_2608_muxgate_11654
* NET 377 = abc_11867_auto_rtlil_cc_2608_muxgate_11622
* NET 388 = subckt_1634_sff1_x4.sff_s
* NET 389 = subckt_1634_sff1_x4.y
* NET 393 = subckt_1634_sff1_x4.sff_m
* NET 394 = subckt_1634_sff1_x4.ckr
* NET 395 = subckt_1634_sff1_x4.u
* NET 396 = subckt_1634_sff1_x4.nckr
* NET 397 = abc_11867_auto_rtlil_cc_2608_muxgate_11652
* NET 407 = subckt_1649_sff1_x4.sff_s
* NET 411 = subckt_1649_sff1_x4.y
* NET 412 = subckt_1649_sff1_x4.sff_m
* NET 414 = subckt_1649_sff1_x4.ckr
* NET 415 = subckt_1649_sff1_x4.u
* NET 416 = subckt_1649_sff1_x4.nckr
* NET 419 = abc_11867_auto_rtlil_cc_2608_muxgate_11620
* NET 428 = subckt_1633_sff1_x4.sff_s
* NET 429 = subckt_1633_sff1_x4.y
* NET 432 = subckt_1633_sff1_x4.sff_m
* NET 434 = subckt_1633_sff1_x4.u
* NET 435 = subckt_1633_sff1_x4.ckr
* NET 436 = subckt_1633_sff1_x4.nckr
* NET 437 = abc_11867_new_n873
* NET 449 = abc_11867_new_n868
* NET 451 = abc_11867_new_n864
* NET 452 = abc_11867_new_n874
* NET 460 = abc_11867_new_n865
* NET 464 = abc_11867_new_n876
* NET 466 = abc_11867_new_n875
* NET 472 = abc_11867_new_n863
* NET 482 = abc_11867_new_n870
* NET 487 = abc_11867_new_n428
* NET 489 = abc_11867_new_n608_hfns_2
* NET 494 = abc_11867_new_n475
* NET 499 = abc_11867_new_n471
* NET 508 = abc_11867_new_n431_hfns_2
* NET 510 = abc_11867_new_n431
* NET 663 = subckt_1744_sff1_x4.sff_s
* NET 664 = subckt_1744_sff1_x4.y
* NET 666 = subckt_1744_sff1_x4.sff_m
* NET 668 = subckt_1744_sff1_x4.u
* NET 669 = subckt_1744_sff1_x4.ckr
* NET 670 = subckt_1744_sff1_x4.nckr
* NET 672 = subckt_1654_sff1_x4.sff_s
* NET 673 = subckt_1654_sff1_x4.y
* NET 676 = subckt_1654_sff1_x4.sff_m
* NET 677 = subckt_1654_sff1_x4.ckr
* NET 678 = subckt_1654_sff1_x4.u
* NET 679 = subckt_1654_sff1_x4.nckr
* NET 680 = subckt_1652_sff1_x4.sff_s
* NET 683 = subckt_1652_sff1_x4.y
* NET 684 = subckt_1652_sff1_x4.sff_m
* NET 686 = subckt_1652_sff1_x4.u
* NET 687 = subckt_1652_sff1_x4.ckr
* NET 688 = subckt_1652_sff1_x4.nckr
* NET 690 = abc_11867_auto_rtlil_cc_2608_muxgate_11662
* NET 691 = mos6502_axys_2_5
* NET 692 = mos6502_axys_3_5
* NET 699 = subckt_1620_sff1_x4.sff_s
* NET 700 = subckt_1620_sff1_x4.y
* NET 701 = subckt_1620_sff1_x4.sff_m
* NET 703 = subckt_1620_sff1_x4.u
* NET 704 = subckt_1620_sff1_x4.ckr
* NET 705 = subckt_1620_sff1_x4.nckr
* NET 706 = mos6502_axys_2_1
* NET 708 = mos6502_axys_0_1
* NET 711 = mos6502_axys_3_1
* NET 712 = subckt_1618_sff1_x4.sff_s
* NET 714 = subckt_1618_sff1_x4.y
* NET 717 = subckt_1618_sff1_x4.sff_m
* NET 718 = subckt_1618_sff1_x4.u
* NET 719 = subckt_1618_sff1_x4.ckr
* NET 720 = subckt_1618_sff1_x4.nckr
* NET 722 = abc_11867_auto_rtlil_cc_2608_muxgate_11606
* NET 723 = mos6502_axys_2_0
* NET 724 = mos6502_axys_3_0
* NET 726 = mos6502_axys_0_0
* NET 729 = mos6502_axys_0_2
* NET 734 = subckt_1619_sff1_x4.sff_s
* NET 735 = subckt_1619_sff1_x4.y
* NET 736 = subckt_1619_sff1_x4.sff_m
* NET 739 = subckt_1619_sff1_x4.u
* NET 740 = subckt_1619_sff1_x4.ckr
* NET 741 = subckt_1619_sff1_x4.nckr
* NET 743 = abc_11867_auto_rtlil_cc_2608_muxgate_11624
* NET 745 = abc_11867_new_n867
* NET 747 = abc_11867_new_n862
* NET 750 = abc_11867_new_n859
* NET 752 = abc_11867_new_n1411
* NET 753 = abc_11867_new_n857
* NET 756 = abc_11867_new_n476
* NET 759 = abc_11867_new_n856
* NET 762 = abc_11867_new_n475_hfns_3
* NET 767 = abc_11867_new_n490
* NET 770 = abc_11867_new_n482
* NET 773 = abc_11867_new_n430
* NET 859 = subckt_1756_sff1_x4.sff_s
* NET 860 = subckt_1756_sff1_x4.sff_m
* NET 861 = subckt_1756_sff1_x4.y
* NET 863 = subckt_1756_sff1_x4.ckr
* NET 864 = subckt_1756_sff1_x4.u
* NET 865 = subckt_1756_sff1_x4.nckr
* NET 867 = abc_11867_auto_rtlil_cc_2608_muxgate_11860
* NET 876 = abc_11867_auto_rtlil_cc_2608_muxgate_11666
* NET 884 = subckt_1624_sff1_x4.sff_s
* NET 885 = subckt_1624_sff1_x4.sff_m
* NET 886 = subckt_1624_sff1_x4.y
* NET 888 = subckt_1624_sff1_x4.ckr
* NET 889 = subckt_1624_sff1_x4.u
* NET 890 = subckt_1624_sff1_x4.nckr
* NET 892 = abc_11867_auto_rtlil_cc_2608_muxgate_11618
* NET 901 = mos6502_axys_2_7
* NET 902 = mos6502_axys_3_7
* NET 915 = subckt_1636_sff1_x4.sff_s
* NET 916 = mos6502_axys_0_5
* NET 917 = subckt_1636_sff1_x4.sff_m
* NET 920 = subckt_1636_sff1_x4.y
* NET 925 = abc_11867_auto_rtlil_cc_2608_muxgate_11630
* NET 926 = subckt_1636_sff1_x4.u
* NET 928 = subckt_1636_sff1_x4.ckr
* NET 929 = subckt_1636_sff1_x4.nckr
* NET 934 = abc_11867_auto_rtlil_cc_2608_muxgate_11658
* NET 951 = mos6502_axys_2_3
* NET 959 = mos6502_axys_0_3
* NET 963 = abc_11867_auto_rtlil_cc_2608_muxgate_11626
* NET 969 = subckt_1640_sff1_x4.sff_s
* NET 970 = subckt_1640_sff1_x4.sff_m
* NET 974 = subckt_1640_sff1_x4.y
* NET 978 = subckt_1640_sff1_x4.u
* NET 980 = subckt_1640_sff1_x4.ckr
* NET 981 = subckt_1640_sff1_x4.nckr
* NET 983 = abc_11867_auto_rtlil_cc_2608_muxgate_11656
* NET 984 = mos6502_axys_2_2
* NET 992 = subckt_1651_sff1_x4.sff_s
* NET 997 = subckt_1651_sff1_x4.sff_m
* NET 998 = subckt_1651_sff1_x4.y
* NET 1002 = subckt_1651_sff1_x4.ckr
* NET 1003 = subckt_1651_sff1_x4.u
* NET 1004 = subckt_1651_sff1_x4.nckr
* NET 1005 = mos6502_axys_3_2
* NET 1008 = abc_11867_auto_rtlil_cc_2608_muxgate_11608
* NET 1020 = subckt_1621_sff1_x4.sff_s
* NET 1022 = subckt_1621_sff1_x4.sff_m
* NET 1023 = subckt_1621_sff1_x4.y
* NET 1025 = abc_11867_auto_rtlil_cc_2608_muxgate_11612
* NET 1026 = subckt_1621_sff1_x4.ckr
* NET 1027 = subckt_1621_sff1_x4.u
* NET 1028 = subckt_1621_sff1_x4.nckr
* NET 1035 = abc_11867_new_n858
* NET 1040 = abc_11867_new_n1424
* NET 1041 = abc_11867_new_n1410
* NET 1042 = abc_11867_new_n640
* NET 1055 = abc_11867_new_n380
* NET 1061 = abc_11867_new_n654
* NET 1067 = abc_11867_new_n471_hfns_3
* NET 1075 = abc_11867_new_n482_hfns_2
* NET 1079 = abc_11867_new_n473
* NET 1195 = subckt_1748_sff1_x4.sff_s
* NET 1196 = subckt_1748_sff1_x4.y
* NET 1198 = subckt_1748_sff1_x4.sff_m
* NET 1200 = subckt_1748_sff1_x4.u
* NET 1201 = subckt_1748_sff1_x4.ckr
* NET 1202 = subckt_1748_sff1_x4.nckr
* NET 1210 = abc_11867_new_n1906
* NET 1213 = subckt_1646_sff1_x4.sff_s
* NET 1214 = subckt_1646_sff1_x4.y
* NET 1216 = subckt_1646_sff1_x4.sff_m
* NET 1218 = subckt_1646_sff1_x4.ckr
* NET 1219 = subckt_1646_sff1_x4.u
* NET 1220 = subckt_1646_sff1_x4.nckr
* NET 1222 = subckt_1644_sff1_x4.sff_s
* NET 1224 = subckt_1644_sff1_x4.y
* NET 1225 = subckt_1644_sff1_x4.sff_m
* NET 1227 = subckt_1644_sff1_x4.u
* NET 1228 = subckt_1644_sff1_x4.ckr
* NET 1229 = subckt_1644_sff1_x4.nckr
* NET 1230 = abc_11867_auto_rtlil_cc_2608_muxgate_11646
* NET 1235 = abc_11867_auto_rtlil_cc_2608_muxgate_11650
* NET 1244 = abc_11867_auto_rtlil_cc_2608_muxgate_11610
* NET 1245 = mos6502_axys_3_3
* NET 1248 = abc_11867_new_n1103
* NET 1252 = subckt_1642_sff1_x4.sff_s
* NET 1253 = subckt_1642_sff1_x4.y
* NET 1256 = subckt_1642_sff1_x4.sff_m
* NET 1257 = subckt_1642_sff1_x4.u
* NET 1258 = subckt_1642_sff1_x4.nckr
* NET 1259 = subckt_1642_sff1_x4.ckr
* NET 1260 = abc_11867_auto_rtlil_cc_2608_muxgate_11638
* NET 1265 = abc_11867_auto_rtlil_cc_2608_muxgate_11660
* NET 1268 = abc_11867_new_n1166
* NET 1272 = subckt_1635_sff1_x4.sff_s
* NET 1274 = subckt_1635_sff1_x4.y
* NET 1276 = subckt_1635_sff1_x4.sff_m
* NET 1277 = subckt_1635_sff1_x4.u
* NET 1278 = subckt_1635_sff1_x4.ckr
* NET 1279 = subckt_1635_sff1_x4.nckr
* NET 1280 = abc_11867_auto_rtlil_cc_2608_muxgate_11628
* NET 1284 = abc_11867_new_n1148
* NET 1287 = abc_11867_new_n1421
* NET 1288 = abc_11867_new_n1426
* NET 1291 = abc_11867_new_n1409
* NET 1292 = abc_11867_new_n1407
* NET 1293 = abc_11867_new_n1412
* NET 1300 = abc_11867_new_n1423
* NET 1301 = abc_11867_new_n1425
* NET 1302 = abc_11867_new_n663
* NET 1308 = abc_11867_new_n426
* NET 1310 = abc_11867_new_n490_hfns_2
* NET 1314 = abc_11867_new_n430_hfns_2
* NET 1363 = subckt_1645_sff1_x4.sff_s
* NET 1365 = subckt_1645_sff1_x4.y
* NET 1369 = subckt_1645_sff1_x4.u
* NET 1370 = subckt_1645_sff1_x4.sff_m
* NET 1372 = subckt_1645_sff1_x4.ckr
* NET 1373 = subckt_1645_sff1_x4.nckr
* NET 1376 = subckt_1738_sff1_x4.sff_s
* NET 1380 = subckt_1738_sff1_x4.y
* NET 1382 = subckt_1738_sff1_x4.sff_m
* NET 1384 = subckt_1738_sff1_x4.ckr
* NET 1385 = subckt_1738_sff1_x4.u
* NET 1386 = subckt_1738_sff1_x4.nckr
* NET 1388 = abc_11867_auto_rtlil_cc_2608_muxgate_11648
* NET 1396 = mos6502_axys_1_6
* NET 1401 = abc_11867_new_n1030
* NET 1403 = mos6502_axys_1_7
* NET 1409 = abc_11867_new_n1022
* NET 1415 = subckt_1721_sff1_x4.sff_s
* NET 1416 = subckt_1721_sff1_x4.y
* NET 1418 = subckt_1721_sff1_x4.sff_m
* NET 1420 = subckt_1721_sff1_x4.u
* NET 1421 = subckt_1721_sff1_x4.ckr
* NET 1422 = subckt_1721_sff1_x4.nckr
* NET 1423 = mos6502_axys_0_7
* NET 1424 = subckt_1638_sff1_x4.sff_s
* NET 1427 = subckt_1638_sff1_x4.y
* NET 1430 = subckt_1638_sff1_x4.sff_m
* NET 1431 = abc_11867_auto_rtlil_cc_2608_muxgate_11634
* NET 1433 = subckt_1638_sff1_x4.u
* NET 1434 = subckt_1638_sff1_x4.nckr
* NET 1435 = subckt_1638_sff1_x4.ckr
* NET 1437 = abc_11867_auto_rtlil_cc_2608_muxgate_11642
* NET 1445 = subckt_1639_sff1_x4.sff_s
* NET 1449 = subckt_1639_sff1_x4.y
* NET 1451 = subckt_1639_sff1_x4.sff_m
* NET 1453 = subckt_1639_sff1_x4.ckr
* NET 1454 = subckt_1639_sff1_x4.u
* NET 1455 = subckt_1639_sff1_x4.nckr
* NET 1456 = mos6502_axys_1_1
* NET 1461 = abc_11867_auto_rtlil_cc_2608_muxgate_11636
* NET 1472 = subckt_1643_sff1_x4.sff_s
* NET 1474 = subckt_1643_sff1_x4.y
* NET 1477 = subckt_1643_sff1_x4.sff_m
* NET 1479 = subckt_1643_sff1_x4.u
* NET 1480 = subckt_1643_sff1_x4.ckr
* NET 1481 = subckt_1643_sff1_x4.nckr
* NET 1489 = abc_11867_new_n881
* NET 1490 = mos6502_axys_2_4
* NET 1493 = mos6502_axys_0_4
* NET 1494 = abc_11867_new_n882
* NET 1495 = abc_11867_new_n883
* NET 1496 = mos6502_axys_3_4
* NET 1500 = abc_11867_new_n1414
* NET 1501 = abc_11867_new_n1427
* NET 1504 = abc_11867_new_n1102
* NET 1519 = abc_11867_new_n1101
* NET 1520 = abc_11867_new_n959
* NET 1528 = abc_11867_new_n1413
* NET 1529 = abc_11867_new_n639
* NET 1537 = abc_11867_new_n1100
* NET 1542 = abc_11867_new_n766
* NET 1545 = abc_11867_new_n861
* NET 1552 = abc_11867_new_n656
* NET 1556 = abc_11867_new_n517
* NET 1573 = abc_11867_new_n606
* NET 1574 = abc_11867_new_n602
* NET 1575 = abc_11867_new_n599
* NET 1583 = abc_11867_new_n605
* NET 1601 = abc_11867_new_n426_hfns_2
* NET 1610 = abc_11867_new_n473_hfns_3
* NET 1793 = abc_11867_new_n1914
* NET 1796 = abc_11867_new_n1907
* NET 1801 = abc_11867_new_n1909
* NET 1802 = abc_11867_new_n1723
* NET 1804 = abc_11867_new_n1724
* NET 1805 = abc_11867_new_n1910
* NET 1806 = abc_11867_new_n1920
* NET 1807 = abc_11867_new_n1913
* NET 1810 = abc_11867_new_n1725
* NET 1813 = mos6502_axys_1_5
* NET 1815 = do[3]
* NET 1816 = abc_11867_auto_rtlil_cc_2608_muxgate_11790
* NET 1822 = abc_11867_new_n909
* NET 1824 = abc_11867_new_n999
* NET 1826 = mos6502_axys_1_3
* NET 1834 = abc_11867_new_n917
* NET 1837 = abc_11867_new_n914
* NET 1839 = abc_11867_auto_rtlil_cc_2608_muxgate_11644
* NET 1841 = abc_11867_new_n1157
* NET 1844 = mos6502_axys_1_4
* NET 1847 = subckt_1717_sff1_x4.sff_s
* NET 1848 = subckt_1717_sff1_x4.y
* NET 1851 = subckt_1717_sff1_x4.sff_m
* NET 1852 = subckt_1717_sff1_x4.u
* NET 1853 = subckt_1717_sff1_x4.ckr
* NET 1854 = subckt_1717_sff1_x4.nckr
* NET 1855 = abc_11867_new_n915
* NET 1857 = abc_11867_new_n916
* NET 1861 = abc_11867_new_n479
* NET 1862 = abc_11867_new_n383
* NET 1864 = abc_11867_new_n951
* NET 1865 = abc_11867_new_n1467
* NET 1866 = abc_11867_new_n1668
* NET 1867 = abc_11867_new_n1422
* NET 1868 = abc_11867_new_n1408
* NET 1870 = abc_11867_new_n1434
* NET 1871 = abc_11867_new_n855
* NET 1873 = abc_11867_new_n658
* NET 1874 = abc_11867_new_n966
* NET 1877 = we
* NET 1881 = abc_11867_new_n524
* NET 1884 = abc_11867_new_n690
* NET 1886 = abc_11867_new_n689
* NET 1890 = abc_11867_new_n641
* NET 1893 = abc_11867_new_n638
* NET 1898 = abc_11867_new_n659
* NET 1899 = abc_11867_new_n660
* NET 1958 = abc_11867_new_n1357
* NET 1964 = abc_11867_new_n1720
* NET 1973 = abc_11867_new_n1718
* NET 1991 = abc_11867_new_n1670
* NET 1993 = abc_11867_new_n1676
* NET 2000 = abc_11867_new_n1014
* NET 2003 = a[5]
* NET 2004 = abc_11867_new_n942
* NET 2006 = abc_11867_new_n943
* NET 2009 = subckt_1719_sff1_x4.sff_s
* NET 2011 = subckt_1719_sff1_x4.y
* NET 2014 = subckt_1719_sff1_x4.sff_m
* NET 2016 = subckt_1719_sff1_x4.u
* NET 2017 = subckt_1719_sff1_x4.ckr
* NET 2018 = subckt_1719_sff1_x4.nckr
* NET 2019 = abc_11867_auto_rtlil_cc_2608_muxgate_11786
* NET 2024 = a[3]
* NET 2035 = abc_11867_new_n983
* NET 2038 = mos6502_axys_1_2
* NET 2039 = subckt_1641_sff1_x4.sff_s
* NET 2043 = subckt_1641_sff1_x4.y
* NET 2046 = subckt_1641_sff1_x4.sff_m
* NET 2047 = abc_11867_auto_rtlil_cc_2608_muxgate_11640
* NET 2048 = subckt_1641_sff1_x4.ckr
* NET 2049 = subckt_1641_sff1_x4.u
* NET 2050 = subckt_1641_sff1_x4.nckr
* NET 2053 = subckt_1720_sff1_x4.sff_s
* NET 2054 = subckt_1720_sff1_x4.y
* NET 2057 = subckt_1720_sff1_x4.sff_m
* NET 2059 = subckt_1720_sff1_x4.u
* NET 2060 = subckt_1720_sff1_x4.ckr
* NET 2061 = subckt_1720_sff1_x4.nckr
* NET 2062 = abc_11867_auto_rtlil_cc_2608_muxgate_11788
* NET 2073 = a[4]
* NET 2074 = abc_11867_auto_rtlil_cc_2608_muxgate_11782
* NET 2081 = a[1]
* NET 2090 = abc_11867_new_n1420
* NET 2093 = abc_11867_new_n1417
* NET 2094 = abc_11867_new_n1415
* NET 2098 = abc_11867_new_n1418
* NET 2099 = abc_11867_new_n604
* NET 2102 = abc_11867_new_n1465
* NET 2104 = abc_11867_new_n1466
* NET 2105 = abc_11867_new_n1468
* NET 2109 = abc_11867_new_n965
* NET 2114 = abc_11867_new_n768
* NET 2119 = abc_11867_new_n1667
* NET 2121 = abc_11867_new_n598
* NET 2133 = abc_11867_new_n608_hfns_1
* NET 2138 = abc_11867_new_n509
* NET 2140 = abc_11867_new_n484
* NET 2147 = abc_11867_new_n774
* NET 2158 = abc_11867_new_n777
* NET 2165 = abc_11867_new_n613
* NET 2166 = abc_11867_new_n567
* NET 2167 = abc_11867_new_n603
* NET 2168 = abc_11867_new_n691
* NET 2172 = abc_11867_new_n580
* NET 2177 = abc_11867_new_n578
* NET 2203 = abc_11867_new_n725
* NET 2208 = abc_11867_new_n657
* NET 2209 = abc_11867_new_n652
* NET 2211 = abc_11867_new_n726
* NET 2212 = abc_11867_new_n729
* NET 2213 = abc_11867_new_n730
* NET 2216 = subckt_1630_sff1_x4.y
* NET 2217 = subckt_1630_sff1_x4.sff_s
* NET 2221 = subckt_1630_sff1_x4.sff_m
* NET 2222 = subckt_1630_sff1_x4.ckr
* NET 2223 = subckt_1630_sff1_x4.u
* NET 2224 = subckt_1630_sff1_x4.nckr
* NET 2373 = nmi
* NET 2375 = subckt_1749_sff1_x4.sff_s
* NET 2376 = subckt_1749_sff1_x4.y
* NET 2378 = subckt_1749_sff1_x4.sff_m
* NET 2380 = subckt_1749_sff1_x4.u
* NET 2381 = subckt_1749_sff1_x4.ckr
* NET 2382 = subckt_1749_sff1_x4.nckr
* NET 2384 = abc_11867_new_n1717
* NET 2385 = abc_11867_new_n1740
* NET 2393 = abc_11867_new_n1728
* NET 2401 = abc_11867_new_n1760
* NET 2403 = abc_11867_new_n1699
* NET 2406 = abc_11867_new_n1698
* NET 2412 = abc_11867_new_n927
* NET 2413 = abc_11867_new_n926
* NET 2415 = abc_11867_new_n895
* NET 2416 = do[1]
* NET 2417 = abc_11867_new_n935
* NET 2418 = abc_11867_new_n936
* NET 2420 = spare_buffer_19.q
* NET 2426 = abc_11867_new_n902
* NET 2427 = do[2]
* NET 2432 = mos6502_axys_1_0
* NET 2434 = abc_11867_new_n893
* NET 2435 = abc_11867_new_n894
* NET 2440 = subckt_1718_sff1_x4.sff_s
* NET 2441 = subckt_1718_sff1_x4.y
* NET 2442 = subckt_1718_sff1_x4.sff_m
* NET 2444 = subckt_1718_sff1_x4.u
* NET 2446 = clk_root_tr_2
* NET 2447 = subckt_1718_sff1_x4.nckr
* NET 2448 = subckt_1718_sff1_x4.ckr
* NET 2450 = abc_11867_new_n954
* NET 2452 = abc_11867_new_n953
* NET 2454 = abc_11867_new_n949
* NET 2456 = abc_11867_new_n1419
* NET 2459 = abc_11867_new_n1429
* NET 2462 = abc_11867_new_n1688
* NET 2464 = abc_11867_new_n1442
* NET 2466 = abc_11867_new_n1435
* NET 2469 = abc_11867_new_n1436
* NET 2470 = abc_11867_new_n625
* NET 2472 = abc_11867_new_n500
* NET 2473 = mos6502_state[5]
* NET 2474 = abc_11867_new_n429
* NET 2480 = abc_11867_new_n569
* NET 2481 = reset_root_tl_0
* NET 2483 = spare_buffer_14.q
* NET 2487 = abc_11867_new_n809
* NET 2490 = abc_11867_new_n829
* NET 2491 = abc_11867_new_n830
* NET 2492 = abc_11867_new_n832
* NET 2493 = abc_11867_new_n831
* NET 2495 = abc_11867_new_n775
* NET 2499 = abc_11867_new_n665
* NET 2500 = abc_11867_new_n664
* NET 2554 = subckt_1740_sff1_x4.y
* NET 2555 = subckt_1740_sff1_x4.sff_m
* NET 2572 = abc_11867_new_n583
* NET 2575 = abc_11867_new_n1437
* NET 2576 = abc_11867_new_n1441
* NET 2578 = abc_11867_new_n565
* NET 2581 = abc_11867_new_n581
* NET 2582 = abc_11867_new_n584
* NET 2589 = abc_11867_new_n644
* NET 2590 = abc_11867_new_n645
* NET 2592 = abc_11867_new_n823
* NET 2597 = abc_11867_new_n825
* NET 2601 = abc_11867_new_n525
* NET 2602 = abc_11867_new_n521
* NET 2609 = abc_11867_new_n1598
* NET 2610 = abc_11867_auto_rtlil_cc_2608_muxgate_11836
* NET 2614 = subckt_1740_sff1_x4.sff_s
* NET 2622 = subckt_1740_sff1_x4.nckr
* NET 2623 = subckt_1740_sff1_x4.ckr
* NET 2624 = subckt_1740_sff1_x4.u
* NET 2630 = abc_11867_new_n1745
* NET 2632 = abc_11867_new_n1739
* NET 2636 = abc_11867_new_n1908
* NET 2637 = abc_11867_new_n1746
* NET 2640 = abc_11867_new_n1738
* NET 2646 = abc_11867_new_n1697
* NET 2657 = abc_11867_new_n1696
* NET 2673 = clk_root_tr_1
* NET 2679 = abc_11867_new_n1912
* NET 2680 = abc_11867_new_n907
* NET 2681 = abc_11867_new_n908
* NET 2688 = abc_11867_new_n1669
* NET 2691 = abc_11867_new_n900
* NET 2692 = abc_11867_new_n901
* NET 2693 = abc_11867_new_n991
* NET 2697 = abc_11867_new_n954_hfns_2
* NET 2709 = abc_11867_auto_rtlil_cc_2608_muxgate_11784
* NET 2717 = a[2]
* NET 2727 = abc_11867_new_n1687
* NET 2728 = abc_11867_new_n530
* NET 2736 = abc_11867_new_n600
* NET 2741 = abc_11867_new_n563
* NET 2746 = abc_11867_new_n958
* NET 2750 = abc_11867_new_n1430
* NET 2752 = abc_11867_new_n1440
* NET 2753 = abc_11867_new_n850
* NET 2761 = abc_11867_new_n851
* NET 2763 = abc_11867_new_n853
* NET 2773 = spare_buffer_13.q
* NET 2776 = abc_11867_new_n776
* NET 2782 = abc_11867_new_n646
* NET 2788 = abc_11867_new_n738
* NET 2791 = abc_11867_new_n661
* NET 2792 = abc_11867_new_n666
* NET 2796 = abc_11867_new_n519
* NET 2799 = abc_11867_new_n527
* NET 2801 = abc_11867_new_n522
* NET 2956 = abc_11867_auto_rtlil_cc_2608_muxgate_11844
* NET 2957 = mos6502_alu_bi7
* NET 2962 = abc_11867_new_n1700
* NET 2964 = abc_11867_new_n1719
* NET 2965 = abc_11867_new_n1693
* NET 2967 = abc_11867_new_n1741
* NET 2968 = abc_11867_new_n1905
* NET 2971 = abc_11867_new_n1743
* NET 2973 = abc_11867_new_n1762
* NET 2974 = abc_11867_new_n1729
* NET 2982 = abc_11867_new_n1737
* NET 2984 = abc_11867_new_n1695
* NET 2985 = abc_11867_new_n1694
* NET 2986 = abc_11867_new_n1691
* NET 2989 = abc_11867_new_n1747
* NET 2996 = abc_11867_new_n1829
* NET 2997 = abc_11867_new_n1791
* NET 2998 = abc_11867_new_n1911
* NET 3000 = abc_11867_new_n1862
* NET 3003 = abc_11867_new_n885
* NET 3004 = abc_11867_new_n1816
* NET 3007 = abc_11867_new_n1817
* NET 3008 = abc_11867_new_n880
* NET 3009 = abc_11867_new_n884
* NET 3011 = abc_11867_new_n955
* NET 3012 = a[0]
* NET 3014 = subckt_1716_sff1_x4.sff_s
* NET 3015 = subckt_1716_sff1_x4.y
* NET 3018 = subckt_1716_sff1_x4.sff_m
* NET 3019 = abc_11867_auto_rtlil_cc_2608_muxgate_11780
* NET 3020 = subckt_1716_sff1_x4.u
* NET 3021 = subckt_1716_sff1_x4.ckr
* NET 3022 = subckt_1716_sff1_x4.nckr
* NET 3028 = abc_11867_new_n1039
* NET 3029 = abc_11867_new_n950
* NET 3032 = abc_11867_new_n952
* NET 3033 = abc_11867_new_n615
* NET 3035 = abc_11867_new_n1661
* NET 3036 = abc_11867_new_n1663
* NET 3037 = abc_11867_new_n1662
* NET 3040 = abc_11867_new_n579
* NET 3044 = abc_11867_new_n1689
* NET 3046 = abc_11867_new_n1439
* NET 3047 = abc_11867_new_n1438
* NET 3050 = abc_11867_new_n852
* NET 3057 = abc_11867_new_n614
* NET 3062 = abc_11867_new_n571
* NET 3063 = abc_11867_new_n566
* NET 3064 = abc_11867_new_n620
* NET 3065 = abc_11867_new_n616
* NET 3066 = abc_11867_new_n612
* NET 3068 = abc_11867_new_n810
* NET 3069 = abc_11867_new_n834
* NET 3070 = abc_11867_new_n572
* NET 3071 = abc_11867_new_n622
* NET 3072 = abc_11867_new_n817
* NET 3076 = abc_11867_new_n621
* NET 3077 = abc_11867_new_n607
* NET 3079 = abc_11867_new_n642
* NET 3081 = abc_11867_new_n650
* NET 3082 = abc_11867_new_n735
* NET 3084 = abc_11867_new_n736
* NET 3086 = abc_11867_new_n518
* NET 3088 = abc_11867_new_n516
* NET 3092 = mos6502_state[2]
* NET 3094 = subckt_1627_sff1_x4.sff_s
* NET 3095 = subckt_1627_sff1_x4.y
* NET 3096 = subckt_1627_sff1_x4.sff_m
* NET 3099 = subckt_1627_sff1_x4.ckr
* NET 3100 = subckt_1627_sff1_x4.u
* NET 3101 = subckt_1627_sff1_x4.nckr
* NET 3151 = abc_11867_new_n523
* NET 3152 = abc_11867_new_n1026
* NET 3155 = abc_11867_new_n1722
* NET 3158 = abc_11867_auto_rtlil_cc_2608_muxgate_11846
* NET 3160 = subckt_1757_sff1_x4.sff_s
* NET 3164 = subckt_1757_sff1_x4.y
* NET 3166 = subckt_1757_sff1_x4.sff_m
* NET 3167 = subckt_1757_sff1_x4.u
* NET 3168 = subckt_1757_sff1_x4.ckr
* NET 3169 = subckt_1757_sff1_x4.nckr
* NET 3175 = abc_11867_new_n1756
* NET 3179 = abc_11867_new_n1761
* NET 3183 = abc_11867_new_n1757
* NET 3188 = abc_11867_new_n1765
* NET 3193 = abc_11867_new_n1759
* NET 3198 = abc_11867_new_n1796
* NET 3202 = abc_11867_new_n1830
* NET 3213 = abc_11867_new_n1792
* NET 3219 = abc_11867_new_n1831
* NET 3230 = abc_11867_new_n1832
* NET 3236 = abc_11867_new_n1649
* NET 3242 = abc_11867_new_n1822
* NET 3246 = abc_11867_new_n1855
* NET 3263 = a[8]
* NET 3266 = subckt_1724_sff1_x4.y
* NET 3267 = subckt_1724_sff1_x4.sff_s
* NET 3270 = subckt_1724_sff1_x4.sff_m
* NET 3272 = abc_11867_auto_rtlil_cc_2608_muxgate_11796
* NET 3273 = subckt_1724_sff1_x4.ckr
* NET 3274 = subckt_1724_sff1_x4.u
* NET 3275 = subckt_1724_sff1_x4.nckr
* NET 3277 = abc_11867_new_n1104
* NET 3285 = abc_11867_new_n961
* NET 3288 = abc_11867_new_n1046
* NET 3292 = abc_11867_new_n1041
* NET 3295 = abc_11867_new_n1044
* NET 3306 = abc_11867_new_n956
* NET 3311 = abc_11867_new_n960
* NET 3322 = abc_11867_new_n957
* NET 3331 = abc_11867_new_n1431
* NET 3337 = abc_11867_new_n1433
* NET 3338 = abc_11867_new_n1432
* NET 3349 = abc_11867_new_n724
* NET 3355 = abc_11867_new_n649
* NET 3370 = abc_11867_new_n556
* NET 3375 = abc_11867_new_n835
* NET 3377 = abc_11867_new_n833
* NET 3379 = abc_11867_new_n505
* NET 3382 = abc_11867_new_n824
* NET 3391 = abc_11867_new_n800
* NET 3396 = abc_11867_new_n526
* NET 3402 = abc_11867_new_n651
* NET 3403 = abc_11867_new_n667
* NET 3410 = abc_11867_new_n485
* NET 3413 = mos6502_state[4]
* NET 3416 = subckt_1629_sff1_x4.y
* NET 3417 = subckt_1629_sff1_x4.sff_s
* NET 3420 = subckt_1629_sff1_x4.sff_m
* NET 3422 = subckt_1629_sff1_x4.ckr
* NET 3423 = subckt_1629_sff1_x4.u
* NET 3424 = subckt_1629_sff1_x4.nckr
* NET 3425 = do[0]
* NET 3606 = abc_11867_new_n1763
* NET 3607 = abc_11867_new_n1767
* NET 3610 = abc_11867_new_n1768
* NET 3611 = abc_11867_new_n1904
* NET 3612 = abc_11867_new_n1902
* NET 3615 = abc_11867_new_n1716
* NET 3617 = abc_11867_new_n1766
* NET 3618 = abc_11867_new_n1734
* NET 3621 = abc_11867_new_n1735
* NET 3625 = abc_11867_new_n1736
* NET 3626 = abc_11867_new_n1758
* NET 3628 = abc_11867_new_n1744
* NET 3630 = abc_11867_new_n1754
* NET 3632 = abc_11867_new_n1683
* NET 3635 = abc_11867_new_n1750
* NET 3637 = abc_11867_new_n1783
* NET 3646 = abc_11867_new_n1834
* NET 3647 = abc_11867_new_n1833
* NET 3651 = abc_11867_new_n1835
* NET 3652 = abc_11867_new_n1837
* NET 3654 = abc_11867_new_n1821
* NET 3658 = abc_11867_new_n1854
* NET 3664 = abc_11867_new_n1846
* NET 3668 = abc_11867_new_n1876
* NET 3675 = abc_11867_new_n1925
* NET 3677 = abc_11867_new_n1926
* NET 3679 = subckt_1750_sff1_x4.sff_s
* NET 3680 = subckt_1750_sff1_x4.y
* NET 3683 = subckt_1750_sff1_x4.sff_m
* NET 3684 = abc_11867_auto_rtlil_cc_2608_muxgate_11848
* NET 3685 = subckt_1750_sff1_x4.u
* NET 3686 = subckt_1750_sff1_x4.ckr
* NET 3687 = subckt_1750_sff1_x4.nckr
* NET 3688 = abc_11867_new_n1666
* NET 3693 = abc_11867_new_n972
* NET 3694 = abc_11867_new_n1042
* NET 3695 = abc_11867_new_n1659
* NET 3698 = abc_11867_new_n491
* NET 3703 = abc_11867_new_n382
* NET 3704 = abc_11867_new_n483
* NET 3706 = abc_11867_new_n381
* NET 3709 = abc_11867_new_n493
* NET 3710 = abc_11867_new_n767
* NET 3712 = abc_11867_new_n769
* NET 3714 = abc_11867_new_n515
* NET 3716 = abc_11867_new_n591
* NET 3718 = abc_11867_new_n590
* NET 3719 = abc_11867_new_n550
* NET 3721 = abc_11867_new_n836
* NET 3722 = abc_11867_new_n655
* NET 3723 = abc_11867_new_n506
* NET 3726 = abc_11867_new_n555
* NET 3728 = abc_11867_new_n573
* NET 3734 = abc_11867_new_n508
* NET 3735 = abc_11867_new_n653
* NET 3738 = abc_11867_new_n551
* NET 3739 = abc_11867_new_n549
* NET 3744 = subckt_1625_sff1_x4.sff_s
* NET 3745 = subckt_1625_sff1_x4.y
* NET 3748 = subckt_1625_sff1_x4.sff_m
* NET 3749 = subckt_1625_sff1_x4.u
* NET 3750 = subckt_1625_sff1_x4.ckr
* NET 3751 = subckt_1625_sff1_x4.nckr
* NET 3804 = abc_11867_new_n374
* NET 3814 = abc_11867_new_n1903
* NET 3817 = abc_11867_new_n1692
* NET 3822 = abc_11867_new_n1713
* NET 3830 = abc_11867_new_n1742
* NET 3832 = abc_11867_new_n1028
* NET 3833 = abc_11867_new_n1027
* NET 3837 = abc_11867_new_n1732
* NET 3844 = abc_11867_new_n1751
* NET 3849 = abc_11867_new_n1784
* NET 3860 = abc_11867_new_n1685
* NET 3871 = abc_11867_new_n1782
* NET 3872 = abc_11867_new_n1841
* NET 3875 = abc_11867_new_n1889
* NET 3879 = abc_11867_new_n1825
* NET 3884 = abc_11867_new_n1828
* NET 3889 = abc_11867_new_n1827
* NET 3890 = abc_11867_new_n1856
* NET 3893 = abc_11867_new_n1853
* NET 3905 = abc_11867_new_n1875
* NET 3917 = abc_11867_new_n1877
* NET 3922 = abc_11867_new_n1881
* NET 3925 = abc_11867_new_n1883
* NET 3928 = abc_11867_new_n1874
* NET 3938 = abc_11867_new_n1878
* NET 3941 = abc_11867_new_n1880
* NET 3945 = abc_11867_new_n1884
* NET 3952 = abc_11867_new_n1924
* NET 3956 = abc_11867_new_n1045
* NET 3958 = abc_11867_new_n1660
* NET 3959 = abc_11867_new_n1664
* NET 3961 = abc_11867_new_n967
* NET 3962 = abc_11867_new_n962
* NET 3967 = abc_11867_new_n499
* NET 3969 = abc_11867_new_n486
* NET 3974 = abc_11867_new_n575
* NET 3976 = abc_11867_new_n487
* NET 3982 = abc_11867_new_n770
* NET 3983 = abc_11867_new_n1428
* NET 3993 = abc_11867_new_n488
* NET 3994 = abc_11867_new_n477
* NET 4000 = abc_11867_new_n771
* NET 4003 = abc_11867_new_n701
* NET 4005 = abc_11867_new_n700
* NET 4010 = abc_11867_new_n495
* NET 4012 = abc_11867_new_n570
* NET 4013 = abc_11867_new_n806
* NET 4014 = abc_11867_new_n427
* NET 4023 = abc_11867_new_n560
* NET 4029 = abc_11867_new_n561
* NET 4030 = abc_11867_new_n763
* NET 4031 = abc_11867_new_n662
* NET 4036 = abc_11867_new_n574
* NET 4037 = abc_11867_new_n592
* NET 4038 = abc_11867_new_n562
* NET 4042 = abc_11867_new_n635
* NET 4043 = abc_11867_new_n634
* NET 4047 = abc_11867_new_n797
* NET 4048 = abc_11867_new_n798
* NET 4054 = abc_11867_new_n668
* NET 4057 = abc_11867_new_n623
* NET 4058 = abc_11867_new_n593
* NET 4063 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[5]
* NET 4064 = abc_11867_new_n837
* NET 4066 = mos6502_state[0]
* NET 4070 = mos6502_state[1]
* NET 4073 = subckt_1626_sff1_x4.y
* NET 4074 = subckt_1626_sff1_x4.sff_s
* NET 4078 = subckt_1626_sff1_x4.sff_m
* NET 4079 = subckt_1626_sff1_x4.ckr
* NET 4080 = subckt_1626_sff1_x4.u
* NET 4081 = subckt_1626_sff1_x4.nckr
* NET 4142 = abc_11867_new_n1665
* NET 4183 = abc_11867_new_n632
* NET 4240 = a[7]
* NET 4250 = abc_11867_new_n733
* NET 4254 = mos6502_pc[12]
* NET 4255 = abc_11867_new_n1024
* NET 4258 = subckt_1755_sff1_x4.sff_s
* NET 4260 = subckt_1755_sff1_x4.ckr
* NET 4261 = subckt_1755_sff1_x4.y
* NET 4262 = subckt_1755_sff1_x4.sff_m
* NET 4265 = subckt_1755_sff1_x4.u
* NET 4268 = subckt_1755_sff1_x4.nckr
* NET 4272 = abc_11867_new_n1785
* NET 4274 = abc_11867_new_n1764
* NET 4275 = abc_11867_new_n1786
* NET 4277 = abc_11867_new_n1789
* NET 4279 = abc_11867_new_n1788
* NET 4281 = abc_11867_new_n1779
* NET 4285 = abc_11867_new_n1836
* NET 4286 = abc_11867_new_n1840
* NET 4288 = abc_11867_new_n1839
* NET 4290 = abc_11867_new_n1838
* NET 4291 = abc_11867_new_n1826
* NET 4295 = abc_11867_new_n1861
* NET 4298 = abc_11867_new_n1886
* NET 4301 = abc_11867_new_n1859
* NET 4304 = abc_11867_new_n1851
* NET 4305 = abc_11867_new_n1863
* NET 4306 = abc_11867_new_n1867
* NET 4307 = abc_11867_new_n1879
* NET 4311 = abc_11867_new_n1842
* NET 4312 = abc_11867_new_n1845
* NET 4314 = abc_11867_new_n1710
* NET 4316 = abc_11867_new_n1870
* NET 4318 = abc_11867_new_n1871
* NET 4320 = abc_11867_new_n1872
* NET 4322 = abc_11867_new_n1873
* NET 4323 = abc_11867_new_n1869
* NET 4325 = abc_11867_new_n848
* NET 4327 = abc_11867_new_n503
* NET 4333 = abc_11867_new_n778
* NET 4335 = abc_11867_new_n588
* NET 4342 = abc_11867_new_n779
* NET 4344 = abc_11867_new_n772
* NET 4347 = abc_11867_new_n504
* NET 4348 = abc_11867_new_n510
* NET 4349 = abc_11867_new_n597
* NET 4352 = abc_11867_new_n428_hfns_5
* NET 4354 = abc_11867_new_n811
* NET 4356 = abc_11867_new_n485_hfns_4
* NET 4359 = abc_11867_new_n528
* NET 4361 = abc_11867_new_n737
* NET 4363 = abc_11867_new_n669
* NET 4364 = abc_11867_new_n554
* NET 4368 = abc_11867_new_n790
* NET 4369 = abc_11867_new_n781
* NET 4370 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[2]
* NET 4374 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[1]
* NET 4405 = subckt_1723_sff1_x4.y
* NET 4407 = subckt_1723_sff1_x4.sff_m
* NET 4410 = abc_11867_new_n1684
* NET 4436 = subckt_1685_sff1_x4.y
* NET 4438 = subckt_1685_sff1_x4.sff_m
* NET 4439 = abc_11867_new_n773
* NET 4450 = abc_11867_new_n511
* NET 4451 = abc_11867_new_n489
* NET 4452 = abc_11867_new_n502
* NET 4453 = abc_11867_new_n711
* NET 4463 = abc_11867_new_n839
* NET 4465 = abc_11867_new_n780
* NET 4467 = abc_11867_new_n529
* NET 4472 = abc_11867_new_n816
* NET 4476 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[0]
* NET 4478 = abc_11867_new_n815
* NET 4481 = subckt_1628_sff1_x4.y
* NET 4484 = subckt_1628_sff1_x4.sff_m
* NET 4488 = abc_11867_new_n1918
* NET 4489 = abc_11867_new_n1917
* NET 4494 = subckt_1723_sff1_x4.sff_s
* NET 4496 = abc_11867_auto_rtlil_cc_2608_muxgate_11794
* NET 4497 = subckt_1723_sff1_x4.ckr
* NET 4498 = subckt_1723_sff1_x4.u
* NET 4499 = subckt_1723_sff1_x4.nckr
* NET 4500 = abc_11867_new_n1790
* NET 4501 = abc_11867_new_n1901
* NET 4508 = abc_11867_new_n1733
* NET 4524 = a[6]
* NET 4530 = abc_11867_new_n1780
* NET 4535 = abc_11867_new_n1781
* NET 4539 = abc_11867_new_n1888
* NET 4543 = abc_11867_new_n1890
* NET 4553 = abc_11867_new_n1680
* NET 4555 = abc_11867_new_n1804
* NET 4567 = abc_11867_new_n1730
* NET 4584 = abc_11867_new_n1850
* NET 4587 = abc_11867_new_n1852
* NET 4602 = abc_11867_new_n1882
* NET 4617 = abc_11867_new_n1682
* NET 4628 = abc_11867_new_n1679
* NET 4631 = abc_11867_new_n1708
* NET 4640 = abc_11867_new_n1678
* NET 4653 = abc_11867_new_n636
* NET 4654 = abc_11867_new_n474
* NET 4658 = abc_11867_new_n520
* NET 4665 = abc_11867_new_n643
* NET 4666 = abc_11867_new_n637
* NET 4672 = subckt_1685_sff1_x4.sff_s
* NET 4673 = mos6502_src_reg[0]
* NET 4675 = subckt_1685_sff1_x4.ckr
* NET 4676 = subckt_1685_sff1_x4.u
* NET 4677 = subckt_1685_sff1_x4.nckr
* NET 4679 = abc_11867_new_n709
* NET 4680 = abc_11867_new_n386
* NET 4684 = abc_11867_new_n869
* NET 4694 = abc_11867_new_n596
* NET 4700 = abc_11867_new_n803
* NET 4701 = abc_11867_new_n807
* NET 4708 = abc_11867_new_n512
* NET 4710 = abc_11867_new_n513
* NET 4717 = abc_11867_new_n552
* NET 4720 = abc_11867_new_n553
* NET 4723 = abc_11867_new_n820
* NET 4724 = subckt_1628_sff1_x4.sff_s
* NET 4726 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[3]
* NET 4727 = subckt_1628_sff1_x4.u
* NET 4728 = subckt_1628_sff1_x4.ckr
* NET 4729 = subckt_1628_sff1_x4.nckr
* NET 4880 = abc_11867_new_n1549
* NET 4881 = abc_11867_auto_rtlil_cc_2608_muxgate_11828
* NET 4885 = abc_11867_auto_rtlil_cc_2608_muxgate_11826
* NET 4887 = subckt_1722_sff1_x4.sff_s
* NET 4888 = subckt_1722_sff1_x4.y
* NET 4890 = subckt_1722_sff1_x4.sff_m
* NET 4892 = abc_11867_auto_rtlil_cc_2608_muxgate_11792
* NET 4893 = subckt_1722_sff1_x4.u
* NET 4894 = subckt_1722_sff1_x4.ckr
* NET 4895 = subckt_1722_sff1_x4.nckr
* NET 4896 = subckt_1754_sff1_x4.sff_s
* NET 4899 = subckt_1754_sff1_x4.y
* NET 4900 = subckt_1754_sff1_x4.sff_m
* NET 4902 = subckt_1754_sff1_x4.u
* NET 4903 = subckt_1754_sff1_x4.nckr
* NET 4904 = subckt_1754_sff1_x4.ckr
* NET 4905 = abc_11867_new_n1140
* NET 4910 = abc_11867_new_n1146
* NET 4915 = abc_11867_new_n1686
* NET 4916 = abc_11867_new_n1787
* NET 4919 = abc_11867_new_n1806
* NET 4925 = abc_11867_new_n1712
* NET 4926 = abc_11867_new_n1715
* NET 4929 = abc_11867_new_n1650
* NET 4932 = abc_11867_new_n1805
* NET 4936 = abc_11867_new_n1797
* NET 4939 = abc_11867_new_n1731
* NET 4940 = abc_11867_new_n1857
* NET 4942 = abc_11867_new_n1858
* NET 4943 = abc_11867_new_n1860
* NET 4944 = abc_11867_new_n1849
* NET 4948 = abc_11867_new_n1885
* NET 4950 = abc_11867_new_n1887
* NET 4952 = abc_11867_new_n1701
* NET 4954 = abc_11867_new_n1702
* NET 4955 = abc_11867_new_n847
* NET 4956 = abc_11867_new_n845
* NET 4959 = abc_11867_new_n1709
* NET 4960 = abc_11867_new_n1707
* NET 4966 = subckt_1715_sff1_x4.sff_s
* NET 4968 = subckt_1715_sff1_x4.y
* NET 4969 = abc_11867_auto_rtlil_cc_2608_muxgate_11778
* NET 4971 = subckt_1715_sff1_x4.sff_m
* NET 4972 = subckt_1715_sff1_x4.u
* NET 4973 = subckt_1715_sff1_x4.nckr
* NET 4974 = subckt_1715_sff1_x4.ckr
* NET 4975 = abc_11867_new_n356
* NET 4976 = abc_11867_new_n1654
* NET 4979 = abc_11867_new_n1658
* NET 4981 = abc_11867_new_n765
* NET 4983 = abc_11867_new_n1647
* NET 4984 = abc_11867_new_n1653
* NET 4986 = abc_11867_new_n1652
* NET 4991 = abc_11867_new_n740
* NET 4995 = abc_11867_new_n866
* NET 4996 = abc_11867_new_n501
* NET 4997 = abc_11867_new_n713
* NET 4998 = abc_11867_new_n710
* NET 5001 = abc_11867_new_n712
* NET 5002 = abc_11867_new_n714
* NET 5008 = abc_11867_new_n703
* NET 5009 = abc_11867_new_n702
* NET 5012 = abc_11867_new_n589
* NET 5014 = abc_11867_new_n808
* NET 5015 = abc_11867_new_n826
* NET 5017 = abc_11867_new_n789
* NET 5018 = abc_11867_new_n788
* NET 5023 = abc_11867_new_n716
* NET 5024 = abc_11867_new_n715
* NET 5029 = abc_11867_new_n818
* NET 5032 = abc_11867_new_n819
* NET 5033 = abc_11867_new_n827
* NET 5034 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[4]
* NET 5035 = abc_11867_new_n478
* NET 5037 = abc_11867_new_n814
* NET 5038 = abc_11867_new_n792
* NET 5040 = abc_11867_new_n802
* NET 5075 = subckt_1759_sff1_x4.sff_s
* NET 5076 = subckt_1759_sff1_x4.y
* NET 5080 = subckt_1759_sff1_x4.sff_m
* NET 5081 = subckt_1759_sff1_x4.u
* NET 5083 = clk_root_tr_0
* NET 5084 = subckt_1759_sff1_x4.nckr
* NET 5085 = subckt_1759_sff1_x4.ckr
* NET 5086 = abc_11867_new_n1036
* NET 5091 = abc_11867_new_n1031
* NET 5093 = abc_11867_new_n355
* NET 5094 = abc_11867_new_n1932
* NET 5097 = abc_11867_auto_rtlil_cc_2608_muxgate_11856
* NET 5098 = abc_11867_new_n1900
* NET 5100 = abc_11867_new_n1933
* NET 5103 = abc_11867_new_n1023
* NET 5105 = abc_11867_new_n1752
* NET 5119 = abc_11867_new_n1753
* NET 5123 = abc_11867_new_n1755
* NET 5124 = abc_11867_new_n1711
* NET 5128 = abc_11867_new_n1809
* NET 5131 = abc_11867_new_n1714
* NET 5132 = abc_11867_new_n1810
* NET 5140 = abc_11867_new_n1801
* NET 5142 = abc_11867_new_n1921
* NET 5143 = abc_11867_new_n1919
* NET 5144 = abc_11867_new_n1922
* NET 5148 = abc_11867_new_n1803
* NET 5150 = abc_11867_new_n1774
* NET 5153 = abc_11867_new_n1824
* NET 5159 = abc_11867_new_n1848
* NET 5162 = abc_11867_new_n1539
* NET 5165 = abc_11867_new_n1865
* NET 5168 = abc_11867_new_n968
* NET 5175 = abc_11867_new_n1703
* NET 5177 = abc_11867_new_n841
* NET 5181 = abc_11867_new_n1648
* NET 5183 = abc_11867_new_n1704
* NET 5185 = abc_11867_new_n1706
* NET 5191 = mos6502_backwards
* NET 5194 = abc_11867_new_n1705
* NET 5199 = reset
* NET 5202 = abc_11867_new_n846
* NET 5207 = abc_11867_new_n974
* NET 5214 = abc_11867_new_n969
* NET 5216 = abc_11867_new_n1657
* NET 5220 = abc_11867_new_n1655
* NET 5226 = abc_11867_new_n564
* NET 5229 = abc_11867_new_n624
* NET 5240 = abc_11867_new_n1651
* NET 5253 = abc_11867_new_n494
* NET 5255 = subckt_1684_sff1_x4.sff_s
* NET 5256 = subckt_1684_sff1_x4.y
* NET 5261 = subckt_1684_sff1_x4.sff_m
* NET 5262 = clk_root_tl_0
* NET 5263 = subckt_1684_sff1_x4.ckr
* NET 5264 = subckt_1684_sff1_x4.u
* NET 5265 = subckt_1684_sff1_x4.nckr
* NET 5269 = abc_11867_new_n497
* NET 5271 = abc_11867_new_n784
* NET 5273 = abc_11867_new_n568
* NET 5275 = abc_11867_new_n594
* NET 5279 = abc_11867_new_n692
* NET 5283 = abc_11867_new_n693
* NET 5286 = abc_11867_new_n694
* NET 5288 = abc_11867_new_n787
* NET 5292 = abc_11867_new_n739
* NET 5293 = abc_11867_new_n426_hfns_0
* NET 5295 = abc_11867_new_n732
* NET 5297 = abc_11867_new_n762
* NET 5302 = abc_11867_new_n731
* NET 5304 = abc_11867_new_n838
* NET 5307 = abc_11867_new_n785
* NET 5309 = abc_11867_new_n786
* NET 5312 = abc_11867_new_n813
* NET 5313 = abc_11867_new_n812
* NET 5320 = abc_11867_new_n801
* NET 5321 = abc_11867_new_n799
* NET 5487 = abc_11867_auto_rtlil_cc_2608_muxgate_11866
* NET 5488 = mos6502_alu_ai7
* NET 5490 = abc_11867_new_n1677
* NET 5494 = abc_11867_auto_rtlil_cc_2608_muxgate_11858
* NET 5496 = abc_11867_new_n1916
* NET 5500 = abc_11867_new_n1136
* NET 5501 = abc_11867_new_n1020
* NET 5503 = abc_11867_new_n1931
* NET 5504 = abc_11867_new_n1015
* NET 5510 = abc_11867_new_n1132
* NET 5518 = abc_11867_new_n1807
* NET 5519 = abc_11867_new_n1777
* NET 5521 = abc_11867_new_n1778
* NET 5522 = abc_11867_new_n1776
* NET 5523 = abc_11867_new_n1800
* NET 5525 = abc_11867_new_n1775
* NET 5527 = abc_11867_new_n1773
* NET 5528 = abc_11867_new_n1769
* NET 5531 = abc_11867_new_n1110
* NET 5535 = abc_11867_new_n1819
* NET 5539 = abc_11867_new_n1868
* NET 5541 = abc_11867_new_n353
* NET 5544 = abc_11867_new_n1126
* NET 5550 = abc_11867_new_n1043
* NET 5552 = abc_11867_new_n727
* NET 5554 = clk
* NET 5556 = abc_11867_new_n849
* NET 5557 = abc_11867_new_n918
* NET 5561 = abc_11867_new_n919
* NET 5562 = abc_11867_new_n357
* NET 5564 = abc_11867_new_n347
* NET 5565 = abc_11867_new_n1656
* NET 5568 = subckt_1675_sff1_x4.sff_s
* NET 5569 = subckt_1675_sff1_x4.y
* NET 5571 = subckt_1675_sff1_x4.sff_m
* NET 5573 = subckt_1675_sff1_x4.u
* NET 5574 = subckt_1675_sff1_x4.ckr
* NET 5575 = subckt_1675_sff1_x4.nckr
* NET 5577 = abc_11867_new_n514
* NET 5579 = abc_11867_new_n496
* NET 5580 = abc_11867_new_n498
* NET 5581 = abc_11867_new_n514_hfns_2
* NET 5583 = abc_11867_new_n485_hfns_3
* NET 5586 = subckt_1687_sff1_x4.sff_s
* NET 5587 = subckt_1687_sff1_x4.y
* NET 5589 = subckt_1687_sff1_x4.sff_m
* NET 5591 = subckt_1687_sff1_x4.u
* NET 5592 = subckt_1687_sff1_x4.ckr
* NET 5593 = abc_11867_new_n492
* NET 5594 = subckt_1687_sff1_x4.nckr
* NET 5599 = abc_11867_new_n471_hfns_1
* NET 5600 = abc_11867_new_n482_hfns_0
* NET 5601 = abc_11867_new_n699
* NET 5603 = abc_11867_new_n704
* NET 5606 = abc_11867_new_n822
* NET 5607 = abc_11867_new_n426_hfns_1
* NET 5608 = abc_11867_new_n478_hfns_3
* NET 5610 = abc_11867_new_n683
* NET 5611 = rdy
* NET 5655 = subckt_1741_sff1_x4.sff_s
* NET 5657 = subckt_1741_sff1_x4.y
* NET 5660 = subckt_1741_sff1_x4.sff_m
* NET 5662 = subckt_1741_sff1_x4.u
* NET 5663 = subckt_1741_sff1_x4.ckr
* NET 5664 = subckt_1741_sff1_x4.nckr
* NET 5665 = abc_11867_new_n1032
* NET 5667 = abc_11867_new_n1035
* NET 5670 = abc_11867_new_n1034
* NET 5671 = abc_11867_new_n375
* NET 5672 = abc_11867_new_n1005
* NET 5681 = abc_11867_new_n1808
* NET 5684 = abc_11867_new_n1811
* NET 5693 = abc_11867_new_n1815
* NET 5698 = abc_11867_new_n1893
* NET 5702 = abc_11867_new_n1812
* NET 5703 = abc_11867_new_n1898
* NET 5704 = abc_11867_new_n1813
* NET 5707 = abc_11867_new_n1124
* NET 5718 = abc_11867_new_n1823
* NET 5719 = abc_11867_new_n473_hfns_2
* NET 5726 = abc_11867_new_n1795
* NET 5727 = abc_11867_new_n1416
* NET 5728 = abc_11867_new_n1690
* NET 5732 = abc_11867_new_n1118
* NET 5736 = abc_11867_new_n610
* NET 5743 = abc_11867_new_n1820
* NET 5746 = abc_11867_new_n997
* NET 5748 = abc_11867_new_n928
* NET 5753 = abc_11867_new_n1866
* NET 5755 = abc_11867_new_n933
* NET 5756 = abc_11867_new_n931
* NET 5757 = abc_11867_new_n932
* NET 5764 = abc_11867_new_n968_hfns_2
* NET 5766 = abc_11867_new_n1012
* NET 5770 = abc_11867_new_n920
* NET 5771 = abc_11867_new_n843
* NET 5774 = abc_11867_new_n921
* NET 5776 = abc_11867_new_n924
* NET 5777 = abc_11867_new_n923
* NET 5782 = abc_11867_new_n922
* NET 5801 = abc_11867_new_n1497
* NET 5809 = abc_11867_new_n728
* NET 5811 = irq
* NET 5816 = abc_11867_new_n1392
* NET 5818 = abc_11867_new_n1337
* NET 5824 = subckt_1709_sff1_x4.sff_s
* NET 5826 = subckt_1709_sff1_x4.y
* NET 5829 = abc_11867_auto_rtlil_cc_2608_muxgate_11768
* NET 5831 = subckt_1709_sff1_x4.u
* NET 5832 = subckt_1709_sff1_x4.sff_m
* NET 5833 = subckt_1709_sff1_x4.ckr
* NET 5834 = subckt_1709_sff1_x4.nckr
* NET 5837 = abc_11867_new_n385
* NET 5841 = abc_11867_auto_rtlil_cc_2608_muxgate_11708
* NET 5842 = mos6502_shift_right
* NET 5851 = abc_11867_new_n346
* NET 5853 = subckt_1680_sff1_x4.sff_s
* NET 5857 = subckt_1680_sff1_x4.y
* NET 5858 = subckt_1680_sff1_x4.sff_m
* NET 5860 = subckt_1680_sff1_x4.ckr
* NET 5861 = subckt_1680_sff1_x4.u
* NET 5862 = subckt_1680_sff1_x4.nckr
* NET 5863 = mos6502_index_y
* NET 5866 = abc_11867_auto_rtlil_cc_2608_muxgate_11728
* NET 5873 = abc_11867_new_n805
* NET 5878 = abc_11867_new_n783
* NET 5890 = abc_11867_new_n684
* NET 5891 = abc_11867_new_n686
* NET 5897 = abc_11867_new_n782
* NET 5898 = abc_11867_new_n475_hfns_0
* NET 5901 = abc_11867_new_n514_hfns_0
* NET 5906 = abc_11867_new_n717
* NET 5908 = abc_11867_new_n720
* NET 5911 = abc_11867_new_n475_hfns_1
* NET 5918 = abc_11867_new_n471_hfns_0
* NET 5919 = abc_11867_new_n608_hfns_0
* NET 5926 = abc_11867_new_n548
* NET 5927 = abc_11867_new_n531
* NET 5931 = abc_11867_new_n796
* NET 5933 = abc_11867_new_n794
* NET 5934 = abc_11867_new_n795
* NET 6105 = abc_11867_new_n1134
* NET 6106 = abc_11867_new_n1139
* NET 6108 = abc_11867_new_n1000
* NET 6109 = abc_11867_new_n351
* NET 6116 = abc_11867_new_n354
* NET 6117 = abc_11867_new_n1123
* NET 6119 = abc_11867_new_n1897
* NET 6121 = abc_11867_new_n1033
* NET 6127 = abc_11867_new_n1847
* NET 6128 = abc_11867_new_n1802
* NET 6130 = abc_11867_new_n891
* NET 6131 = abc_11867_new_n992
* NET 6132 = abc_11867_new_n954_hfns_1
* NET 6137 = abc_11867_new_n1038
* NET 6140 = abc_11867_new_n905
* NET 6141 = abc_11867_new_n930
* NET 6142 = abc_11867_new_n1007
* NET 6150 = abc_11867_new_n1399
* NET 6151 = abc_11867_new_n1366
* NET 6152 = abc_11867_new_n1368
* NET 6163 = mos6502_dst_reg[0]
* NET 6164 = abc_11867_auto_rtlil_cc_2608_muxgate_11734
* NET 6171 = abc_11867_new_n630
* NET 6173 = abc_11867_new_n633
* NET 6175 = abc_11867_new_n679
* NET 6176 = abc_11867_new_n719
* NET 6177 = abc_11867_new_n682
* NET 6179 = abc_11867_new_n723
* NET 6180 = abc_11867_new_n678
* NET 6182 = abc_11867_new_n793
* NET 6183 = subckt_1745_sff1_x4.sff_s
* NET 6184 = subckt_1745_sff1_x4.y
* NET 6185 = subckt_1745_sff1_x4.sff_m
* NET 6186 = subckt_1745_sff1_x4.u
* NET 6187 = subckt_1745_sff1_x4.ckr
* NET 6188 = subckt_1745_sff1_x4.nckr
* NET 6192 = abc_11867_new_n1138
* NET 6194 = subckt_1615_nmx2_x1.q
* NET 6195 = abc_11867_new_n1899
* NET 6200 = abc_11867_new_n1814
* NET 6201 = abc_11867_new_n1891
* NET 6205 = abc_11867_new_n1895
* NET 6206 = abc_11867_new_n1894
* NET 6210 = abc_11867_new_n423
* NET 6213 = abc_11867_new_n1681
* NET 6214 = abc_11867_new_n1799
* NET 6215 = abc_11867_new_n1798
* NET 6220 = abc_11867_new_n609
* NET 6221 = abc_11867_new_n647
* NET 6228 = abc_11867_new_n619
* NET 6230 = abc_11867_new_n577
* NET 6232 = abc_11867_new_n1471
* NET 6233 = abc_11867_new_n434
* NET 6234 = subckt_1689_sff1_x4.sff_s
* NET 6235 = subckt_1689_sff1_x4.sff_m
* NET 6236 = subckt_1689_sff1_x4.u
* NET 6237 = subckt_1689_sff1_x4.ckr
* NET 6238 = subckt_1689_sff1_x4.y
* NET 6239 = subckt_1689_sff1_x4.nckr
* NET 6240 = abc_11867_new_n1404
* NET 6241 = mos6502_nmi_edge
* NET 6243 = abc_11867_new_n617
* NET 6245 = subckt_1672_sff1_x4.sff_s
* NET 6246 = mos6502_op[2]
* NET 6247 = subckt_1672_sff1_x4.y
* NET 6248 = subckt_1672_sff1_x4.sff_m
* NET 6249 = subckt_1672_sff1_x4.u
* NET 6250 = subckt_1672_sff1_x4.ckr
* NET 6251 = abc_11867_new_n587
* NET 6252 = subckt_1672_sff1_x4.nckr
* NET 6255 = abc_11867_new_n1181
* NET 6259 = abc_11867_new_n358
* NET 6260 = subckt_1686_sff1_x4.sff_s
* NET 6261 = mos6502_src_reg[1]
* NET 6262 = subckt_1686_sff1_x4.y
* NET 6263 = subckt_1686_sff1_x4.sff_m
* NET 6264 = subckt_1686_sff1_x4.u
* NET 6265 = subckt_1686_sff1_x4.ckr
* NET 6266 = subckt_1686_sff1_x4.nckr
* NET 6267 = subckt_1682_sff1_x4.sff_s
* NET 6268 = subckt_1682_sff1_x4.sff_m
* NET 6269 = subckt_1682_sff1_x4.u
* NET 6270 = subckt_1682_sff1_x4.ckr
* NET 6271 = subckt_1682_sff1_x4.y
* NET 6272 = subckt_1682_sff1_x4.nckr
* NET 6273 = abc_11867_auto_rtlil_cc_2608_muxgate_11724
* NET 6275 = abc_11867_new_n475_hfns_2
* NET 6276 = abc_11867_new_n482_hfns_1
* NET 6277 = abc_11867_new_n473_hfns_0
* NET 6278 = abc_11867_new_n514_hfns_1
* NET 6280 = abc_11867_new_n626
* NET 6282 = abc_11867_new_n680
* NET 6285 = abc_11867_new_n671
* NET 6286 = abc_11867_new_n533
* NET 6320 = subckt_1758_sff1_x4.y
* NET 6323 = subckt_1758_sff1_x4.sff_m
* NET 6324 = subckt_1758_sff1_x4.ckr
* NET 6331 = subckt_1751_sff1_x4.y
* NET 6332 = subckt_1751_sff1_x4.sff_m
* NET 6333 = subckt_1751_sff1_x4.ckr
* NET 6341 = subckt_1697_sff1_x4.y
* NET 6344 = subckt_1697_sff1_x4.sff_m
* NET 6345 = subckt_1697_sff1_x4.ckr
* NET 6353 = subckt_1674_sff1_x4.y
* NET 6356 = subckt_1674_sff1_x4.sff_m
* NET 6357 = subckt_1674_sff1_x4.ckr
* NET 6358 = abc_11867_new_n387
* NET 6370 = abc_11867_auto_rtlil_cc_2608_muxgate_11862
* NET 6376 = abc_11867_new_n1915
* NET 6379 = abc_11867_new_n1016
* NET 6381 = abc_11867_new_n1019
* NET 6387 = abc_11867_new_n1130
* NET 6394 = abc_11867_new_n1142
* NET 6401 = abc_11867_new_n1145
* NET 6402 = abc_11867_new_n1144
* NET 6403 = subckt_1758_sff1_x4.sff_s
* NET 6404 = abc_11867_auto_rtlil_cc_2608_muxgate_11864
* NET 6406 = subckt_1758_sff1_x4.u
* NET 6407 = subckt_1758_sff1_x4.nckr
* NET 6413 = abc_11867_new_n1122
* NET 6425 = subckt_1751_sff1_x4.sff_s
* NET 6427 = abc_11867_auto_rtlil_cc_2608_muxgate_11850
* NET 6429 = subckt_1751_sff1_x4.u
* NET 6430 = subckt_1751_sff1_x4.nckr
* NET 6431 = abc_11867_new_n1794
* NET 6435 = abc_11867_new_n1772
* NET 6437 = abc_11867_new_n1771
* NET 6440 = abc_11867_new_n981
* NET 6449 = abc_11867_new_n1109
* NET 6451 = abc_11867_new_n422
* NET 6452 = subckt_1697_sff1_x4.sff_s
* NET 6454 = subckt_1697_sff1_x4.u
* NET 6455 = abc_11867_new_n352
* NET 6456 = subckt_1697_sff1_x4.nckr
* NET 6457 = abc_11867_new_n1474
* NET 6465 = di[7]
* NET 6468 = mos6502_dihold[7]
* NET 6469 = subckt_101_nmx2_x1.q
* NET 6473 = abc_11867_new_n1488
* NET 6476 = mos6502_res
* NET 6477 = abc_11867_new_n323
* NET 6478 = abc_11867_auto_rtlil_cc_2608_muxgate_11740
* NET 6483 = abc_11867_new_n1393
* NET 6486 = abc_11867_new_n1401
* NET 6487 = abc_11867_new_n1400
* NET 6489 = abc_11867_new_n363
* NET 6490 = abc_11867_new_n324
* NET 6493 = mos6502_write_back
* NET 6496 = abc_11867_new_n1394
* NET 6497 = abc_11867_new_n1339
* NET 6498 = abc_11867_new_n1338
* NET 6499 = abc_11867_new_n331
* NET 6503 = abc_11867_new_n328
* NET 6506 = abc_11867_new_n1398
* NET 6518 = abc_11867_new_n1365
* NET 6520 = subckt_1674_sff1_x4.sff_s
* NET 6522 = subckt_1674_sff1_x4.u
* NET 6523 = subckt_1674_sff1_x4.nckr
* NET 6524 = abc_11867_new_n1298
* NET 6525 = abc_11867_auto_rtlil_cc_2608_muxgate_11730
* NET 6527 = mos6502_rotate
* NET 6530 = abc_11867_auto_rtlil_cc_2608_muxgate_11706
* NET 6537 = abc_11867_new_n1300
* NET 6538 = abc_11867_auto_rtlil_cc_2608_muxgate_11732
* NET 6543 = abc_11867_auto_rtlil_cc_2608_muxgate_11720
* NET 6545 = mos6502_inc
* NET 6560 = abc_11867_new_n470
* NET 6564 = abc_11867_new_n458
* NET 6569 = abc_11867_new_n457
* NET 6571 = abc_11867_new_n1291
* NET 6574 = abc_11867_new_n532
* NET 6579 = abc_11867_new_n688
* NET 6585 = abc_11867_new_n718
* NET 6586 = abc_11867_new_n761
* NET 6590 = abc_11867_new_n746
* NET 6591 = abc_11867_new_n722
* NET 6592 = abc_11867_new_n744
* NET 6749 = abc_11867_new_n1547
* NET 6751 = subckt_1753_sff1_x4.sff_s
* NET 6752 = subckt_1753_sff1_x4.y
* NET 6755 = subckt_1753_sff1_x4.sff_m
* NET 6756 = subckt_1753_sff1_x4.ckr
* NET 6757 = subckt_1753_sff1_x4.u
* NET 6758 = subckt_1753_sff1_x4.nckr
* NET 6759 = abc_11867_new_n1143
* NET 6760 = abc_11867_new_n341
* NET 6762 = abc_11867_new_n1004
* NET 6764 = abc_11867_new_n1121
* NET 6765 = abc_11867_new_n336
* NET 6766 = abc_11867_new_n335
* NET 6769 = subckt_1752_sff1_x4.sff_s
* NET 6770 = subckt_1752_sff1_x4.y
* NET 6773 = subckt_1752_sff1_x4.sff_m
* NET 6774 = subckt_1752_sff1_x4.u
* NET 6775 = subckt_1752_sff1_x4.ckr
* NET 6776 = subckt_1752_sff1_x4.nckr
* NET 6777 = abc_11867_auto_rtlil_cc_2608_muxgate_11852
* NET 6778 = abc_11867_new_n1896
* NET 6784 = abc_11867_new_n1112
* NET 6788 = abc_11867_new_n1117
* NET 6789 = abc_11867_new_n1116
* NET 6791 = abc_11867_new_n944
* NET 6793 = do[7]
* NET 6796 = abc_11867_new_n890
* NET 6798 = abc_11867_new_n976
* NET 6803 = abc_11867_new_n333
* NET 6806 = abc_11867_new_n929
* NET 6809 = abc_11867_new_n887
* NET 6811 = abc_11867_new_n1844
* NET 6815 = abc_11867_new_n619_hfns_2
* NET 6817 = abc_11867_new_n888
* NET 6819 = mos6502_i
* NET 6820 = abc_11867_new_n903
* NET 6822 = subckt_1713_sff1_x4.sff_s
* NET 6824 = subckt_1713_sff1_x4.y
* NET 6826 = subckt_1713_sff1_x4.sff_m
* NET 6827 = abc_11867_auto_rtlil_cc_2608_muxgate_11776
* NET 6829 = subckt_1713_sff1_x4.u
* NET 6830 = subckt_1713_sff1_x4.nckr
* NET 6831 = subckt_1713_sff1_x4.ckr
* NET 6833 = subckt_1670_sff1_x4.sff_s
* NET 6835 = subckt_1670_sff1_x4.y
* NET 6837 = subckt_1670_sff1_x4.sff_m
* NET 6838 = subckt_1670_sff1_x4.u
* NET 6839 = subckt_1670_sff1_x4.ckr
* NET 6840 = subckt_1670_sff1_x4.nckr
* NET 6842 = subckt_1699_sff1_x4.sff_s
* NET 6843 = subckt_1699_sff1_x4.y
* NET 6845 = subckt_1699_sff1_x4.sff_m
* NET 6847 = abc_11867_auto_rtlil_cc_2608_muxgate_11746
* NET 6848 = subckt_1699_sff1_x4.u
* NET 6849 = subckt_1699_sff1_x4.ckr
* NET 6850 = subckt_1699_sff1_x4.nckr
* NET 6851 = abc_11867_new_n1367
* NET 6859 = abc_11867_new_n1181_hfns_2
* NET 6861 = abc_11867_new_n764
* NET 6862 = abc_11867_new_n1363
* NET 6863 = abc_11867_new_n344
* NET 6864 = abc_11867_new_n384
* NET 6866 = abc_11867_new_n1297
* NET 6867 = mos6502_php
* NET 6869 = subckt_1661_sff1_x4.sff_s
* NET 6870 = subckt_1661_sff1_x4.y
* NET 6872 = subckt_1661_sff1_x4.sff_m
* NET 6874 = subckt_1661_sff1_x4.u
* NET 6875 = subckt_1661_sff1_x4.ckr
* NET 6876 = subckt_1661_sff1_x4.nckr
* NET 6877 = abc_11867_new_n1221
* NET 6879 = mos6502_dst_reg[1]
* NET 6881 = subckt_1688_sff1_x4.sff_s
* NET 6882 = subckt_1688_sff1_x4.y
* NET 6884 = subckt_1688_sff1_x4.sff_m
* NET 6886 = subckt_1688_sff1_x4.ckr
* NET 6887 = subckt_1688_sff1_x4.u
* NET 6888 = subckt_1688_sff1_x4.nckr
* NET 6889 = abc_11867_new_n388
* NET 6890 = abc_11867_new_n1317
* NET 6891 = abc_11867_auto_rtlil_cc_2608_muxgate_11736
* NET 6894 = abc_11867_new_n1315
* NET 6895 = abc_11867_new_n685
* NET 6896 = abc_11867_new_n697
* NET 6898 = abc_11867_new_n760
* NET 6900 = abc_11867_new_n748
* NET 6901 = abc_11867_new_n681
* NET 6902 = abc_11867_new_n677
* NET 6904 = abc_11867_new_n759
* NET 6905 = abc_11867_new_n756
* NET 6906 = abc_11867_new_n687
* NET 6908 = abc_11867_new_n628
* NET 6941 = abc_11867_new_n1559
* NET 6942 = abc_11867_new_n1546
* NET 6959 = abc_11867_new_n1001
* NET 6963 = abc_11867_auto_rtlil_cc_2608_muxgate_11854
* NET 6967 = abc_11867_new_n1892
* NET 6978 = abc_11867_new_n1675
* NET 6992 = mos6502_alu_hc
* NET 6993 = abc_11867_new_n1120
* NET 6994 = abc_11867_new_n1114
* NET 6997 = abc_11867_new_n1115
* NET 6998 = abc_11867_new_n1113
* NET 7004 = abc_11867_new_n1108
* NET 7006 = abc_11867_new_n1107
* NET 7007 = abc_11867_new_n1106
* NET 7012 = abc_11867_new_n1674
* NET 7019 = abc_11867_new_n372
* NET 7022 = abc_11867_new_n980
* NET 7023 = abc_11867_new_n977
* NET 7027 = abc_11867_new_n989
* NET 7031 = abc_11867_new_n985
* NET 7033 = abc_11867_new_n988
* NET 7036 = abc_11867_new_n1481
* NET 7037 = mos6502_abl[0]
* NET 7041 = abc_11867_new_n648
* NET 7042 = abc_11867_new_n611
* NET 7045 = abc_11867_new_n1011
* NET 7046 = abc_11867_new_n1010
* NET 7050 = abc_11867_new_n1008
* NET 7058 = abc_11867_new_n1496
* NET 7059 = abc_11867_new_n1498
* NET 7061 = abc_11867_new_n1499
* NET 7063 = abc_11867_new_n1673
* NET 7068 = abc_11867_new_n595
* NET 7069 = abc_11867_new_n631
* NET 7082 = abc_11867_new_n1099
* NET 7084 = abc_11867_new_n329
* NET 7085 = mos6502_op[0]
* NET 7089 = abc_11867_auto_rtlil_cc_2608_muxgate_11698
* NET 7096 = subckt_1673_sff1_x4.sff_s
* NET 7098 = rdy_hfns_4
* NET 7099 = subckt_1673_sff1_x4.y
* NET 7101 = subckt_1673_sff1_x4.sff_m
* NET 7104 = subckt_1673_sff1_x4.u
* NET 7105 = subckt_1673_sff1_x4.nckr
* NET 7106 = subckt_1673_sff1_x4.ckr
* NET 7108 = abc_11867_auto_rtlil_cc_2608_muxgate_11704
* NET 7109 = mos6502_op[3]
* NET 7117 = mos6502_cli
* NET 7119 = subckt_1666_sff1_x4.sff_s
* NET 7122 = subckt_1666_sff1_x4.y
* NET 7124 = subckt_1666_sff1_x4.sff_m
* NET 7126 = subckt_1666_sff1_x4.ckr
* NET 7127 = subckt_1666_sff1_x4.u
* NET 7128 = subckt_1666_sff1_x4.nckr
* NET 7129 = abc_11867_new_n1237
* NET 7131 = abc_11867_auto_rtlil_cc_2608_muxgate_11702
* NET 7132 = subckt_1667_sff1_x4.sff_s
* NET 7136 = subckt_1667_sff1_x4.y
* NET 7139 = subckt_1667_sff1_x4.sff_m
* NET 7140 = subckt_1667_sff1_x4.ckr
* NET 7141 = subckt_1667_sff1_x4.u
* NET 7142 = abc_11867_new_n1185
* NET 7143 = subckt_1667_sff1_x4.nckr
* NET 7144 = abc_11867_auto_rtlil_cc_2608_muxgate_11680
* NET 7147 = mos6502_load_only
* NET 7149 = subckt_1681_sff1_x4.sff_s
* NET 7153 = subckt_1681_sff1_x4.y
* NET 7154 = abc_11867_auto_rtlil_cc_2608_muxgate_11722
* NET 7156 = subckt_1681_sff1_x4.sff_m
* NET 7157 = subckt_1681_sff1_x4.ckr
* NET 7158 = subckt_1681_sff1_x4.u
* NET 7160 = subckt_1681_sff1_x4.nckr
* NET 7161 = abc_11867_new_n757
* NET 7165 = abc_11867_new_n1278
* NET 7167 = abc_11867_new_n1314
* NET 7176 = abc_11867_new_n629
* NET 7177 = abc_11867_new_n1313
* NET 7190 = abc_11867_new_n750
* NET 7201 = abc_11867_new_n459
* NET 7204 = abc_11867_new_n547
* NET 7212 = abc_11867_new_n698
* NET 7217 = abc_11867_new_n758
* NET 7403 = abc_11867_new_n1025
* NET 7404 = abc_11867_new_n419
* NET 7408 = abc_11867_new_n1137
* NET 7410 = abc_11867_new_n1018
* NET 7411 = abc_11867_new_n373
* NET 7414 = abc_11867_new_n1135
* NET 7415 = abc_11867_new_n1128
* NET 7418 = mos6502_abl[6]
* NET 7419 = abc_11867_new_n1531
* NET 7421 = abc_11867_new_n1129
* NET 7422 = abc_11867_new_n1131
* NET 7425 = mos6502_abl[5]
* NET 7426 = abc_11867_new_n1727
* NET 7430 = abc_11867_new_n904
* NET 7432 = abc_11867_new_n1749
* NET 7437 = abc_11867_new_n1671
* NET 7439 = abc_11867_new_n984
* NET 7444 = abc_11867_new_n349
* NET 7445 = abc_11867_new_n1491
* NET 7447 = abc_11867_new_n1500
* NET 7448 = abc_11867_new_n350
* NET 7450 = mos6502_abl[4]
* NET 7451 = abc_11867_new_n979
* NET 7452 = abc_11867_new_n368
* NET 7455 = abc_11867_new_n1480
* NET 7457 = abc_11867_new_n1461
* NET 7459 = abc_11867_new_n1482
* NET 7460 = abc_11867_new_n348
* NET 7463 = abc_11867_new_n1478
* NET 7465 = abc_11867_new_n585
* NET 7466 = mos6502_abl[2]
* NET 7467 = abc_11867_new_n1490
* NET 7468 = abc_11867_new_n1489
* NET 7471 = abc_11867_new_n987
* NET 7474 = mos6502_abl[1]
* NET 7475 = abc_11867_new_n369
* NET 7476 = abc_11867_new_n1098
* NET 7478 = abc_11867_new_n431_hfns_1
* NET 7480 = abc_11867_new_n1403
* NET 7484 = mos6502_alu_co
* NET 7490 = subckt_1671_sff1_x4.sff_s
* NET 7492 = subckt_1671_sff1_x4.y
* NET 7494 = subckt_1671_sff1_x4.sff_m
* NET 7495 = subckt_1671_sff1_x4.u
* NET 7496 = subckt_1671_sff1_x4.ckr
* NET 7497 = subckt_1671_sff1_x4.nckr
* NET 7498 = abc_11867_new_n1397
* NET 7501 = subckt_1676_sff1_x4.sff_s
* NET 7503 = subckt_1676_sff1_x4.y
* NET 7505 = subckt_1676_sff1_x4.sff_m
* NET 7506 = subckt_1676_sff1_x4.u
* NET 7507 = subckt_1676_sff1_x4.nckr
* NET 7508 = subckt_1676_sff1_x4.ckr
* NET 7509 = abc_11867_auto_rtlil_cc_2608_muxgate_11710
* NET 7514 = abc_11867_new_n430_hfns_0
* NET 7516 = mos6502_sei
* NET 7517 = abc_11867_new_n1204
* NET 7518 = abc_11867_auto_rtlil_cc_2608_muxgate_11690
* NET 7520 = abc_11867_new_n1207
* NET 7521 = abc_11867_auto_rtlil_cc_2608_muxgate_11692
* NET 7523 = abc_11867_new_n557
* NET 7525 = abc_11867_new_n1205
* NET 7526 = abc_11867_new_n1257
* NET 7527 = abc_11867_new_n559
* NET 7529 = abc_11867_new_n1256
* NET 7531 = abc_11867_new_n1305
* NET 7532 = abc_11867_new_n1306
* NET 7533 = abc_11867_new_n1277
* NET 7534 = abc_11867_new_n1239
* NET 7535 = abc_11867_new_n1320
* NET 7536 = abc_11867_new_n749
* NET 7538 = abc_11867_new_n1319
* NET 7539 = abc_11867_new_n1318
* NET 7540 = abc_11867_new_n747
* NET 7583 = abc_11867_new_n418
* NET 7585 = abc_11867_new_n1532
* NET 7594 = abc_11867_new_n1358
* NET 7600 = abc_11867_new_n1540
* NET 7601 = mos6502_abl[7]
* NET 7605 = abc_11867_new_n1003
* NET 7606 = abc_11867_new_n371
* NET 7611 = mos6502_abl[3]
* NET 7615 = abc_11867_new_n619_hfns_1
* NET 7618 = abc_11867_new_n1506
* NET 7622 = subckt_1733_sff1_x4.sff_s
* NET 7623 = subckt_1733_sff1_x4.y
* NET 7627 = subckt_1733_sff1_x4.sff_m
* NET 7628 = subckt_1733_sff1_x4.ckr
* NET 7629 = subckt_1733_sff1_x4.u
* NET 7630 = subckt_1733_sff1_x4.nckr
* NET 7631 = abc_11867_new_n1487
* NET 7633 = abc_11867_new_n1493
* NET 7634 = abc_11867_auto_rtlil_cc_2608_muxgate_11814
* NET 7638 = subckt_1732_sff1_x4.sff_s
* NET 7639 = subckt_1732_sff1_x4.y
* NET 7643 = subckt_1732_sff1_x4.sff_m
* NET 7644 = subckt_1732_sff1_x4.ckr
* NET 7645 = subckt_1732_sff1_x4.u
* NET 7646 = subckt_1732_sff1_x4.nckr
* NET 7648 = abc_11867_new_n947
* NET 7652 = mos6502_pc[0]
* NET 7655 = mos6502_adj_bcd
* NET 7657 = subckt_1714_sff1_x4.sff_s
* NET 7661 = subckt_1714_sff1_x4.y
* NET 7662 = subckt_1714_sff1_x4.sff_m
* NET 7664 = subckt_1714_sff1_x4.ckr
* NET 7665 = subckt_1714_sff1_x4.u
* NET 7666 = subckt_1714_sff1_x4.nckr
* NET 7667 = abc_11867_new_n1484
* NET 7670 = abc_11867_new_n1464
* NET 7672 = abc_11867_new_n1470
* NET 7673 = abc_11867_new_n1469
* NET 7678 = abc_11867_new_n471_hfns_2
* NET 7684 = abc_11867_new_n1476
* NET 7685 = abc_11867_new_n1463
* NET 7689 = abc_11867_new_n370
* NET 7690 = abc_11867_new_n973
* NET 7695 = abc_11867_new_n1351
* NET 7701 = abc_11867_new_n879
* NET 7702 = abc_11867_new_n1375
* NET 7704 = abc_11867_new_n1378
* NET 7711 = abc_11867_new_n473_hfns_1
* NET 7719 = abc_11867_new_n376
* NET 7721 = abc_11867_new_n431_hfns_0
* NET 7727 = abc_11867_new_n1402
* NET 7739 = mos6502_compare
* NET 7740 = abc_11867_new_n1395
* NET 7747 = abc_11867_new_n1364
* NET 7748 = subckt_1041_nmx2_x1.q
* NET 7749 = mos6502_op[1]
* NET 7752 = abc_11867_auto_rtlil_cc_2608_muxgate_11700
* NET 7766 = abc_11867_new_n435
* NET 7770 = abc_11867_new_n1396
* NET 7773 = subckt_1662_sff1_x4.sff_s
* NET 7774 = subckt_1662_sff1_x4.y
* NET 7777 = subckt_1662_sff1_x4.sff_m
* NET 7779 = subckt_1662_sff1_x4.u
* NET 7780 = subckt_1662_sff1_x4.ckr
* NET 7781 = subckt_1662_sff1_x4.nckr
* NET 7784 = abc_11867_new_n1230
* NET 7786 = abc_11867_new_n1251
* NET 7798 = abc_11867_new_n1296
* NET 7802 = abc_11867_auto_rtlil_cc_2608_muxgate_11682
* NET 7805 = abc_11867_new_n1254
* NET 7813 = abc_11867_new_n1190
* NET 7817 = abc_11867_new_n1261
* NET 7824 = abc_11867_new_n558
* NET 7825 = abc_11867_new_n468
* NET 7828 = abc_11867_new_n1276
* NET 7835 = abc_11867_new_n1244
* NET 7837 = abc_11867_new_n469
* NET 7840 = abc_11867_new_n745
* NET 7848 = abc_11867_new_n721
* NET 7852 = abc_11867_new_n439
* NET 8000 = abc_11867_new_n1017
* NET 8007 = abc_11867_new_n1524
* NET 8009 = abc_11867_new_n1523
* NET 8012 = abc_11867_new_n912
* NET 8014 = abc_11867_new_n898
* NET 8015 = spare_buffer_11.q
* NET 8016 = spare_buffer_10.q
* NET 8017 = do[6]
* NET 8019 = abc_11867_auto_rtlil_cc_2608_muxgate_11812
* NET 8021 = abc_11867_new_n996
* NET 8022 = abc_11867_new_n945
* NET 8026 = abc_11867_new_n1377
* NET 8030 = abc_11867_flatten_mos6502_0_adj_bcd_0_0
* NET 8038 = abc_11867_new_n1354
* NET 8042 = abc_11867_new_n1235
* NET 8046 = abc_11867_new_n1187
* NET 8047 = reset_root_bl_0
* NET 8048 = clk_root_bl_2
* NET 8049 = abc_11867_new_n1229
* NET 8050 = abc_11867_new_n1208
* NET 8051 = abc_11867_new_n804
* NET 8052 = abc_11867_new_n465
* NET 8053 = abc_11867_new_n1250
* NET 8054 = abc_11867_new_n1245
* NET 8056 = abc_11867_new_n1311
* NET 8059 = abc_11867_new_n695
* NET 8060 = abc_11867_new_n461
* NET 8062 = abc_11867_new_n443
* NET 8063 = abc_11867_new_n446
* NET 8064 = di[6]
* NET 8065 = subckt_97_nmx2_x1.q
* NET 8070 = abc_11867_new_n1541
* NET 8071 = subckt_1696_sff1_x4.sff_s
* NET 8072 = mos6502_dihold[6]
* NET 8073 = subckt_1696_sff1_x4.y
* NET 8074 = subckt_1696_sff1_x4.sff_m
* NET 8075 = subckt_1696_sff1_x4.u
* NET 8076 = subckt_1696_sff1_x4.ckr
* NET 8077 = subckt_1696_sff1_x4.nckr
* NET 8080 = abc_11867_new_n1522
* NET 8081 = abc_11867_new_n1507
* NET 8082 = mos6502_pc[1]
* NET 8084 = abc_11867_new_n910
* NET 8086 = abc_11867_new_n897
* NET 8089 = abc_11867_new_n937
* NET 8090 = mos6502_pc[8]
* NET 8091 = abc_11867_new_n586
* NET 8092 = abc_11867_new_n481
* NET 8093 = abc_11867_new_n1460
* NET 8094 = abc_11867_new_n1485
* NET 8095 = abc_11867_new_n1483
* NET 8096 = abc_11867_new_n995
* NET 8097 = abc_11867_new_n993
* NET 8100 = abc_11867_new_n432
* NET 8101 = abc_11867_new_n896
* NET 8103 = abc_11867_new_n1359
* NET 8106 = abc_11867_new_n1376
* NET 8107 = abc_11867_new_n1379
* NET 8112 = abc_11867_new_n1355
* NET 8113 = abc_11867_new_n1350
* NET 8114 = subckt_1677_sff1_x4.sff_s
* NET 8115 = subckt_1677_sff1_x4.sff_m
* NET 8116 = subckt_1677_sff1_x4.u
* NET 8117 = subckt_1677_sff1_x4.ckr
* NET 8118 = subckt_1677_sff1_x4.y
* NET 8119 = subckt_1677_sff1_x4.nckr
* NET 8120 = abc_11867_auto_rtlil_cc_2608_muxgate_11714
* NET 8121 = abc_11867_new_n1264
* NET 8122 = mos6502_adc_bcd
* NET 8123 = abc_11867_new_n1265
* NET 8124 = mos6502_state[3]
* NET 8126 = abc_11867_new_n430_hfns_1
* NET 8128 = abc_11867_new_n1274
* NET 8130 = subckt_1669_sff1_x4.sff_s
* NET 8131 = subckt_1669_sff1_x4.y
* NET 8132 = subckt_1669_sff1_x4.sff_m
* NET 8133 = subckt_1669_sff1_x4.u
* NET 8134 = subckt_1669_sff1_x4.ckr
* NET 8135 = subckt_1669_sff1_x4.nckr
* NET 8136 = subckt_1678_sff1_x4.sff_s
* NET 8138 = subckt_1678_sff1_x4.y
* NET 8139 = subckt_1678_sff1_x4.sff_m
* NET 8141 = subckt_1678_sff1_x4.u
* NET 8142 = subckt_1678_sff1_x4.ckr
* NET 8144 = subckt_1678_sff1_x4.nckr
* NET 8145 = reset_root_0
* NET 8151 = abc_11867_new_n1246
* NET 8152 = abc_11867_new_n460
* NET 8155 = abc_11867_new_n1255
* NET 8192 = subckt_1737_sff1_x4.y
* NET 8196 = subckt_1737_sff1_x4.sff_m
* NET 8197 = subckt_1737_sff1_x4.ckr
* NET 8206 = abc_11867_new_n1360
* NET 8212 = abc_11867_new_n1352
* NET 8220 = subckt_1679_sff1_x4.y
* NET 8221 = subckt_1679_sff1_x4.sff_m
* NET 8222 = subckt_1679_sff1_x4.ckr
* NET 8225 = subckt_1668_sff1_x4.y
* NET 8228 = subckt_1668_sff1_x4.sff_m
* NET 8229 = subckt_1668_sff1_x4.ckr
* NET 8244 = abc_11867_new_n755
* NET 8245 = subckt_1737_sff1_x4.sff_s
* NET 8247 = subckt_1737_sff1_x4.u
* NET 8248 = subckt_1737_sff1_x4.nckr
* NET 8252 = abc_11867_auto_rtlil_cc_2608_muxgate_11822
* NET 8261 = abc_11867_new_n1528
* NET 8262 = abc_11867_new_n1525
* NET 8267 = abc_11867_new_n1508
* NET 8277 = abc_11867_new_n946
* NET 8286 = spare_buffer_9.q
* NET 8290 = abc_11867_new_n1387
* NET 8291 = abc_11867_new_n1388
* NET 8297 = mos6502_alu_out[0]
* NET 8305 = mos6502_abh[0]
* NET 8309 = abc_11867_new_n1536
* NET 8310 = abc_11867_new_n1530
* NET 8312 = abc_11867_auto_rtlil_cc_2608_muxgate_11824
* NET 8313 = abc_11867_new_n1537
* NET 8316 = abc_11867_new_n618
* NET 8318 = abc_11867_new_n886
* NET 8327 = abc_11867_new_n1380
* NET 8328 = abc_11867_new_n1381
* NET 8340 = abc_11867_new_n1356
* NET 8341 = abc_11867_new_n1361
* NET 8358 = abc_11867_new_n1353
* NET 8385 = subckt_1679_sff1_x4.sff_s
* NET 8388 = mos6502_adc_sbc
* NET 8390 = abc_11867_auto_rtlil_cc_2608_muxgate_11718
* NET 8392 = subckt_1679_sff1_x4.u
* NET 8393 = subckt_1679_sff1_x4.nckr
* NET 8394 = abc_11867_new_n1268
* NET 8395 = abc_11867_new_n1267
* NET 8402 = abc_11867_new_n1266
* NET 8403 = abc_11867_new_n1263
* NET 8407 = mos6502_clc
* NET 8408 = abc_11867_new_n325
* NET 8409 = mos6502_shift
* NET 8410 = subckt_1668_sff1_x4.sff_s
* NET 8411 = mos6502_clv
* NET 8419 = subckt_1668_sff1_x4.u
* NET 8420 = subckt_1668_sff1_x4.nckr
* NET 8424 = clk_root_0
* NET 8426 = abc_11867_new_n1220
* NET 8429 = abc_11867_new_n1227
* NET 8430 = abc_11867_new_n1222
* NET 8431 = abc_11867_new_n1226
* NET 8437 = abc_11867_new_n1223
* NET 8443 = abc_11867_new_n1218
* NET 8453 = abc_11867_new_n540
* NET 8458 = abc_11867_new_n1243
* NET 8459 = abc_11867_new_n1312
* NET 8460 = abc_11867_new_n1308
* NET 8472 = abc_11867_new_n754
* NET 8475 = abc_11867_new_n696
* NET 8477 = abc_11867_new_n753
* NET 8610 = abc_11867_new_n1543
* NET 8612 = abc_11867_new_n1545
* NET 8613 = abc_11867_new_n1527
* NET 8615 = abc_11867_new_n1534
* NET 8616 = abc_11867_new_n1533
* NET 8617 = mos6502_pc[6]
* NET 8620 = abc_11867_new_n415
* NET 8621 = abc_11867_new_n414
* NET 8623 = mos6502_pc[5]
* NET 8624 = abc_11867_new_n1521
* NET 8627 = abc_11867_new_n1505
* NET 8629 = abc_11867_new_n1511
* NET 8633 = abc_11867_new_n889
* NET 8635 = abc_11867_new_n842
* NET 8636 = abc_11867_new_n844
* NET 8638 = abc_11867_new_n911
* NET 8642 = mos6502_alu_out[7]
* NET 8643 = abc_11867_new_n428_hfns_2
* NET 8644 = abc_11867_new_n1473
* NET 8645 = abc_11867_new_n1516
* NET 8647 = abc_11867_new_n1515
* NET 8648 = abc_11867_new_n1514
* NET 8650 = abc_11867_new_n938
* NET 8651 = abc_11867_new_n940
* NET 8652 = abc_11867_new_n939
* NET 8654 = abc_11867_new_n359
* NET 8657 = abc_11867_new_n1552
* NET 8658 = abc_11867_new_n1551
* NET 8659 = abc_11867_new_n1553
* NET 8661 = abc_11867_new_n490_hfns_1
* NET 8662 = abc_11867_new_n432_hfns_2
* NET 8664 = subckt_1711_sff1_x4.sff_s
* NET 8667 = subckt_1711_sff1_x4.y
* NET 8668 = subckt_1711_sff1_x4.sff_m
* NET 8670 = abc_11867_auto_rtlil_cc_2608_muxgate_11772
* NET 8671 = subckt_1711_sff1_x4.u
* NET 8672 = subckt_1711_sff1_x4.ckr
* NET 8673 = subckt_1711_sff1_x4.nckr
* NET 8675 = abc_11867_new_n1383
* NET 8679 = abc_11867_new_n1390
* NET 8682 = abc_11867_new_n1389
* NET 8684 = abc_11867_new_n1385
* NET 8685 = abc_11867_new_n1384
* NET 8690 = abc_11867_new_n1386
* NET 8691 = mos6502_c
* NET 8694 = mos6502_n
* NET 8697 = abc_11867_new_n1372
* NET 8699 = mos6502_alu_out[3]
* NET 8703 = abc_11867_new_n1373
* NET 8708 = abc_11867_new_n326
* NET 8709 = abc_11867_new_n582
* NET 8712 = abc_11867_new_n1371
* NET 8713 = abc_11867_new_n433
* NET 8714 = subckt_1048_nmx2_x1.q
* NET 8716 = subckt_1657_sff1_x4.sff_s
* NET 8717 = subckt_1657_sff1_x4.y
* NET 8720 = subckt_1657_sff1_x4.sff_m
* NET 8721 = subckt_1657_sff1_x4.u
* NET 8722 = subckt_1657_sff1_x4.ckr
* NET 8723 = subckt_1657_sff1_x4.nckr
* NET 8724 = abc_11867_auto_rtlil_cc_2608_muxgate_11696
* NET 8725 = mos6502_bit_ins
* NET 8728 = abc_11867_new_n1217
* NET 8731 = abc_11867_new_n327
* NET 8733 = abc_11867_new_n1181_hfns_1
* NET 8734 = abc_11867_auto_rtlil_cc_2608_muxgate_11716
* NET 8735 = subckt_950_nmx2_x1.q
* NET 8738 = subckt_1663_sff1_x4.sff_s
* NET 8740 = subckt_1663_sff1_x4.sff_m
* NET 8741 = subckt_1663_sff1_x4.y
* NET 8743 = subckt_1663_sff1_x4.u
* NET 8744 = subckt_1663_sff1_x4.nckr
* NET 8745 = subckt_1663_sff1_x4.ckr
* NET 8746 = abc_11867_new_n546
* NET 8748 = mos6502_sec
* NET 8749 = abc_11867_new_n1192
* NET 8750 = abc_11867_new_n1195
* NET 8751 = abc_11867_auto_rtlil_cc_2608_muxgate_11684
* NET 8753 = abc_11867_new_n1228
* NET 8754 = abc_11867_new_n1260
* NET 8756 = abc_11867_new_n1238
* NET 8758 = abc_11867_new_n1249
* NET 8760 = abc_11867_new_n1248
* NET 8762 = abc_11867_new_n1295
* NET 8765 = abc_11867_new_n1304
* NET 8767 = abc_11867_new_n1290
* NET 8768 = abc_11867_new_n1303
* NET 8770 = abc_11867_new_n535
* NET 8816 = do[5]
* NET 8817 = abc_11867_new_n1526
* NET 8821 = abc_11867_new_n1608
* NET 8824 = abc_11867_new_n1535
* NET 8831 = abc_11867_new_n1556
* NET 8833 = abc_11867_new_n1544
* NET 8834 = abc_11867_new_n1479
* NET 8835 = abc_11867_new_n1542
* NET 8839 = mos6502_pc[7]
* NET 8840 = di[5]
* NET 8846 = subckt_93_nmx2_x1.q
* NET 8848 = mos6502_pc[3]
* NET 8850 = subckt_1735_sff1_x4.sff_s
* NET 8852 = subckt_1735_sff1_x4.y
* NET 8855 = subckt_1735_sff1_x4.sff_m
* NET 8856 = abc_11867_auto_rtlil_cc_2608_muxgate_11818
* NET 8858 = subckt_1735_sff1_x4.u
* NET 8859 = subckt_1735_sff1_x4.ckr
* NET 8860 = subckt_1735_sff1_x4.nckr
* NET 8862 = abc_11867_new_n1517
* NET 8864 = abc_11867_new_n1503
* NET 8865 = abc_11867_new_n1502
* NET 8866 = abc_11867_new_n1495
* NET 8869 = mos6502_pc[2]
* NET 8870 = subckt_1734_sff1_x4.sff_s
* NET 8873 = subckt_1734_sff1_x4.y
* NET 8876 = subckt_1734_sff1_x4.sff_m
* NET 8878 = abc_11867_auto_rtlil_cc_2608_muxgate_11816
* NET 8879 = subckt_1734_sff1_x4.ckr
* NET 8880 = subckt_1734_sff1_x4.u
* NET 8881 = subckt_1734_sff1_x4.nckr
* NET 8882 = abc_11867_new_n1726
* NET 8885 = mos6502_alu_out[6]
* NET 8893 = abc_11867_new_n343
* NET 8903 = abc_11867_new_n1009
* NET 8906 = abc_11867_new_n411
* NET 8912 = abc_11867_new_n1555
* NET 8913 = abc_11867_new_n1554
* NET 8915 = abc_11867_new_n1550
* NET 8918 = mos6502_alu_out[4]
* NET 8921 = abc_11867_new_n428_hfns_4
* NET 8922 = abc_11867_new_n485_hfns_0
* NET 8930 = mos6502_alu_out[1]
* NET 8937 = abc_11867_new_n1864
* NET 8938 = abc_11867_new_n1040
* NET 8942 = subckt_1712_sff1_x4.y
* NET 8943 = subckt_1712_sff1_x4.sff_s
* NET 8948 = subckt_1712_sff1_x4.sff_m
* NET 8949 = abc_11867_auto_rtlil_cc_2608_muxgate_11774
* NET 8950 = subckt_1712_sff1_x4.ckr
* NET 8951 = subckt_1712_sff1_x4.u
* NET 8952 = subckt_1712_sff1_x4.nckr
* NET 8954 = mos6502_z
* NET 8970 = mos6502_d
* NET 8971 = subckt_1710_sff1_x4.sff_s
* NET 8973 = subckt_1710_sff1_x4.y
* NET 8977 = abc_11867_auto_rtlil_cc_2608_muxgate_11770
* NET 8979 = subckt_1710_sff1_x4.sff_m
* NET 8980 = subckt_1710_sff1_x4.u
* NET 8981 = subckt_1710_sff1_x4.ckr
* NET 8982 = subckt_1710_sff1_x4.nckr
* NET 8983 = abc_11867_new_n332
* NET 8985 = abc_11867_new_n705
* NET 8989 = abc_11867_new_n706
* NET 8995 = abc_11867_new_n345
* NET 8999 = abc_11867_new_n707
* NET 9002 = abc_11867_new_n708
* NET 9006 = abc_11867_auto_rtlil_cc_2608_muxgate_11672
* NET 9007 = mos6502_cond_code[0]
* NET 9016 = abc_11867_new_n1370
* NET 9020 = abc_11867_new_n478_hfns_1
* NET 9028 = abc_11867_new_n1210
* NET 9029 = abc_11867_new_n1214
* NET 9030 = abc_11867_auto_rtlil_cc_2608_muxgate_11694
* NET 9033 = mos6502_plp
* NET 9035 = subckt_1660_sff1_x4.sff_s
* NET 9039 = subckt_1660_sff1_x4.y
* NET 9041 = subckt_1660_sff1_x4.sff_m
* NET 9042 = subckt_1660_sff1_x4.ckr
* NET 9043 = subckt_1660_sff1_x4.u
* NET 9044 = abc_11867_new_n1182
* NET 9045 = subckt_1660_sff1_x4.nckr
* NET 9046 = abc_11867_new_n1183
* NET 9047 = abc_11867_auto_rtlil_cc_2608_muxgate_11678
* NET 9051 = abc_11867_new_n538
* NET 9057 = abc_11867_new_n674
* NET 9061 = abc_11867_new_n676
* NET 9066 = abc_11867_new_n1232
* NET 9073 = abc_11867_new_n545
* NET 9074 = abc_11867_new_n1282
* NET 9080 = abc_11867_new_n675
* NET 9081 = abc_11867_new_n1294
* NET 9083 = abc_11867_new_n1188
* NET 9087 = abc_11867_new_n1247
* NET 9095 = abc_11867_new_n464
* NET 9100 = abc_11867_new_n751
* NET 9103 = abc_11867_new_n1310
* NET 9104 = abc_11867_new_n1309
* NET 9107 = abc_11867_new_n534_hfns_1
* NET 9266 = subckt_1743_sff1_x4.sff_s
* NET 9267 = subckt_1743_sff1_x4.y
* NET 9270 = subckt_1743_sff1_x4.sff_m
* NET 9271 = subckt_1743_sff1_x4.u
* NET 9272 = subckt_1743_sff1_x4.ckr
* NET 9273 = subckt_1743_sff1_x4.nckr
* NET 9275 = abc_11867_new_n1002
* NET 9280 = subckt_1736_sff1_x4.sff_s
* NET 9281 = subckt_1736_sff1_x4.y
* NET 9284 = subckt_1736_sff1_x4.sff_m
* NET 9285 = subckt_1736_sff1_x4.u
* NET 9286 = subckt_1736_sff1_x4.ckr
* NET 9287 = mos6502_pc[4]
* NET 9288 = subckt_1736_sff1_x4.nckr
* NET 9290 = abc_11867_new_n1518
* NET 9291 = abc_11867_new_n1513
* NET 9292 = abc_11867_auto_rtlil_cc_2608_muxgate_11820
* NET 9293 = abc_11867_new_n1519
* NET 9295 = abc_11867_new_n1510
* NET 9296 = abc_11867_new_n1501
* NET 9297 = abc_11867_new_n1492
* NET 9298 = abc_11867_new_n1509
* NET 9300 = abc_11867_new_n1748
* NET 9304 = mos6502_alu_out[5]
* NET 9305 = abc_11867_new_n342
* NET 9306 = abc_11867_new_n1085
* NET 9308 = abc_11867_new_n428_hfns_3
* NET 9309 = abc_11867_new_n485_hfns_1
* NET 9310 = abc_11867_new_n1793
* NET 9313 = mos6502_alu_out[2]
* NET 9314 = abc_11867_new_n490_hfns_0
* NET 9315 = abc_11867_new_n410
* NET 9316 = di[4]
* NET 9320 = subckt_89_nmx2_x1.q
* NET 9321 = abc_11867_new_n1770
* NET 9323 = abc_11867_new_n1818
* NET 9329 = abc_11867_new_n1070
* NET 9332 = abc_11867_new_n1073
* NET 9333 = abc_11867_new_n339
* NET 9335 = mos6502_v
* NET 9336 = subckt_1708_sff1_x4.sff_s
* NET 9338 = subckt_1708_sff1_x4.y
* NET 9339 = subckt_1708_sff1_x4.sff_m
* NET 9341 = abc_11867_auto_rtlil_cc_2608_muxgate_11764
* NET 9343 = subckt_1708_sff1_x4.u
* NET 9344 = subckt_1708_sff1_x4.nckr
* NET 9345 = subckt_1708_sff1_x4.ckr
* NET 9346 = abc_11867_new_n1843
* NET 9347 = abc_11867_new_n1672
* NET 9350 = mos6502_cond_code[2]
* NET 9352 = subckt_1659_sff1_x4.sff_s
* NET 9354 = subckt_1659_sff1_x4.y
* NET 9355 = abc_11867_auto_rtlil_cc_2608_muxgate_11676
* NET 9357 = subckt_1659_sff1_x4.sff_m
* NET 9358 = subckt_1659_sff1_x4.u
* NET 9359 = subckt_1659_sff1_x4.nckr
* NET 9360 = subckt_1659_sff1_x4.ckr
* NET 9362 = abc_11867_new_n424
* NET 9367 = subckt_1658_sff1_x4.sff_s
* NET 9368 = subckt_1658_sff1_x4.y
* NET 9370 = subckt_1658_sff1_x4.sff_m
* NET 9372 = subckt_1658_sff1_x4.u
* NET 9373 = subckt_1658_sff1_x4.ckr
* NET 9374 = subckt_1658_sff1_x4.nckr
* NET 9375 = abc_11867_auto_rtlil_cc_2608_muxgate_11674
* NET 9376 = mos6502_cond_code[1]
* NET 9379 = abc_11867_new_n330
* NET 9382 = mos6502_cld
* NET 9384 = subckt_1664_sff1_x4.sff_s
* NET 9385 = subckt_1664_sff1_x4.y
* NET 9388 = subckt_1664_sff1_x4.sff_m
* NET 9389 = subckt_1664_sff1_x4.u
* NET 9390 = subckt_1664_sff1_x4.nckr
* NET 9391 = subckt_1664_sff1_x4.ckr
* NET 9392 = abc_11867_new_n1197
* NET 9394 = abc_11867_auto_rtlil_cc_2608_muxgate_11686
* NET 9395 = mos6502_load_reg
* NET 9397 = subckt_1698_sff1_x4.sff_s
* NET 9398 = subckt_1698_sff1_x4.y
* NET 9401 = subckt_1698_sff1_x4.sff_m
* NET 9402 = subckt_1698_sff1_x4.u
* NET 9403 = subckt_1698_sff1_x4.nckr
* NET 9404 = subckt_1698_sff1_x4.ckr
* NET 9405 = abc_11867_new_n437
* NET 9409 = abc_11867_new_n1323
* NET 9411 = abc_11867_auto_rtlil_cc_2608_muxgate_11742
* NET 9412 = abc_11867_new_n441
* NET 9417 = abc_11867_new_n1224
* NET 9418 = abc_11867_new_n1225
* NET 9419 = abc_11867_new_n462
* NET 9421 = abc_11867_new_n1198
* NET 9424 = abc_11867_new_n743
* NET 9426 = abc_11867_new_n672
* NET 9427 = abc_11867_new_n1326
* NET 9429 = abc_11867_new_n1289
* NET 9430 = abc_11867_new_n673
* NET 9432 = abc_11867_new_n454
* NET 9433 = abc_11867_new_n534_hfns_0
* NET 9475 = subckt_1742_sff1_x4.sff_s
* NET 9479 = subckt_1742_sff1_x4.y
* NET 9482 = subckt_1742_sff1_x4.sff_m
* NET 9483 = subckt_1742_sff1_x4.ckr
* NET 9484 = subckt_1742_sff1_x4.u
* NET 9485 = subckt_1742_sff1_x4.nckr
* NET 9486 = abc_11867_new_n407
* NET 9489 = mos6502_dihold[5]
* NET 9491 = subckt_1695_sff1_x4.sff_s
* NET 9493 = subckt_1695_sff1_x4.y
* NET 9497 = subckt_1695_sff1_x4.u
* NET 9498 = subckt_1695_sff1_x4.sff_m
* NET 9499 = subckt_1695_sff1_x4.ckr
* NET 9500 = subckt_1695_sff1_x4.nckr
* NET 9503 = abc_11867_new_n406
* NET 9505 = di[3]
* NET 9509 = abc_11867_new_n408
* NET 9513 = subckt_85_nmx2_x1.q
* NET 9514 = mos6502_dihold[3]
* NET 9516 = subckt_1693_sff1_x4.sff_s
* NET 9520 = subckt_1693_sff1_x4.y
* NET 9521 = subckt_1693_sff1_x4.sff_m
* NET 9523 = subckt_1693_sff1_x4.ckr
* NET 9524 = subckt_1693_sff1_x4.u
* NET 9525 = subckt_1693_sff1_x4.nckr
* NET 9526 = abc_11867_new_n1639
* NET 9532 = abc_11867_new_n1627
* NET 9533 = abc_11867_new_n1626
* NET 9540 = abc_11867_new_n1638
* NET 9541 = abc_11867_new_n1092
* NET 9547 = abc_11867_new_n1628
* NET 9552 = abc_11867_new_n340
* NET 9559 = abc_11867_new_n1078
* NET 9560 = abc_11867_new_n478_hfns_0
* NET 9566 = abc_11867_new_n338
* NET 9571 = abc_11867_new_n1591
* NET 9572 = abc_11867_new_n1589
* NET 9579 = abc_11867_new_n1588
* NET 9582 = abc_11867_new_n432_hfns_1
* NET 9586 = abc_11867_new_n1590
* NET 9594 = abc_11867_new_n1064
* NET 9597 = abc_11867_new_n428_hfns_1
* NET 9603 = abc_11867_new_n1071
* NET 9605 = abc_11867_new_n337
* NET 9609 = abc_11867_new_n971
* NET 9610 = abc_11867_new_n334
* NET 9612 = abc_11867_new_n412
* NET 9613 = abc_11867_new_n1050
* NET 9620 = subckt_81_nmx2_x1.q
* NET 9624 = abc_11867_new_n986
* NET 9633 = abc_11867_new_n420
* NET 9639 = abc_11867_new_n377
* NET 9642 = subckt_1707_sff1_x4.y
* NET 9643 = subckt_1707_sff1_x4.sff_s
* NET 9647 = subckt_1707_sff1_x4.sff_m
* NET 9648 = subckt_1707_sff1_x4.ckr
* NET 9649 = subckt_1707_sff1_x4.u
* NET 9650 = subckt_1707_sff1_x4.nckr
* NET 9667 = mos6502_sed
* NET 9669 = subckt_1665_sff1_x4.sff_s
* NET 9673 = subckt_1665_sff1_x4.y
* NET 9674 = subckt_1665_sff1_x4.sff_m
* NET 9676 = subckt_1665_sff1_x4.ckr
* NET 9677 = subckt_1665_sff1_x4.u
* NET 9678 = abc_11867_new_n1202
* NET 9679 = subckt_1665_sff1_x4.nckr
* NET 9680 = abc_11867_new_n1200
* NET 9682 = abc_11867_auto_rtlil_cc_2608_muxgate_11688
* NET 9686 = abc_11867_new_n1189
* NET 9688 = abc_11867_new_n393
* NET 9692 = abc_11867_new_n1194
* NET 9701 = abc_11867_new_n392
* NET 9702 = abc_11867_new_n1216
* NET 9710 = abc_11867_new_n1234
* NET 9716 = abc_11867_new_n447
* NET 9724 = abc_11867_new_n1242
* NET 9729 = abc_11867_new_n467
* NET 9732 = abc_11867_new_n1270
* NET 9743 = abc_11867_new_n1212
* NET 9746 = abc_11867_new_n1293
* NET 9747 = abc_11867_new_n440
* NET 9750 = abc_11867_new_n627
* NET 9760 = abc_11867_new_n1241
* NET 9916 = abc_11867_auto_rtlil_cc_2608_muxgate_11832
* NET 9922 = mos6502_pc[10]
* NET 9925 = abc_11867_new_n1640
* NET 9927 = abc_11867_new_n1587
* NET 9932 = abc_11867_new_n1072
* NET 9938 = abc_11867_new_n399
* NET 9939 = abc_11867_new_n398
* NET 9945 = abc_11867_new_n378
* NET 9946 = abc_11867_auto_rtlil_cc_2608_muxgate_11762
* NET 9947 = mos6502_irhold[7]
* NET 9955 = abc_11867_new_n416
* NET 9958 = abc_11867_new_n544
* NET 9971 = abc_11867_new_n1233
* NET 9972 = abc_11867_new_n1335
* NET 9974 = abc_11867_new_n752
* NET 9975 = abc_11867_new_n1334
* NET 9976 = abc_11867_new_n1199
* NET 9977 = abc_11867_new_n1302
* NET 9979 = abc_11867_new_n1324
* NET 9980 = abc_11867_new_n541
* NET 9984 = abc_11867_new_n1582
* NET 9985 = abc_11867_new_n1584
* NET 9986 = abc_11867_new_n1573
* NET 9987 = rdy_hfns_0
* NET 9989 = abc_11867_new_n1583
* NET 9991 = abc_11867_new_n1580
* NET 9993 = abc_11867_new_n1558
* NET 9994 = abc_11867_new_n1616
* NET 9996 = abc_11867_new_n1629
* NET 9997 = abc_11867_new_n1625
* NET 9998 = abc_11867_new_n1611
* NET 10000 = abc_11867_new_n1615
* NET 10002 = abc_11867_new_n1614
* NET 10003 = abc_11867_new_n1613
* NET 10004 = abc_11867_new_n1612
* NET 10005 = abc_11867_new_n1603
* NET 10006 = abc_11867_new_n1599
* NET 10008 = abc_11867_new_n1576
* NET 10009 = abc_11867_new_n1575
* NET 10011 = abc_11867_new_n1577
* NET 10013 = abc_11867_new_n1601
* NET 10014 = abc_11867_new_n1600
* NET 10015 = abc_11867_new_n1602
* NET 10017 = abc_11867_new_n1057
* NET 10018 = abc_11867_new_n619_hfns_0
* NET 10019 = subckt_1694_sff1_x4.sff_s
* NET 10020 = mos6502_dihold[4]
* NET 10021 = subckt_1694_sff1_x4.y
* NET 10022 = subckt_1694_sff1_x4.sff_m
* NET 10023 = subckt_1694_sff1_x4.u
* NET 10024 = mos6502_dimux[4]
* NET 10025 = subckt_1694_sff1_x4.ckr
* NET 10026 = subckt_1694_sff1_x4.nckr
* NET 10027 = abc_11867_new_n432_hfns_0
* NET 10028 = abc_11867_new_n428_hfns_0
* NET 10029 = abc_11867_new_n478_hfns_2
* NET 10031 = abc_11867_new_n485_hfns_2
* NET 10032 = abc_11867_new_n1056
* NET 10033 = abc_11867_new_n1058
* NET 10034 = abc_11867_new_n1059
* NET 10036 = abc_11867_new_n436
* NET 10042 = abc_11867_new_n1049
* NET 10043 = abc_11867_new_n1051
* NET 10044 = abc_11867_new_n1052
* NET 10053 = subckt_1704_sff1_x4.sff_s
* NET 10054 = mos6502_irhold[4]
* NET 10055 = subckt_1704_sff1_x4.y
* NET 10056 = subckt_1704_sff1_x4.sff_m
* NET 10057 = subckt_1704_sff1_x4.nckr
* NET 10058 = subckt_1704_sff1_x4.u
* NET 10059 = abc_11867_auto_rtlil_cc_2608_muxgate_11756
* NET 10060 = subckt_1704_sff1_x4.ckr
* NET 10063 = subckt_1703_sff1_x4.sff_s
* NET 10064 = subckt_1703_sff1_x4.ckr
* NET 10065 = subckt_1703_sff1_x4.nckr
* NET 10066 = subckt_1703_sff1_x4.y
* NET 10067 = subckt_1703_sff1_x4.sff_m
* NET 10068 = subckt_1703_sff1_x4.u
* NET 10073 = abc_11867_new_n543
* NET 10074 = abc_11867_new_n1327
* NET 10075 = abc_11867_new_n1325
* NET 10078 = abc_11867_new_n542
* NET 10080 = abc_11867_new_n1280
* NET 10081 = do[4]
* NET 10083 = abc_11867_new_n438
* NET 10137 = abc_11867_new_n1630
* NET 10139 = abc_11867_new_n1087
* NET 10142 = abc_11867_new_n1074
* NET 10147 = abc_11867_new_n1060
* NET 10153 = subckt_1692_sff1_x4.y
* NET 10155 = subckt_1692_sff1_x4.sff_m
* NET 10156 = subckt_1692_sff1_x4.ckr
* NET 10158 = abc_11867_new_n1053
* NET 10164 = subckt_1706_sff1_x4.y
* NET 10166 = subckt_1706_sff1_x4.sff_m
* NET 10167 = subckt_1706_sff1_x4.ckr
* NET 10170 = abc_11867_new_n451
* NET 10171 = abc_11867_new_n1570
* NET 10172 = abc_11867_new_n1561
* NET 10176 = abc_11867_new_n1586
* NET 10177 = abc_11867_auto_rtlil_cc_2608_muxgate_11834
* NET 10179 = abc_11867_new_n1596
* NET 10182 = abc_11867_new_n1617
* NET 10184 = abc_11867_new_n1595
* NET 10186 = abc_11867_auto_rtlil_cc_2608_muxgate_11830
* NET 10194 = abc_11867_new_n1605
* NET 10197 = rdy_hfns_3
* NET 10200 = abc_11867_new_n1568
* NET 10206 = abc_11867_new_n1641
* NET 10212 = abc_11867_new_n1637
* NET 10213 = mos6502_pc[11]
* NET 10214 = abc_11867_new_n1624
* NET 10215 = abc_11867_new_n1592
* NET 10218 = abc_11867_new_n1593
* NET 10222 = abc_11867_new_n1578
* NET 10225 = abc_11867_new_n1574
* NET 10228 = abc_11867_new_n1086
* NET 10231 = mos6502_dimux[6]
* NET 10232 = abc_11867_new_n1084
* NET 10239 = abc_11867_new_n978
* NET 10247 = abc_11867_new_n1564
* NET 10248 = abc_11867_new_n1565
* NET 10249 = abc_11867_new_n1563
* NET 10255 = abc_11867_new_n994
* NET 10256 = abc_11867_new_n472
* NET 10257 = mos6502_dimux[7]
* NET 10258 = abc_11867_new_n507
* NET 10259 = abc_11867_new_n402
* NET 10267 = subckt_1692_sff1_x4.sff_s
* NET 10268 = mos6502_dihold[2]
* NET 10269 = abc_11867_new_n601
* NET 10271 = subckt_1692_sff1_x4.nckr
* NET 10272 = subckt_1692_sff1_x4.u
* NET 10273 = subckt_77_nmx2_x1.q
* NET 10279 = abc_11867_new_n1048
* NET 10288 = subckt_1706_sff1_x4.sff_s
* NET 10289 = mos6502_irhold[6]
* NET 10291 = subckt_1706_sff1_x4.nckr
* NET 10292 = abc_11867_auto_rtlil_cc_2608_muxgate_11760
* NET 10293 = subckt_1706_sff1_x4.u
* NET 10302 = abc_11867_new_n379
* NET 10312 = mos6502_dimux[5]
* NET 10323 = abc_11867_new_n400
* NET 10332 = abc_11867_new_n390
* NET 10348 = abc_11867_auto_rtlil_cc_2608_muxgate_11754
* NET 10350 = mos6502_irhold[3]
* NET 10366 = abc_11867_new_n404
* NET 10378 = abc_11867_new_n452
* NET 10382 = abc_11867_new_n1272
* NET 10392 = abc_11867_new_n1271
* NET 10395 = abc_11867_new_n444
* NET 10399 = abc_11867_new_n741
* NET 10408 = abc_11867_new_n1240
* NET 10414 = abc_11867_new_n453
* NET 10418 = abc_11867_new_n534_hfns_2
* NET 10419 = abc_11867_new_n534
* NET 10540 = abc_11867_new_n1571
* NET 10541 = abc_11867_new_n1557
* NET 10542 = abc_11867_new_n1569
* NET 10545 = abc_11867_new_n1607
* NET 10546 = abc_11867_new_n1618
* NET 10547 = abc_11867_new_n1594
* NET 10550 = abc_11867_new_n1633
* NET 10551 = abc_11867_new_n1631
* NET 10554 = abc_11867_new_n1604
* NET 10555 = abc_11867_new_n1606
* NET 10558 = abc_11867_new_n1645
* NET 10559 = abc_11867_new_n1632
* NET 10560 = abc_11867_new_n1644
* NET 10561 = abc_11867_new_n1635
* NET 10564 = abc_11867_new_n1477
* NET 10565 = abc_11867_new_n1579
* NET 10566 = abc_11867_new_n1581
* NET 10567 = mos6502_pc[9]
* NET 10568 = abc_11867_new_n360
* NET 10570 = abc_11867_new_n1642
* NET 10571 = abc_11867_new_n1643
* NET 10575 = abc_11867_new_n367
* NET 10576 = abc_11867_new_n1636
* NET 10577 = abc_11867_new_n1462
* NET 10578 = abc_11867_new_n1475
* NET 10582 = abc_11867_new_n1055
* NET 10583 = abc_11867_new_n361
* NET 10584 = abc_11867_new_n1094
* NET 10585 = abc_11867_new_n1091
* NET 10589 = abc_11867_new_n1088
* NET 10590 = abc_11867_new_n1083
* NET 10591 = abc_11867_new_n1093
* NET 10594 = mos6502_dimux[3]
* NET 10595 = abc_11867_new_n963
* NET 10596 = abc_11867_new_n964
* NET 10599 = abc_11867_new_n1080
* NET 10600 = abc_11867_new_n1077
* NET 10604 = abc_11867_new_n968_hfns_0
* NET 10605 = abc_11867_new_n1079
* NET 10606 = abc_11867_new_n480
* NET 10608 = abc_11867_new_n970
* NET 10610 = abc_11867_new_n1567
* NET 10611 = abc_11867_new_n1566
* NET 10613 = abc_11867_new_n1562
* NET 10614 = abc_11867_new_n1472
* NET 10615 = abc_11867_new_n576
* NET 10618 = abc_11867_new_n1069
* NET 10619 = abc_11867_new_n364
* NET 10620 = di[2]
* NET 10621 = abc_11867_new_n403
* NET 10623 = subckt_1690_sff1_x4.sff_s
* NET 10624 = subckt_1690_sff1_x4.y
* NET 10627 = subckt_1690_sff1_x4.sff_m
* NET 10628 = subckt_1690_sff1_x4.u
* NET 10629 = subckt_1690_sff1_x4.ckr
* NET 10630 = subckt_1690_sff1_x4.nckr
* NET 10631 = subckt_1727_sff1_x4.sff_s
* NET 10634 = subckt_1727_sff1_x4.y
* NET 10635 = subckt_1727_sff1_x4.sff_m
* NET 10637 = subckt_1727_sff1_x4.u
* NET 10638 = clk_root_bl_1
* NET 10639 = subckt_1727_sff1_x4.ckr
* NET 10640 = subckt_1727_sff1_x4.nckr
* NET 10641 = mos6502_abh[2]
* NET 10643 = subckt_1726_sff1_x4.sff_s
* NET 10644 = subckt_1726_sff1_x4.y
* NET 10646 = abc_11867_auto_rtlil_cc_2608_muxgate_11800
* NET 10648 = subckt_1726_sff1_x4.sff_m
* NET 10649 = subckt_1726_sff1_x4.u
* NET 10650 = subckt_1726_sff1_x4.ckr
* NET 10651 = subckt_1726_sff1_x4.nckr
* NET 10652 = mos6502_dihold[1]
* NET 10654 = subckt_1691_sff1_x4.sff_s
* NET 10655 = subckt_1691_sff1_x4.y
* NET 10658 = subckt_1691_sff1_x4.sff_m
* NET 10659 = subckt_1691_sff1_x4.u
* NET 10660 = subckt_1691_sff1_x4.ckr
* NET 10661 = subckt_1691_sff1_x4.nckr
* NET 10662 = mos6502_irhold[5]
* NET 10663 = subckt_1705_sff1_x4.sff_s
* NET 10665 = subckt_1705_sff1_x4.y
* NET 10666 = subckt_1705_sff1_x4.sff_m
* NET 10668 = abc_11867_auto_rtlil_cc_2608_muxgate_11758
* NET 10670 = subckt_1705_sff1_x4.u
* NET 10671 = subckt_1705_sff1_x4.ckr
* NET 10672 = subckt_1705_sff1_x4.nckr
* NET 10675 = abc_11867_new_n389
* NET 10680 = mos6502_dimux[1]
* NET 10684 = mos6502_irhold_valid
* NET 10686 = abc_11867_new_n435_hfns_3
* NET 10687 = abc_11867_new_n1181_hfns_0
* NET 10689 = abc_11867_new_n1193
* NET 10691 = abc_11867_new_n1213
* NET 10692 = abc_11867_new_n1329
* NET 10693 = abc_11867_new_n448
* NET 10694 = abc_11867_new_n742
* NET 10695 = abc_11867_new_n1328
* NET 10697 = abc_11867_new_n1180
* NET 10698 = abc_11867_new_n537
* NET 10699 = abc_11867_new_n539
* NET 10700 = abc_11867_new_n435_hfns_1
* NET 10701 = abc_11867_new_n463
* NET 10702 = abc_11867_new_n456
* NET 10704 = abc_11867_new_n455
* NET 10705 = abc_11867_new_n449
* NET 10706 = abc_11867_new_n1284
* NET 10707 = abc_11867_new_n1330
* NET 10708 = abc_11867_new_n435_hfns_0
* NET 10709 = abc_11867_new_n536
* NET 10710 = abc_11867_new_n442
* NET 10771 = mos6502_pc[13]
* NET 10772 = abc_11867_new_n365
* NET 10773 = abc_11867_new_n1623
* NET 10774 = rdy_hfns_2
* NET 10777 = abc_11867_new_n1610
* NET 10780 = abc_11867_new_n1620
* NET 10781 = abc_11867_auto_rtlil_cc_2608_muxgate_11838
* NET 10783 = abc_11867_new_n1619
* NET 10786 = abc_11867_new_n1621
* NET 10787 = subckt_1746_sff1_x4.sff_s
* NET 10789 = di[1]
* NET 10792 = subckt_1746_sff1_x4.y
* NET 10795 = subckt_1746_sff1_x4.sff_m
* NET 10796 = abc_11867_auto_rtlil_cc_2608_muxgate_11840
* NET 10797 = subckt_1746_sff1_x4.ckr
* NET 10798 = subckt_1746_sff1_x4.u
* NET 10799 = subckt_1746_sff1_x4.nckr
* NET 10800 = mos6502_pc[15]
* NET 10803 = subckt_1747_sff1_x4.sff_s
* NET 10804 = subckt_1747_sff1_x4.y
* NET 10807 = subckt_1747_sff1_x4.sff_m
* NET 10808 = abc_11867_auto_rtlil_cc_2608_muxgate_11842
* NET 10810 = subckt_1747_sff1_x4.u
* NET 10811 = subckt_1747_sff1_x4.ckr
* NET 10812 = subckt_1747_sff1_x4.nckr
* NET 10813 = subckt_1731_sff1_x4.sff_s
* NET 10815 = subckt_1731_sff1_x4.y
* NET 10819 = subckt_1731_sff1_x4.u
* NET 10820 = subckt_1731_sff1_x4.sff_m
* NET 10822 = subckt_1731_sff1_x4.ckr
* NET 10823 = subckt_1731_sff1_x4.nckr
* NET 10824 = abc_11867_auto_rtlil_cc_2608_muxgate_11810
* NET 10825 = mos6502_abh[7]
* NET 10832 = abc_11867_new_n1090
* NET 10836 = abc_11867_new_n1095
* NET 10838 = mos6502_pc[14]
* NET 10839 = abc_11867_new_n366
* NET 10841 = subckt_1730_sff1_x4.sff_s
* NET 10843 = subckt_1730_sff1_x4.y
* NET 10846 = subckt_1730_sff1_x4.sff_m
* NET 10847 = a[15]
* NET 10849 = subckt_1730_sff1_x4.u
* NET 10850 = subckt_1730_sff1_x4.ckr
* NET 10851 = subckt_1730_sff1_x4.nckr
* NET 10853 = abc_11867_auto_rtlil_cc_2608_muxgate_11808
* NET 10854 = mos6502_abh[6]
* NET 10861 = abc_11867_new_n1076
* NET 10865 = abc_11867_new_n1081
* NET 10868 = subckt_1729_sff1_x4.sff_s
* NET 10869 = subckt_1729_sff1_x4.y
* NET 10873 = subckt_1729_sff1_x4.sff_m
* NET 10874 = subckt_1729_sff1_x4.ckr
* NET 10875 = subckt_1729_sff1_x4.u
* NET 10876 = subckt_1729_sff1_x4.nckr
* NET 10877 = a[14]
* NET 10879 = abc_11867_auto_rtlil_cc_2608_muxgate_11806
* NET 10880 = mos6502_abh[5]
* NET 10888 = abc_11867_new_n954_hfns_0
* NET 10890 = abc_11867_new_n362
* NET 10891 = abc_11867_new_n968_hfns_1
* NET 10892 = abc_11867_new_n975
* NET 10896 = abc_11867_new_n395
* NET 10897 = abc_11867_new_n1063
* NET 10899 = abc_11867_new_n1065
* NET 10900 = abc_11867_new_n1066
* NET 10901 = di[0]
* NET 10908 = abc_11867_new_n396
* NET 10909 = mos6502_dihold[0]
* NET 10912 = subckt_73_nmx2_x1.q
* NET 10913 = abc_11867_new_n394
* NET 10914 = clk_root_br_0
* NET 10915 = rdy_hfns_1
* NET 10917 = a[13]
* NET 10918 = abc_11867_new_n1067
* NET 10919 = abc_11867_new_n1062
* NET 10923 = abc_11867_auto_rtlil_cc_2608_muxgate_11802
* NET 10924 = mos6502_abh[3]
* NET 10934 = subckt_1728_sff1_x4.y
* NET 10935 = subckt_1728_sff1_x4.sff_s
* NET 10939 = subckt_1728_sff1_x4.sff_m
* NET 10940 = subckt_1728_sff1_x4.ckr
* NET 10941 = subckt_1728_sff1_x4.u
* NET 10942 = subckt_1728_sff1_x4.nckr
* NET 10944 = abc_11867_auto_rtlil_cc_2608_muxgate_11804
* NET 10945 = mos6502_abh[4]
* NET 10951 = a[12]
* NET 10959 = abc_11867_new_n1443
* NET 10963 = mos6502_abh[1]
* NET 10965 = subckt_1725_sff1_x4.sff_s
* NET 10969 = subckt_1725_sff1_x4.y
* NET 10970 = abc_11867_auto_rtlil_cc_2608_muxgate_11798
* NET 10971 = subckt_1725_sff1_x4.sff_m
* NET 10973 = subckt_1725_sff1_x4.ckr
* NET 10974 = subckt_1725_sff1_x4.u
* NET 10975 = subckt_1725_sff1_x4.nckr
* NET 10977 = a[11]
* NET 10979 = subckt_1700_sff1_x4.sff_s
* NET 10980 = subckt_1700_sff1_x4.y
* NET 10984 = subckt_1700_sff1_x4.sff_m
* NET 10985 = subckt_1700_sff1_x4.ckr
* NET 10986 = subckt_1700_sff1_x4.u
* NET 10987 = subckt_1700_sff1_x4.nckr
* NET 10989 = abc_11867_auto_rtlil_cc_2608_muxgate_11748
* NET 10990 = mos6502_irhold[0]
* NET 10995 = mos6502_dimux[0]
* NET 10999 = mos6502_irhold[1]
* NET 11001 = subckt_1701_sff1_x4.sff_s
* NET 11005 = subckt_1701_sff1_x4.y
* NET 11006 = abc_11867_auto_rtlil_cc_2608_muxgate_11750
* NET 11007 = subckt_1701_sff1_x4.sff_m
* NET 11009 = subckt_1701_sff1_x4.ckr
* NET 11010 = subckt_1701_sff1_x4.u
* NET 11011 = subckt_1701_sff1_x4.nckr
* NET 11012 = a[10]
* NET 11013 = abc_11867_new_n391
* NET 11018 = mos6502_dimux[2]
* NET 11019 = abc_11867_new_n1341
* NET 11024 = vdd
* NET 11026 = abc_11867_new_n435_hfns_4
* NET 11028 = mos6502_irhold[2]
* NET 11030 = subckt_1702_sff1_x4.sff_s
* NET 11032 = subckt_1702_sff1_x4.y
* NET 11035 = subckt_1702_sff1_x4.sff_m
* NET 11036 = abc_11867_auto_rtlil_cc_2608_muxgate_11752
* NET 11038 = subckt_1702_sff1_x4.u
* NET 11039 = a[9]
* NET 11040 = subckt_1702_sff1_x4.ckr
* NET 11041 = subckt_1702_sff1_x4.nckr
* NET 11042 = mos6502_store
* NET 11044 = subckt_1683_sff1_x4.sff_s
* NET 11048 = subckt_1683_sff1_x4.y
* NET 11049 = subckt_1683_sff1_x4.sff_m
* NET 11051 = clk_root_bl_0
* NET 11052 = subckt_1683_sff1_x4.ckr
* NET 11053 = subckt_1683_sff1_x4.u
* NET 11054 = abc_11867_new_n1287
* NET 11056 = subckt_1683_sff1_x4.nckr
* NET 11057 = abc_11867_new_n1285
* NET 11058 = abc_11867_new_n1286
* NET 11059 = abc_11867_auto_rtlil_cc_2608_muxgate_11726
* NET 11061 = abc_11867_new_n1331
* NET 11063 = abc_11867_new_n1333
* NET 11066 = abc_11867_new_n1211
* NET 11067 = abc_11867_new_n1301
* NET 11071 = abc_11867_new_n1332
* NET 11072 = abc_11867_new_n435_hfns_2
* NET 11074 = vss
* NET 11075 = abc_11867_new_n450
* NET 11076 = abc_11867_new_n445
* NET 11077 = abc_11867_new_n466
Mtr_16868 11024 10011 10010 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16867 10010 10008 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16866 11024 10009 10010 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16865 10222 10010 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16864 11024 875 876 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16863 875 1268 781 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16862 780 880 875 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16861 11024 1268 880 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16860 781 4910 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16859 11024 901 780 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16858 876 875 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16857 11024 325 320 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16856 325 1268 272 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16855 271 328 325 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16854 11024 1268 328 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16853 272 4905 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16852 11024 338 271 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16851 320 325 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16850 4665 7711 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16849 4665 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16848 11024 5898 4665 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16847 11024 9408 9405 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16846 9408 10684 9407 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16845 9406 9410 9408 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16844 11024 10684 9410 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16843 9407 9612 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16842 11024 9688 9406 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16841 9405 9408 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16840 11024 9698 10083 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16839 9698 10684 9457 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16838 9456 9700 9698 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16837 11024 10684 9700 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16836 9457 10024 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16835 11024 10054 9456 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16834 10083 9698 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16833 2158 8126 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16832 2158 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16831 11024 7721 2158 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16830 11024 9597 2158 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16829 11024 1973 1800 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16828 1800 2384 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16827 11024 2403 1800 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16826 1802 1800 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16825 5047 5100 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16824 5097 5094 5047 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16823 11024 5503 5097 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16822 9077 9732 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16821 11024 9743 9077 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16820 9074 9077 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16819 8384 10036 8183 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16818 8183 9419 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16817 11024 8970 8384 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16816 8395 8384 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16815 10690 11066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16814 11024 10689 10690 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16813 10691 10690 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16812 5508 5541 5509 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16811 5506 10604 5508 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16810 5507 10892 5506 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16809 11024 10888 5507 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16808 5504 5509 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16807 11024 6277 3866 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16806 3866 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16805 3866 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16804 11024 8839 3866 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16803 3860 3866 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16802 7035 7471 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16801 11024 7031 7035 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16800 7033 7035 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16799 11024 1793 116 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16798 6376 2636 117 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16797 117 1793 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16796 117 116 6376 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16795 11024 115 117 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16794 115 2636 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16793 10174 10540 10084 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16792 11024 10172 10084 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16791 10084 10171 10174 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16790 10186 10174 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16789 3345 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16788 11024 8126 3345 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16787 3967 3345 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16786 1286 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16785 11024 7721 1286 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16784 1861 1286 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16783 6439 7437 6294 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16782 6294 9333 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16781 11024 9321 6439 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16780 6437 6439 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16779 755 756 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16778 1040 1042 755 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16777 11024 1873 1040 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16776 6500 6498 6304 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16775 6304 6497 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16774 11024 6499 6500 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16773 6847 6500 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16772 11024 8430 7791 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16771 7791 8431 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16770 7791 8443 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16769 11024 10697 7791 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16768 7786 7791 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16767 6920 10891 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16766 7050 8091 6920 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16765 11024 8918 7050 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16764 4046 6173 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16763 11024 4183 4046 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16762 4043 4046 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16761 11024 9309 6794 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16760 6794 9560 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16759 11024 8921 6794 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16758 8091 6794 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16757 7854 10083 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16756 11024 10700 7854 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16755 7852 7854 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16754 11024 4701 4355 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16753 4355 4354 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16752 4355 5873 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16751 11024 4700 4355 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16750 5313 4355 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16749 11024 5600 2757 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16748 2757 6277 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16747 11024 3413 2757 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16746 2753 2757 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16745 11024 750 221 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16744 221 753 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16743 11024 1871 221 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16742 219 221 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16741 6149 6236 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16740 6147 6237 6234 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16739 11024 6476 6147 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16738 6237 6239 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16737 11024 8048 6239 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16736 11024 6478 6236 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16735 6235 6237 6149 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16734 6148 6239 6235 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16733 11024 6238 6148 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16732 6238 6235 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16731 6234 6239 6238 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16730 11024 6234 6476 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16729 6476 6234 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16728 11024 9314 7683 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16727 7683 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16726 11024 7678 7683 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16725 10615 7683 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16724 2166 2578 1362 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16723 1361 3714 2166 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16722 11024 2741 1361 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16721 1362 4014 11024 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16720 11024 10073 8747 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16719 8747 9419 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16718 11024 10708 8747 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16717 8746 8747 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16716 11024 7721 3087 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16715 3087 5898 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16714 3087 7514 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16713 11024 5293 3087 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16712 3086 3087 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16711 11024 5583 4690 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16710 4690 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16709 4690 9560 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16708 11024 7678 4690 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16707 5008 4690 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16706 3170 3188 3106 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16705 3106 3617 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16704 11024 3606 3170 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16703 3612 3170 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16702 11024 8424 8088 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16701 8016 8088 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16700 11024 8088 8016 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16699 11024 8088 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16698 11024 8088 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16697 11024 8145 8087 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16696 8015 8087 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16695 11024 8087 8015 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16694 11024 8087 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16693 11024 8087 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16692 11024 8424 2775 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16691 5262 2775 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16690 11024 2775 5262 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16689 11024 2775 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16688 11024 2775 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16687 11024 8424 2771 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16686 2773 2771 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16685 11024 2771 2773 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16684 11024 2771 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16683 11024 2771 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16682 11024 8424 2484 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16681 2483 2484 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16680 11024 2484 2483 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16679 11024 2484 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16678 11024 2484 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16677 11024 8145 2482 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16676 2481 2482 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16675 11024 2482 2481 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16674 11024 2482 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16673 11024 2482 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16672 11024 8424 2676 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16671 5083 2676 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16670 11024 2676 5083 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16669 11024 2676 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16668 11024 2676 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16667 11024 8424 2674 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16666 2673 2674 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16665 11024 2674 2673 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16664 11024 2674 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16663 11024 2674 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16662 11024 8424 2422 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16661 2446 2422 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16660 11024 2422 2446 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16659 11024 2422 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16658 11024 2422 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16657 11024 8145 2421 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16656 2420 2421 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16655 11024 2421 2420 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16654 11024 2421 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16653 11024 2421 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16652 8186 8460 8185 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16651 8185 9103 8463 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16650 8463 9107 8186 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16649 8186 9750 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16648 11024 9087 8186 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16647 8459 8463 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16646 11024 244 243 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16645 242 243 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16644 11024 2373 242 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16643 241 242 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16642 11024 242 241 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16641 11024 2799 2547 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16640 2547 2796 4359 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16639 675 678 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16638 671 677 672 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16637 11024 901 671 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16636 677 679 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16635 11024 2673 679 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16634 11024 876 678 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16633 676 677 675 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16632 674 679 676 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16631 11024 673 674 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16630 673 676 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16629 672 679 673 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16628 11024 672 901 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16627 901 672 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16626 9443 9524 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16625 9441 9523 9516 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16624 11024 9514 9441 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16623 9523 9525 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16622 11024 10914 9525 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16621 11024 10594 9524 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16620 9521 9523 9443 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16619 9442 9525 9521 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16618 11024 9520 9442 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16617 9520 9521 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16616 9516 9525 9520 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16615 11024 9516 9514 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16614 9514 9516 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16613 2003 5501 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16612 11024 2000 2003 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16611 1344 1495 1345 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16610 1345 1494 1488 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16609 1488 1493 1345 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16608 1344 1490 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16607 11024 1489 1344 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16606 1345 1496 1344 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16605 1834 1488 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16604 10086 10184 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16603 10783 10194 10086 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16602 11024 10182 10783 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16601 3817 10257 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16600 3817 5728 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16599 11024 5727 3817 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16598 9448 9649 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16597 9446 9648 9643 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16596 11024 9947 9446 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16595 9648 9650 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16594 11024 10638 9650 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16593 11024 9946 9649 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16592 9647 9648 9448 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16591 9447 9650 9647 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16590 11024 9642 9447 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16589 9642 9647 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16588 9643 9650 9642 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16587 11024 9643 9947 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16586 9947 9643 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16585 10598 10595 10597 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16584 10597 10596 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16583 11024 10594 10598 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16582 10897 10598 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16581 11012 10147 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16580 11024 10582 11012 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16579 4476 4363 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16578 11024 4364 4476 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16577 1355 4014 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16576 1557 3057 1355 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16575 1354 1556 1557 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16574 11024 3714 1354 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16573 2776 1557 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16572 6818 8318 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16571 6817 8316 6818 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16570 11024 8691 6817 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16569 10715 10798 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16568 10713 10797 10787 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16567 11024 10838 10713 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16566 10797 10799 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16565 11024 10914 10799 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16564 11024 10796 10798 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16563 10795 10797 10715 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16562 10714 10799 10795 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16561 11024 10792 10714 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16560 10792 10795 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16559 10787 10799 10792 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16558 11024 10787 10838 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16557 10838 10787 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16556 7535 7534 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16555 7535 7538 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16554 11024 7539 7535 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16553 11024 10697 7535 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16552 9686 10700 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16551 9686 10709 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16550 11024 10083 9686 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16549 1302 3735 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16548 11024 9597 1302 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16547 11024 2166 1946 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16546 1944 2167 2597 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16545 1945 2165 1944 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16544 1946 2581 1945 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16543 11024 2209 1948 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16542 1949 2211 2491 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16541 1950 2212 1949 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16540 1948 2208 1950 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16539 4280 4916 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16538 11024 4926 4280 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16537 4279 4280 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16536 8669 8671 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16535 8665 8672 8664 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16534 11024 8694 8665 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16533 8672 8673 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16532 11024 10914 8673 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16531 11024 8670 8671 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16530 8668 8672 8669 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16529 8666 8673 8668 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16528 11024 8667 8666 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16527 8667 8668 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16526 8664 8673 8667 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16525 11024 8664 8694 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16524 8694 8664 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16523 3682 3685 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16522 3678 3686 3679 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16521 11024 8297 3678 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16520 3686 3687 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16519 11024 5083 3687 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16518 11024 3684 3685 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16517 3683 3686 3682 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16516 3681 3687 3683 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16515 11024 3680 3681 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16514 3680 3683 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16513 3679 3687 3680 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16512 11024 3679 8297 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16511 8297 3679 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16510 8264 9290 8162 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16509 8162 8262 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16508 11024 9987 8264 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16507 8261 8264 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16506 7458 7685 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16505 11024 7457 7458 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16504 7670 7458 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16503 7567 7701 7566 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16502 7566 7719 7697 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16501 7697 7702 7567 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16500 7567 7695 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16499 11024 7704 7567 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16498 8327 7697 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16497 7539 9433 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16496 7539 9421 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16495 11024 9057 7539 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16494 11024 9716 7539 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16493 9046 9716 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16492 9046 10697 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16491 11024 9433 9046 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16490 11039 10158 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16489 11024 10279 11039 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16488 10693 11072 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16487 10693 10395 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16486 11024 10710 10693 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16485 11024 4631 4315 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16484 4315 4952 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16483 11024 4955 4315 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16482 4314 4315 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16481 1804 2403 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16480 1804 1973 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16479 11024 2384 1804 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16478 1808 7426 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16477 11024 1810 1808 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16476 2393 1808 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16475 5147 6214 5056 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16474 11024 6213 5056 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16473 5056 6215 5147 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16472 5148 5147 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16471 4589 5159 4387 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16470 11024 6213 4387 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16469 4387 6127 4589 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16468 4587 4589 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16467 6892 7535 6893 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16466 6893 8459 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16465 11024 6890 6892 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16464 6891 6892 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16463 7177 10399 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16462 7177 11066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16461 11024 9083 7177 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16460 11024 9716 7177 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16459 7784 8426 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16458 7784 8049 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16457 11024 8429 7784 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16456 8753 9051 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16455 8753 9418 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16454 11024 9073 8753 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16453 3375 4349 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16452 3375 3069 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16451 11024 3068 3375 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16450 7530 7534 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16449 11024 10697 7530 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16448 7531 7530 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16447 9417 11072 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16446 9417 10073 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16445 11024 10698 9417 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16444 11024 6764 6408 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16443 6413 9566 6291 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16442 6291 6764 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16441 6291 6408 6413 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16440 11024 6409 6291 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16439 6409 9566 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16438 5026 5610 5027 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16437 5025 5286 5026 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16436 11024 5024 5025 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16435 5023 5027 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16434 11024 4250 4251 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16433 4251 5023 4371 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16432 4374 4371 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16431 10703 10706 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16430 11024 10702 10703 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16429 11057 10703 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16428 11024 9702 8450 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16427 8450 9080 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16426 11024 9057 8450 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16425 8728 8450 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16424 10217 10577 10093 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16423 10093 10578 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16422 11024 10838 10217 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16421 10214 10217 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16420 11024 4950 4951 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16419 6205 4948 4949 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16418 4949 4950 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16417 4949 4951 6205 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16416 11024 4947 4949 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16415 4947 4948 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16414 11024 4352 4008 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16413 10028 4008 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16412 11024 4008 10028 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16411 11024 4008 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16410 11024 4008 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16409 11024 4352 1066 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16408 9597 1066 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16407 11024 1066 9597 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16406 11024 1066 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16405 11024 1066 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16404 11024 4352 4353 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16403 8643 4353 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16402 11024 4353 8643 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16401 11024 4353 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16400 11024 4353 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16399 11024 4352 3361 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16398 9308 3361 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16397 11024 3361 9308 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16396 11024 3361 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16395 11024 3361 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16394 11024 4352 4346 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16393 8921 4346 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16392 11024 4346 8921 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16391 11024 4346 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16390 11024 4346 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16389 11024 487 486 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16388 4352 486 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16387 11024 486 4352 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16386 11024 486 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16385 11024 486 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16384 11024 5275 4351 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16383 4351 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16382 4349 4694 4351 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16381 4350 4347 4349 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16380 4351 4348 4350 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16379 5310 5307 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16378 11024 5897 5310 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16377 5309 5310 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16376 11024 1601 1599 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16375 5293 1599 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16374 11024 1599 5293 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16373 11024 1599 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16372 11024 1599 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16371 11024 1601 1602 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16370 5607 1602 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16369 11024 1602 5607 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16368 11024 1602 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16367 11024 1602 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16366 11024 1308 1309 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16365 1601 1309 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16364 11024 1309 1601 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16363 11024 1309 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16362 11024 1309 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16361 11024 9287 9291 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16360 11024 10197 9289 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16359 9291 9289 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16358 11024 482 214 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16357 214 747 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16356 11024 219 214 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16355 437 214 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16354 11024 9560 3027 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16353 3027 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16352 3027 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16351 11024 8305 3027 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16350 3028 3027 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16349 11024 3969 3786 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16348 3786 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16347 9609 9308 3786 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16346 3785 3974 9609 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16345 3786 3967 3785 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16344 11024 3403 3406 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16343 3406 3402 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16342 11024 4043 3406 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16341 4054 3406 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16340 6432 7437 6292 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16339 6292 9566 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16338 11024 9310 6432 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16337 6431 6432 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16336 8041 8133 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16335 8039 8134 8130 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16334 11024 8725 8039 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16333 8134 8135 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16332 11024 10638 8135 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16331 11024 8724 8133 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16330 8132 8134 8041 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16329 8040 8135 8132 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16328 11024 8131 8040 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16327 8131 8132 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16326 8130 8135 8131 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16325 11024 8130 8725 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16324 8725 8130 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16323 6937 7161 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16322 7144 9046 6937 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16321 11024 7142 7144 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16320 11024 6759 6388 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16319 6402 8893 6289 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16318 6289 6759 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16317 6289 6388 6402 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16316 11024 6389 6289 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16315 6389 8893 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16314 11024 9560 1889 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16313 1889 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16312 1889 7678 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16311 11024 5293 1889 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16310 2172 1889 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16309 11024 5600 1593 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16308 1593 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16307 1593 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16306 11024 5293 1593 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16305 3082 1593 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16304 4959 5185 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16303 11024 5183 4959 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16302 4389 5175 4388 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16301 4388 4960 4603 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16300 4603 4952 4389 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16299 4389 5181 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16298 11024 5842 4389 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16297 4602 4603 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16296 262 395 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16295 260 394 388 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16294 11024 959 260 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16293 394 396 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16292 11024 2446 396 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16291 11024 963 395 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16290 393 394 262 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16289 261 396 393 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16288 11024 389 261 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16287 389 393 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16286 388 396 389 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16285 11024 388 959 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16284 959 388 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16283 6927 7104 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16282 6925 7106 7096 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16281 11024 7109 6925 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16280 7106 7105 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16279 11024 8048 7105 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16278 11024 7108 7104 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16277 7101 7106 6927 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16276 6926 7105 7101 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16275 11024 7099 6926 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16274 7099 7101 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16273 7096 7105 7099 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16272 11024 7096 7109 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16271 7109 7096 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16270 7470 8644 7469 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16269 7469 9610 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16268 11024 7468 7470 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16267 7467 7470 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16266 8206 8885 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16265 11024 9033 8206 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16264 9028 8733 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16263 11024 8411 9028 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16262 6283 6901 6178 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16261 6178 6286 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16260 11024 6282 6283 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16259 6177 6283 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16258 5647 6286 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16257 5931 6905 5647 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16256 11024 5933 5931 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16255 4726 4723 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16254 11024 4472 4726 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16253 5183 5181 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16252 11024 6246 5183 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16251 3844 7432 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16250 11024 2989 3844 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16249 4299 4942 4300 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16248 4300 4301 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16247 11024 4940 4299 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16246 4298 4299 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16245 8050 10689 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16244 11024 8746 8050 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16243 7520 8733 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16242 11024 7516 7520 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16241 7525 9083 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16240 11024 8746 7525 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16239 7517 8733 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16238 11024 7117 7517 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16237 7850 8063 7577 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16236 7577 10704 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16235 11024 8062 7850 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16234 7848 7850 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16233 5037 5312 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16232 11024 5038 5037 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16231 4472 4478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16230 11024 4369 4472 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16229 747 1545 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16228 11024 8713 747 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16227 8013 8082 8011 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16226 8086 10567 8013 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16225 8013 8635 8086 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16224 8011 8636 8013 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16223 8011 8930 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16222 11024 8633 8011 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16221 2637 2630 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16220 11024 2385 2637 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16219 10647 10649 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16218 10642 10650 10643 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16217 11024 10641 10642 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16216 10650 10651 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16215 11024 11051 10651 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16214 11024 10646 10649 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16213 10648 10650 10647 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16212 10645 10651 10648 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16211 11024 10644 10645 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16210 10644 10648 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16209 10643 10651 10644 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16208 11024 10643 10641 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16207 10641 10643 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16206 7419 7418 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16205 7419 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16204 11024 10027 7419 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16203 812 1300 1038 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16202 813 1040 812 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16201 11024 1301 813 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16200 1288 1038 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16199 9461 9566 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16198 10900 9609 9461 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16197 11024 9594 10900 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16196 2121 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16195 2121 8661 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16194 11024 6276 2121 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16193 8052 10701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16192 11024 11072 8052 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16191 5892 6895 5643 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16190 5643 6286 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16189 11024 5890 5892 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16188 5891 5892 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_16187 9999 10000 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16186 11024 9998 9999 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16185 9994 9999 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16184 4317 4323 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16183 11024 5539 4317 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16182 4316 4317 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16181 10726 10849 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16180 10724 10850 10841 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16179 11024 10854 10724 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16178 10850 10851 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16177 11024 10914 10851 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_16176 11024 10853 10849 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16175 10846 10850 10726 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16174 10725 10851 10846 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16173 11024 10843 10725 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16172 10843 10846 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16171 10841 10851 10843 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16170 11024 10841 10854 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16169 10854 10841 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16168 7483 7740 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_16167 7486 10995 7482 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16166 7482 8709 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16165 11024 7481 7488 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16164 7488 7727 7485 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16163 7485 7483 7486 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16162 7486 7740 7487 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16161 7487 7484 7488 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16160 11024 8709 7481 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_16159 7480 7486 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16158 11024 689 690 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16157 689 1268 646 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16156 645 647 689 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16155 11024 1268 647 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16154 646 5510 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16153 11024 691 645 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16152 690 689 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16151 11024 1266 1265 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16150 1266 1268 1269 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16149 1267 1270 1266 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16148 11024 1268 1270 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16147 1269 5544 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16146 11024 1490 1267 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16145 1265 1266 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16144 11024 931 934 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16143 931 1268 793 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16142 792 937 931 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16141 11024 1268 937 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16140 793 5707 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16139 11024 951 792 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16138 934 931 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16137 11024 982 983 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16136 982 1268 802 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16135 801 988 982 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16134 11024 1268 988 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16133 802 5732 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16132 11024 984 801 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16131 983 982 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16130 11024 374 368 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16129 374 1268 280 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16128 279 376 374 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16127 11024 1268 376 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16126 280 5531 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16125 11024 706 279 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16124 368 374 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16123 7068 5898 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16122 7068 8661 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16121 11024 6276 7068 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16120 1877 2763 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16119 11024 4325 1877 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16118 10003 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16117 10003 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16116 11024 9309 10003 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16115 11024 9304 10003 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16114 2995 2996 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16113 11024 4410 2995 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16112 3202 2995 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16111 9928 10614 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16110 9927 10615 9928 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16109 11024 10594 9927 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16108 11024 7684 7464 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16107 7464 7685 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16106 11024 7465 7464 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16105 7463 7464 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16104 11024 402 397 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16103 402 1268 284 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16102 283 405 402 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16101 11024 1268 405 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16100 284 3277 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16099 11024 723 283 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16098 397 402 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16097 11024 1237 1235 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16096 1237 1841 1238 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16095 1236 1239 1237 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16094 11024 1841 1239 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16093 1238 4910 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16092 11024 1403 1236 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16091 1235 1237 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16090 11024 1387 1388 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16089 1387 1841 1324 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16088 1325 1395 1387 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16087 11024 1841 1395 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16086 1324 4905 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16085 11024 1396 1325 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16084 1388 1387 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16083 11024 1232 1230 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16082 1232 1841 1233 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16081 1231 1234 1232 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16080 11024 1841 1234 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16079 1233 5510 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16078 11024 1813 1231 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16077 1230 1232 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16076 6994 8122 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16075 6994 9313 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16074 11024 6992 6994 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16073 11024 7655 6994 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16072 4666 7678 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16071 4666 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16070 11024 5719 4666 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16069 8244 9974 8190 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16068 8189 8475 8244 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16067 11024 9100 8189 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16066 8190 8477 11024 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16065 3074 4036 3073 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16064 3075 3071 3074 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16063 11024 3072 3075 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16062 5029 3073 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16061 5220 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16060 5220 5719 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16059 11024 7478 5220 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16058 11024 7739 5220 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16057 11024 5728 3842 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16056 3842 5727 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16055 11024 10231 3842 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16054 3837 3842 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16053 11024 5131 2510 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16052 2510 3618 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16051 2630 2971 2510 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16050 2509 5124 2630 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16049 2510 2967 2509 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16048 2582 2572 2478 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16047 2477 3714 2582 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16046 11024 8709 2477 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16045 2478 4014 11024 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_16044 9318 9320 9612 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16043 11024 10197 9320 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_16042 9319 10020 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16041 9612 10197 9319 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16040 11024 9316 9318 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16039 3798 4036 4041 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16038 3797 4037 3798 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16037 11024 4042 3797 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_16036 5018 4041 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16035 3223 3242 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_16034 3228 4936 3116 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16033 3116 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16032 11024 3216 3118 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16031 3118 3219 3117 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16030 3117 3223 3228 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16029 3228 3242 3119 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16028 3119 3889 3118 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16027 11024 4929 3216 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_16026 3651 3228 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16025 3209 3242 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_16024 3203 3198 3112 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16023 3112 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16022 11024 3199 3114 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16021 3114 3202 3113 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16020 3113 3209 3203 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16019 3203 3242 3115 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16018 3115 3884 3114 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_16017 11024 4929 3199 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_16016 4285 3203 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16015 11024 5764 5765 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16014 10891 5765 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16013 11024 5765 10891 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16012 11024 5765 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16011 11024 5765 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16010 11024 5168 5170 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16009 5764 5170 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16008 11024 5170 5764 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16007 11024 5170 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16006 11024 5170 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16005 11024 7721 7717 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16004 7717 7711 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16003 7717 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16002 11024 8725 7717 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_16001 8113 7717 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_16000 8776 8846 9955 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15999 11024 10197 8846 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15998 8775 9489 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15997 9955 10197 8775 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15996 11024 8840 8776 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15995 10770 11075 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15994 11077 11076 10770 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15993 11024 11072 11077 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15992 484 1545 289 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15991 289 4680 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15990 11024 4684 484 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15989 482 484 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15988 8085 8086 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15987 11024 8101 8085 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15986 8014 8085 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15985 1856 1857 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15984 11024 1855 1856 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15983 5557 1856 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15982 11024 5764 5540 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15981 10604 5540 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15980 11024 5540 10604 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15979 11024 5540 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15978 11024 5540 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15977 11024 6992 6988 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15976 7007 8122 6915 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15975 6915 6992 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15974 6915 6988 7007 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15973 11024 6983 6915 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15972 6983 8122 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15971 8002 10269 8001 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15970 8001 10256 8068 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15969 8068 10258 8002 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15968 8002 8620 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15967 11024 8621 8002 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15966 8000 8068 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15965 693 1495 695 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15964 695 1494 694 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15963 694 916 695 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15962 693 691 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15961 11024 1489 693 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15960 695 692 693 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15959 2412 694 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15958 9322 9347 9324 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15957 9324 9612 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15956 11024 9603 9322 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15955 9321 9322 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15954 3648 3647 3650 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15953 3650 3879 3649 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15952 3649 5131 3650 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15951 3648 3652 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15950 11024 4290 3648 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15949 3650 3646 3648 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15948 3872 3649 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15947 11024 2964 1795 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15946 1793 2962 1794 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15945 1794 2964 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15944 1794 1795 1793 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15943 11024 1792 1794 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15942 1792 2962 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15941 11024 6815 6463 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15940 10018 6463 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15939 11024 6463 10018 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15938 11024 6463 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15937 11024 6463 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15936 11024 6815 6816 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15935 7615 6816 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15934 11024 6816 7615 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15933 11024 6816 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15932 11024 6816 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15931 11024 6228 6229 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15930 6815 6229 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15929 11024 6229 6815 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15928 11024 6229 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15927 11024 6229 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15926 11024 8753 8148 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15925 8148 8430 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15924 11024 8443 8148 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15923 8049 8148 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15922 10052 10073 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15921 11024 10708 10052 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15920 9958 10052 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15919 3622 4567 3623 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15918 3623 3837 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15917 11024 4553 3622 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15916 3621 3622 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15915 4927 5140 4928 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15914 4928 4925 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15913 11024 4926 4927 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15912 5128 4927 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15911 5228 5226 5061 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15910 5061 5229 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15909 11024 9987 5228 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15908 6497 5228 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15907 8786 8893 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15906 10584 9609 8786 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15905 11024 9541 10584 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15904 7407 10269 7406 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15903 7406 10256 7405 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15902 7405 10258 7407 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15901 7407 7404 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15900 11024 7583 7407 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15899 7403 7405 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15898 1876 2138 1875 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15897 1875 2140 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15896 11024 1873 1876 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15895 1874 1876 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15894 11024 3092 291 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15893 291 8124 770 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15892 5129 5128 5054 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15891 5054 5132 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15890 11024 5681 5129 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15889 5704 5129 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15888 2428 3009 2429 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15887 2429 3008 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15886 11024 2688 2428 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15885 3000 2428 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15884 4503 6195 4377 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15883 4377 5098 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15882 11024 4500 4503 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15881 4501 4503 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15880 265 415 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15879 263 414 407 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15878 11024 984 263 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15877 414 416 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15876 11024 2446 416 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15875 11024 983 415 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15874 412 414 265 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15873 264 416 412 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15872 11024 411 264 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15871 411 412 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15870 407 416 411 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15869 11024 407 984 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15868 984 407 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15867 6885 6887 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15866 6880 6886 6881 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15865 11024 6879 6880 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15864 6886 6888 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15863 11024 8048 6888 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15862 11024 6891 6887 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15861 6884 6886 6885 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15860 6883 6888 6884 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15859 11024 6882 6883 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15858 6882 6884 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15857 6881 6888 6882 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15856 11024 6881 6879 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15855 6879 6881 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15854 8812 9061 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15853 9047 9046 8812 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15852 11024 9044 9047 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15851 6301 6819 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15850 10036 6489 6301 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15849 11024 6490 10036 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15848 11024 3734 1903 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15847 1903 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15846 1903 5600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15845 11024 7711 1903 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15844 2209 1903 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15843 11024 5014 5016 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15842 5016 5015 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15841 5016 5908 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15840 11024 5891 5016 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15839 5033 5016 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15838 11024 7042 754 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15837 754 3033 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15836 754 1881 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15835 11024 1556 754 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15834 753 754 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15833 256 318 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15832 254 317 311 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15831 11024 338 254 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15830 317 319 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15829 11024 2673 319 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15828 11024 320 318 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15827 316 317 256 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15826 255 319 316 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15825 11024 312 255 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15824 312 316 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15823 311 319 312 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15822 11024 311 338 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15821 338 311 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15820 11024 9987 9983 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15819 9982 9983 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15818 11024 10213 9982 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15817 10176 9982 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15816 11024 9982 10176 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15815 10035 10606 9936 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15814 9936 10608 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15813 11024 10641 10035 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15812 10033 10035 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15811 3031 3032 3292 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15810 3030 3028 3031 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15809 11024 3029 3030 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15808 11024 4976 3779 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15807 3780 3958 4142 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15806 3781 3959 3780 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15805 3779 4979 3781 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15804 2970 2971 2969 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15803 2969 3628 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15802 11024 2967 2970 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15801 2968 2970 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15800 10040 10272 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15799 10038 10156 10267 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15798 11024 10268 10038 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15797 10156 10271 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15796 11024 10638 10271 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15795 11024 11018 10272 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15794 10155 10156 10040 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15793 10039 10271 10155 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15792 11024 10153 10039 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15791 10153 10155 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15790 10267 10271 10153 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15789 11024 10267 10268 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15788 10268 10267 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15787 6749 8612 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15786 11024 10915 6749 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15785 9393 9686 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15784 9394 9680 9393 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15783 11024 9392 9394 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15782 2024 5672 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15781 11024 1824 2024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15780 10049 10293 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15779 10047 10167 10288 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15778 11024 10289 10047 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15777 10167 10291 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15776 11024 11051 10291 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15775 11024 10292 10293 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15774 10166 10167 10049 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15773 10048 10291 10166 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15772 11024 10164 10048 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15771 10164 10166 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15770 10288 10291 10164 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15769 11024 10288 10289 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15768 10289 10288 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15767 6104 6186 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15766 6102 6187 6183 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15765 11024 10771 6102 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15764 6187 6188 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15763 11024 10914 6188 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15762 11024 10781 6186 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15761 6185 6187 6104 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15760 6103 6188 6185 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15759 11024 6184 6103 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15758 6184 6185 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15757 6183 6188 6184 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15756 11024 6183 10771 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15755 10771 6183 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15754 11071 11077 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15753 11071 11067 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15752 11024 11066 11071 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15751 10707 10700 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15750 10707 10709 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15749 11024 10701 10707 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15748 1552 3735 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15747 11024 3734 1552 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15746 1873 3735 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15745 11024 5599 1873 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15744 4328 4327 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15743 11024 8713 4328 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15742 4640 4328 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15741 5636 9566 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15740 5726 7437 5636 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15739 11024 9310 5726 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15738 4505 5098 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15737 11024 6195 4505 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15736 5094 4505 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15735 8800 8980 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15734 8798 8981 8971 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15733 11024 8970 8798 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15732 8981 8982 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15731 11024 10638 8982 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15730 11024 8977 8980 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15729 8979 8981 8800 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15728 8799 8982 8979 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15727 11024 8973 8799 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15726 8973 8979 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15725 8971 8982 8973 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15724 11024 8971 8970 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15723 8970 8971 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15722 11024 6274 6164 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15721 6274 10687 6165 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15720 6166 6167 6274 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15719 11024 10687 6167 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15718 6165 6894 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15717 11024 6163 6166 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15716 6164 6274 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15715 8732 8735 8734 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15714 11024 8733 8735 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15713 8736 10382 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15712 8734 8733 8736 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15711 11024 8731 8732 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15710 3263 3288 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15709 11024 6137 3263 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15708 11024 10546 10549 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15707 10549 10555 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15706 11024 10547 10549 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15705 10780 10549 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15704 9543 9541 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15703 11024 10018 9543 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15702 9540 9543 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15701 11024 10576 10573 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15700 10572 10573 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15699 11024 10570 10572 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15698 10571 10572 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15697 11024 10572 10571 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15696 4980 5216 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15695 11024 5564 4980 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15694 4979 4980 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15693 11024 3899 3893 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15692 3899 4584 3758 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15691 3757 3901 3899 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15690 11024 4584 3901 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15689 3758 4617 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15688 11024 4553 3757 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15687 3893 3899 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15686 9915 9985 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15685 9916 9989 9915 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15684 11024 9986 9916 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15683 10079 10080 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15682 11024 10170 10079 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15681 9979 10079 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15680 2523 2691 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15679 2693 2692 2523 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15678 11024 6132 2693 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15677 11024 3086 2546 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15676 2546 3088 2790 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15675 2796 2790 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15674 11024 4066 4069 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15673 4068 4069 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15672 11024 4070 4068 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15671 5035 4068 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15670 11024 4068 5035 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15669 11024 5008 5011 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15668 5011 5009 5010 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15667 5603 5010 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15666 3962 3306 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15665 3962 3311 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15664 11024 3322 3962 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15663 11024 5771 3962 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15662 10196 10564 10087 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15661 10087 10619 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15660 11024 10554 10196 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15659 10194 10196 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15658 6127 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15657 6127 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15656 11024 6277 6127 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15655 11024 8082 6127 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15654 11024 9087 8058 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15653 8058 9750 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15652 8056 9107 8058 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15651 8057 9103 8056 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15650 8058 8460 8057 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15649 8713 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15648 8713 7478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15647 11024 8126 8713 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15646 11024 9729 7576 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15645 7576 8060 7839 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15644 7837 7839 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15643 1925 2006 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15642 6791 2004 1925 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15641 11024 4325 6791 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15640 11024 2121 2120 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15639 2120 2470 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15638 2120 2480 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15637 11024 2578 2120 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15636 2119 2120 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15635 11024 7069 2726 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15634 2726 6221 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15633 2726 3057 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15632 11024 6220 2726 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15631 2727 2726 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15630 11024 4286 4283 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15629 4543 4285 4287 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15628 4287 4286 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15627 4287 4283 4543 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15626 11024 4284 4287 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15625 4284 4285 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15624 8630 8629 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15623 8856 9295 8630 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15622 11024 8627 8856 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15621 5502 6381 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15620 11024 5504 5502 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15619 5501 5502 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15618 6145 6455 6224 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15617 6144 10891 6145 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15616 6143 10892 6144 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15615 11024 10888 6143 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15614 6142 6224 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15613 7025 7451 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15612 11024 7023 7025 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15611 7022 7025 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15610 10739 10912 10908 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15609 11024 10915 10912 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15608 10740 10909 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15607 10908 10915 10740 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15606 11024 10901 10739 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15605 11024 3413 816 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15604 816 2473 1048 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15603 2474 1048 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15602 3800 4064 4065 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15601 3801 5304 3800 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15600 11024 4463 3801 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15599 4063 4065 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15598 3325 8661 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15597 11024 5600 3325 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15596 3698 3325 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15595 6222 6806 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15594 11024 6809 6222 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15593 6141 6222 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15592 8653 8652 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15591 11024 8650 8653 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15590 8651 8653 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15589 2743 2746 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15588 11024 2741 2743 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15587 3311 2743 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15586 3707 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15585 11024 5719 3707 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15584 4653 3707 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15583 11024 5919 5790 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15582 5790 10029 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15581 11024 8643 5790 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15580 8316 5790 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15579 11024 5313 5316 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15578 5316 5320 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15577 11024 6182 5316 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15576 5312 5316 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15575 11024 6192 6191 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15574 6106 6387 6107 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15573 6107 6192 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15572 6107 6191 6106 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15571 11024 6190 6107 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15570 6190 6387 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15569 11024 9560 5007 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15568 5007 7478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15567 11024 10028 5007 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15566 5273 5007 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15565 513 3092 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15564 11024 8124 513 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15563 510 513 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15562 9312 9347 9311 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15561 9311 9509 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15560 11024 9594 9312 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15559 9310 9312 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15558 1803 1802 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15557 1807 1801 1803 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15556 11024 2679 1807 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15555 3142 3423 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15554 3140 3422 3417 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15553 11024 3413 3140 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15552 3422 3424 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15551 11024 5262 3424 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15550 11024 5034 3423 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15549 3420 3422 3142 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15548 3141 3424 3420 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15547 11024 3416 3141 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15546 3416 3420 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15545 3417 3424 3416 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15544 11024 3417 3413 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15543 3413 3417 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15542 8143 8419 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15541 8137 8229 8410 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15540 11024 8411 8137 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15539 8229 8420 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15538 11024 10638 8420 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15537 11024 9030 8419 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15536 8228 8229 8143 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15535 8140 8420 8228 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15534 11024 8225 8140 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15533 8225 8228 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15532 8410 8420 8225 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15531 11024 8410 8411 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15530 8411 8410 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15529 11024 7098 4989 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15528 9987 4989 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15527 11024 4989 9987 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15526 11024 4989 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15525 11024 4989 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15524 11024 7098 5225 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15523 10915 5225 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15522 11024 5225 10915 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15521 11024 5225 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15520 11024 5225 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15519 11024 7098 7073 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15518 10774 7073 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15517 11024 7073 10774 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15516 11024 7073 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15515 11024 7073 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15514 11024 7098 7076 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15513 10197 7076 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15512 11024 7076 10197 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15511 11024 7076 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15510 11024 7076 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15509 11024 5611 5612 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15508 7098 5612 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15507 11024 5612 7098 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15506 11024 5612 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15505 11024 5612 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15504 11024 5600 2498 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15503 2498 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15502 2498 5719 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15501 11024 10028 2498 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15500 2499 2498 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15499 11024 2499 2501 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15498 2501 2500 2792 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15497 8814 9430 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15496 9100 9095 8814 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15495 11024 9747 9100 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15494 2495 6220 1883 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_15493 1882 3714 2495 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_15492 11024 1881 1882 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_15491 1883 4014 11024 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_15490 4954 5181 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15489 11024 7109 4954 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15488 268 434 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15487 266 435 428 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15486 11024 729 266 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15485 435 436 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15484 11024 5262 436 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15483 11024 743 434 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15482 432 435 268 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15481 267 436 432 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15480 11024 429 267 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15479 429 432 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15478 428 436 429 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15477 11024 428 729 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15476 729 428 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15475 10238 10595 10103 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15474 10103 10596 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15473 11024 10312 10238 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15472 10600 10238 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15471 11024 5898 2184 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15470 2184 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15469 2184 7514 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15468 11024 5293 2184 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15467 2590 2184 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15466 3924 3925 3775 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15465 3775 3945 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15464 11024 3922 3924 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15463 4948 3924 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15462 6156 6249 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15461 6154 6250 6245 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15460 11024 6246 6154 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15459 6250 6252 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15458 11024 8048 6252 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15457 11024 7131 6249 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15456 6248 6250 6156 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15455 6155 6252 6248 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15454 11024 6247 6155 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15453 6247 6248 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15452 6245 6252 6247 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15451 11024 6245 6246 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15450 6246 6245 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15449 7036 7037 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15448 7036 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15447 11024 10027 7036 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15446 8212 8709 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15445 11024 8713 8212 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15444 9678 10687 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15443 11024 9667 9678 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15442 9392 10687 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15441 11024 9382 9392 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15440 4338 5191 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15439 11024 5191 4337 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15438 4336 7484 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15437 11024 4336 4338 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15436 4338 4337 4339 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15435 4339 7484 4338 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15434 4335 4339 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15433 11024 4339 4335 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15432 5873 8051 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15431 11024 6574 5873 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15430 10752 10974 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15429 10750 10973 10965 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15428 11024 10963 10750 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15427 10973 10975 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15426 11024 11051 10975 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15425 11024 10970 10974 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15424 10971 10973 10752 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15423 10751 10975 10971 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15422 11024 10969 10751 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15421 10969 10971 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15420 10965 10975 10969 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15419 11024 10965 10963 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15418 10963 10965 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15417 8834 7465 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15416 8834 7684 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15415 11024 7685 8834 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15414 8750 10689 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15413 11024 9080 8750 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15412 11024 1006 1008 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15411 1006 1248 806 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15410 807 1009 1006 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15409 11024 1248 1009 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15408 806 5732 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15407 11024 1005 807 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15406 1008 1006 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15405 11024 5739 5732 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15404 5739 5736 5619 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15403 5618 5742 5739 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15402 11024 5736 5742 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15401 5619 6788 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15400 11024 11018 5618 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15399 5732 5739 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15398 6569 10704 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15397 11024 9716 6569 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15396 11024 5293 5072 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15395 5072 5275 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15394 5279 6278 5072 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15393 5071 10606 5279 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15392 5072 5273 5071 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15391 5542 6221 5543 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15390 11024 5541 5543 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15389 5543 6220 5542 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15388 5756 5542 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15387 2635 2982 2511 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15386 11024 3632 2511 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15385 2511 3625 2635 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15384 2632 2635 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15383 5524 6214 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15382 11024 6215 5524 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15381 5523 5524 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15380 2436 2434 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15379 4311 2435 2436 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15378 11024 2688 4311 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15377 4323 10995 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15376 4323 5728 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15375 11024 5727 4323 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15374 11024 5131 3774 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15373 3774 4316 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15372 3941 4307 3774 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15371 3773 5124 3941 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15370 3774 3917 3773 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15369 8003 8893 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15368 8835 8644 8003 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15367 11024 8070 8835 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15366 7436 7445 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15365 7633 7667 7436 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15364 11024 10774 7633 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15363 10127 10694 10126 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15362 10126 10693 10384 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15361 10384 10392 10127 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15360 10127 10700 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15359 11024 10701 10127 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15358 10382 10384 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15357 8042 9710 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15356 11024 8429 8042 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15355 11024 1842 1839 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15354 1842 1841 1843 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15353 1840 1845 1842 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15352 11024 1841 1845 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15351 1843 5544 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15350 11024 1844 1840 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15349 1839 1842 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15348 11024 1436 1437 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15347 1436 1841 1335 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15346 1334 1442 1436 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15345 11024 1841 1442 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15344 1335 5707 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15343 11024 1826 1334 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15342 1437 1436 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15341 6251 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15340 6251 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15339 11024 9560 6251 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15338 7465 8921 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15337 7465 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15336 11024 8922 7465 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15335 2572 5898 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15334 2572 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15333 11024 9560 2572 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15332 9432 10414 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15331 11024 10686 9432 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15330 5906 9560 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15329 5906 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15328 11024 5600 5906 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15327 11024 5599 5906 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15326 6176 10704 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15325 6176 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15324 11024 6574 6176 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15323 11024 7852 6176 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15322 8636 6221 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15321 11024 6220 8636 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15320 11024 10774 10779 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15319 10776 10779 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15318 11024 10838 10776 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15317 10773 10776 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15316 11024 10776 10773 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15315 5240 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15314 5240 6277 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15313 11024 7478 5240 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15312 11024 5851 5240 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15311 2990 7432 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15310 11024 2989 2990 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15309 3635 2990 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15308 3674 3945 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15307 11024 3925 3674 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15306 3675 3674 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15305 11024 10015 10012 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15304 10012 10013 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15303 11024 10014 10012 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15302 10005 10012 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15301 11024 10566 9990 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15300 9990 10542 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15299 11024 10541 9990 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15298 9989 9990 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15297 11024 1832 2047 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15296 1832 1841 1830 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15295 1831 1833 1832 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15294 11024 1841 1833 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15293 1830 5732 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15292 11024 2038 1831 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15291 2047 1832 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15290 11024 1263 1260 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15289 1263 1841 1262 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15288 1261 1264 1263 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15287 11024 1841 1264 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15286 1262 5531 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15285 11024 1456 1261 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15284 1260 1263 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15283 11024 1460 1461 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15282 1460 1841 1340 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15281 1339 1470 1460 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15280 11024 1841 1470 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15279 1340 3277 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15278 11024 2432 1339 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15277 1461 1460 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15276 11024 1241 1431 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15275 1241 1284 1242 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15274 1240 1243 1241 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15273 11024 1284 1243 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15272 1242 4910 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15271 11024 1423 1240 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15270 1431 1241 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15269 11024 353 347 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15268 353 1284 278 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15267 277 356 353 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15266 11024 1284 356 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15265 278 4905 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15264 11024 348 277 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15263 347 353 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15262 7069 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15261 7069 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15260 11024 6277 7069 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15259 11024 2172 1947 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15258 1947 2177 2174 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15257 2581 2174 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15256 3858 5150 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_15255 3854 3844 3752 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15254 3752 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15253 11024 3846 3754 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15252 3754 3849 3753 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15251 3753 3858 3854 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15250 3854 5150 3755 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15249 3755 4530 3754 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15248 11024 4929 3846 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_15247 4272 3854 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15246 3640 5150 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_15245 3642 3635 3639 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15244 3639 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15243 11024 3636 3643 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15242 3643 3637 3638 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15241 3638 3640 3642 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15240 3642 5150 3641 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15239 3641 4535 3643 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15238 11024 4929 3636 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_15237 4275 3642 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15236 11024 8709 7710 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15235 7710 8092 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15234 11024 8713 7710 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15233 7704 7710 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15232 11024 696 925 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15231 696 1284 649 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15230 648 650 696 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15229 11024 1284 650 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15228 649 5510 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15227 11024 916 648 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15226 925 696 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15225 11024 1283 1280 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15224 1283 1284 1281 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15223 1282 1285 1283 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15222 11024 1284 1285 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15221 1281 5544 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15220 11024 1493 1282 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15219 1280 1283 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15218 2470 6277 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15217 2470 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15216 11024 6275 2470 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15215 8477 9405 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15214 8477 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15213 11024 10710 8477 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15212 11024 10700 8477 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15211 6905 8746 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15210 6905 8059 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15209 11024 9057 6905 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15208 11024 9433 6905 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15207 7217 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15206 7217 9080 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15205 11024 8453 7217 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15204 11024 9433 7217 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15203 11024 6232 6227 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15202 6227 6457 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15201 6227 6251 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15200 11024 6230 6227 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15199 10578 6227 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15198 6540 7532 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15197 11024 6537 6540 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15196 6538 6540 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15195 6865 7798 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15194 11024 10697 6865 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15193 6866 6865 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15192 1507 1519 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15191 11024 10915 1507 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15190 1504 1507 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15189 10530 10619 10617 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15188 10531 10891 10530 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15187 10529 10892 10531 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15186 11024 10888 10529 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_15185 10618 10617 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15184 11024 5131 4945 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15183 4945 4944 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15182 4943 4942 4945 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15181 4941 5124 4943 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15180 4945 4940 4941 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15179 8641 9287 8640 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15178 11024 8645 8640 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15177 8640 8834 8641 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15176 8862 8641 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15175 6258 8733 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15174 11024 6259 6258 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15173 7129 6258 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15172 11024 489 237 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15171 5919 237 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15170 11024 237 5919 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15169 11024 237 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15168 11024 237 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15167 11024 489 490 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15166 2133 490 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15165 11024 490 2133 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15164 11024 490 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15163 11024 490 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15162 11024 238 236 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15161 489 236 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15160 11024 236 489 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15159 11024 236 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15158 11024 236 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15157 11024 2697 2437 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15156 10888 2437 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15155 11024 2437 10888 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15154 11024 2437 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15153 11024 2437 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15152 11024 2697 2698 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15151 6132 2698 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15150 11024 2698 6132 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15149 11024 2698 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15148 11024 2698 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15147 11024 2450 2438 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15146 2697 2438 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15145 11024 2438 2697 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15144 11024 2438 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15143 11024 2438 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15142 3992 5719 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15141 11024 7721 3992 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15140 4654 3992 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15139 1835 1834 1836 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15138 1836 1837 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15137 11024 2688 1835 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15136 5528 1835 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15135 8619 8617 8618 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15134 11024 8616 8618 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15133 8618 8834 8619 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15132 8824 8619 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15131 5820 9379 5642 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15130 5642 5818 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15129 11024 10684 5820 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15128 6498 5820 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15127 3132 3967 3131 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15126 3131 3974 3315 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15125 3315 9308 3132 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15124 3132 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15123 11024 3969 3132 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15122 3693 3315 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15121 10312 9955 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15120 10231 9633 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15119 9075 10701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15118 11024 11072 9075 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15117 9095 9075 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15116 11024 6278 3741 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15115 3741 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15114 3741 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15113 11024 7514 3741 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15112 4047 3741 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15111 11024 6243 1872 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15110 1872 2741 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15109 11024 2728 1872 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15108 1871 1872 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15107 11024 472 470 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15106 470 1545 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15105 11024 5837 470 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15104 466 470 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15103 2613 8821 2505 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15102 11024 2609 2505 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15101 2505 10545 2613 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15100 2610 2613 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15099 11024 5131 3645 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15098 3645 3879 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15097 4286 4290 3645 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15096 3644 5124 4286 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15095 3645 4285 3644 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15094 259 365 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15093 257 366 358 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15092 11024 706 257 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15091 366 367 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15090 11024 2673 367 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15089 11024 368 365 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15088 364 366 259 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15087 258 367 364 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15086 11024 360 258 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15085 360 364 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15084 358 367 360 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15083 11024 358 706 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15082 706 358 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15081 5590 5591 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15080 5585 5592 5586 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15079 11024 6163 5585 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15078 5592 5594 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15077 11024 8048 5594 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15076 11024 6164 5591 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15075 5589 5592 5590 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15074 5588 5594 5589 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15073 11024 5587 5588 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15072 5587 5589 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15071 5586 5594 5587 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15070 11024 5586 6163 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15069 6163 5586 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15068 11024 6413 6203 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15067 6117 6993 6118 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15066 6118 6413 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15065 6118 6203 6117 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15064 11024 6204 6118 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15063 6204 6993 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_15062 11024 9020 1305 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15061 1305 5600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15060 1305 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15059 11024 5293 1305 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15058 1574 1305 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15057 10024 9612 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15056 11024 7514 5596 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15055 5596 7478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15054 5596 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15053 11024 5607 5596 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15052 6574 5596 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15051 5166 7437 5058 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15050 5058 6803 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15049 11024 8937 5166 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15048 5165 5166 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15047 3614 4501 3613 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15046 3613 3612 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15045 11024 3610 3614 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15044 3611 3614 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_15043 685 686 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15042 681 687 680 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15041 11024 691 681 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15040 687 688 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15039 11024 2673 688 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15038 11024 690 686 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15037 684 687 685 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15036 682 688 684 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15035 11024 683 682 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15034 683 684 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15033 680 688 683 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15032 11024 680 691 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15031 691 680 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15030 10657 10659 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15029 10653 10660 10654 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15028 11024 10652 10653 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15027 10660 10661 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15026 11024 11051 10661 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15025 11024 10680 10659 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15024 10658 10660 10657 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15023 10656 10661 10658 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15022 11024 10655 10656 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15021 10655 10658 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15020 10654 10661 10655 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15019 11024 10654 10652 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15018 10652 10654 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15017 2717 5746 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15016 11024 2693 2717 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_15015 11024 5901 5645 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15014 5645 6861 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15013 5897 6574 5645 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15012 5644 7840 5897 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15011 5645 9424 5644 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_15010 10669 10670 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15009 10664 10671 10663 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15008 11024 10662 10664 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15007 10671 10672 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15006 11024 11051 10672 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_15005 11024 10668 10670 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15004 10666 10671 10669 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15003 10667 10672 10666 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15002 11024 10665 10667 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15001 10665 10666 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_15000 10663 10672 10665 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14999 11024 10663 10662 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14998 10662 10663 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14997 8309 8824 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14996 11024 8817 8309 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14995 3694 3693 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14994 11024 8297 3694 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14993 11024 3413 10256 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14992 11024 2473 481 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14991 10256 481 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14990 2688 1864 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14989 2688 1866 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14988 11024 2119 2688 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14987 11024 4554 4555 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14986 4554 5140 4383 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14985 4384 4561 4554 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14984 11024 5140 4561 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14983 4383 4617 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14982 11024 4553 4384 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14981 4555 4554 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14980 667 668 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14979 662 669 663 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14978 11024 4254 662 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14977 669 670 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14976 11024 5083 670 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14975 11024 2610 668 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14974 666 669 667 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14973 665 670 666 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14972 11024 664 665 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14971 664 666 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14970 663 670 664 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14969 11024 663 4254 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14968 4254 663 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14967 9581 9594 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14966 11024 10018 9581 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14965 9579 9581 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14964 11024 10826 10824 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14963 10826 10959 10723 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14962 10722 10835 10826 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14961 11024 10959 10835 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14960 10723 10847 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14959 11024 10825 10722 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14958 10824 10826 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14957 11024 10852 10853 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14956 10852 10959 10728 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14955 10727 10864 10852 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14954 11024 10959 10864 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14953 10728 10877 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14952 11024 10854 10727 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14951 10853 10852 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14950 11024 10878 10879 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14949 10878 10959 10733 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14948 10732 10887 10878 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14947 11024 10959 10887 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14946 10733 10917 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14945 11024 10880 10732 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14944 10879 10878 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14943 11024 10943 10944 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14942 10943 10959 10747 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14941 10746 10953 10943 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14940 11024 10959 10953 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14939 10747 10951 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14938 11024 10945 10746 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14937 10944 10943 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14936 11024 10922 10923 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14935 10922 10959 10742 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14934 10741 10931 10922 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14933 11024 10959 10931 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14932 10742 10977 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14931 11024 10924 10741 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14930 10923 10922 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14929 11024 10280 10646 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14928 10280 10959 10113 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14927 10112 10284 10280 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14926 11024 10959 10284 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14925 10113 11012 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14924 11024 10641 10112 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14923 10646 10280 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14922 4240 5086 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14921 11024 1401 4240 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14920 11024 6468 6451 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14919 11024 9987 6338 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14918 6451 6338 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14917 11024 2473 756 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14916 11024 3413 757 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14915 756 757 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14914 11024 3391 2781 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14913 2777 2781 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14912 11024 2776 2777 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14911 3069 2777 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14910 11024 2777 3069 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14909 3959 3035 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14908 3959 3036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14907 11024 3037 3959 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14906 2972 3830 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14905 11024 4926 2972 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14904 2971 2972 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14903 6215 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14902 6215 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14901 11024 7711 6215 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14900 11024 8848 6215 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14899 3158 5144 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14898 11024 3155 3158 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14897 11024 9298 9299 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14896 9299 9296 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14895 11024 9297 9299 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14894 9295 9299 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14893 11024 10954 10970 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14892 10954 10959 10749 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14891 10748 10962 10954 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14890 11024 10959 10962 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14889 10749 11039 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14888 11024 10963 10748 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14887 10970 10954 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14886 7798 10399 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14885 7798 11066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14884 11024 10689 7798 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14883 11024 9716 7798 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14882 11024 1552 1299 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14881 1299 5809 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14880 1299 7041 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14879 11024 2099 1299 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14878 1867 1299 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14877 11024 6275 5563 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14876 5563 10029 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14875 5563 7478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14874 11024 8409 5563 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14873 5816 5563 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14872 11024 5528 5530 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14871 5529 5530 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14870 11024 6437 5529 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14869 5527 5529 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14868 11024 5529 5527 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14867 11024 8833 8826 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14866 8826 8831 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14865 8826 8824 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14864 11024 8817 8826 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14863 10541 8826 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14862 8010 9566 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14861 8267 8644 8010 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14860 11024 8081 8267 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14859 7000 6998 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14858 11024 9605 7000 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14857 6997 7000 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14856 11024 3092 240 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14855 239 240 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14854 11024 8124 239 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14853 238 239 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14852 11024 239 238 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14851 11024 10709 10711 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14850 10711 10710 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14849 11024 10708 10711 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14848 11067 10711 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14847 2433 7701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14846 11024 2432 2433 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14845 3008 2433 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14844 1829 7701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14843 11024 2038 1829 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14842 2691 1829 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14841 11024 6201 5701 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14840 5698 5693 5634 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14839 5634 6201 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14838 5634 5701 5698 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14837 11024 5694 5634 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14836 5694 5693 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14835 5669 5670 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14834 11024 5665 5669 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14833 5667 5669 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14832 4698 5607 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14831 11024 6493 4698 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14830 4694 4698 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14829 3708 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14828 3994 5911 3708 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14827 11024 4654 3994 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14826 7433 7437 7434 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14825 7434 9552 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14824 11024 9300 7433 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14823 7432 7433 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14822 11024 6105 2423 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14821 6192 9305 2425 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14820 2425 6105 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14819 2425 2423 6192 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14818 11024 2424 2425 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14817 2424 9305 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14816 11024 10078 9425 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14815 9425 10698 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14814 11024 10708 9425 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14813 9430 9425 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14812 11024 5302 5305 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14811 5305 6179 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14810 11024 5908 5305 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14809 5295 5305 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14808 4373 4727 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14807 4367 4728 4724 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14806 11024 8124 4367 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14805 4728 4729 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14804 11024 5262 4729 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14803 11024 4726 4727 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14802 4484 4728 4373 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14801 4372 4729 4484 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14800 11024 4481 4372 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14799 4481 4484 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14798 4724 4729 4481 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14797 11024 4724 8124 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14796 8124 4724 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14795 11024 10774 7579 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14794 7580 7579 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14793 11024 10567 7580 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14792 10172 7580 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14791 11024 7580 10172 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14790 6525 8762 6306 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14789 6306 6866 6525 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14788 11024 6524 6306 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14787 10030 10606 9933 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14786 9933 10608 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14785 11024 10945 10030 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14784 9932 10030 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14783 11024 3076 3078 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14782 3078 3077 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14781 11024 4349 3078 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14780 4057 3078 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14779 11024 9020 1586 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14778 1586 5600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14777 1586 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14776 11024 5293 1586 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14775 1583 1586 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14774 11024 10704 6565 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14773 6565 9716 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14772 11024 9747 6565 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14771 6564 6565 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14770 11024 452 444 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14769 444 464 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14768 444 745 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14767 11024 460 444 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14766 7701 444 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14765 11024 4602 3776 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14764 3776 4142 3926 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14763 3925 3926 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14762 6936 7141 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14761 6934 7140 7132 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14760 11024 7516 6934 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14759 7140 7143 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14758 11024 8048 7143 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14757 11024 7521 7141 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14756 7139 7140 6936 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14755 6935 7143 7139 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14754 11024 7136 6935 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14753 7136 7139 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14752 7132 7143 7136 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14751 11024 7132 7516 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14750 7516 7132 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14749 11024 7478 2503 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14748 2503 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14747 2503 8126 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14746 11024 5607 2503 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14745 2601 2503 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14744 172 174 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14743 168 175 169 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14742 11024 708 168 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14741 175 176 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14740 11024 2673 176 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14739 11024 377 174 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14738 173 175 172 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14737 171 176 173 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14736 11024 170 171 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14735 170 173 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14734 169 176 170 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14733 11024 169 708 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14732 708 169 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14731 7493 7495 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14730 7489 7496 7490 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14729 11024 7749 7489 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14728 7496 7497 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14727 11024 10638 7497 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14726 11024 7752 7495 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14725 7494 7496 7493 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14724 7491 7497 7494 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14723 11024 7492 7491 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14722 7492 7494 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14721 7490 7497 7492 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14720 11024 7490 7749 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14719 7749 7490 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14718 5043 5081 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14717 5041 5085 5075 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14716 11024 5488 5041 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14715 5085 5084 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14714 11024 5083 5084 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14713 11024 5487 5081 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14712 5080 5085 5043 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14711 5042 5084 5080 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14710 11024 5076 5042 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14709 5076 5080 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14708 5075 5084 5076 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14707 11024 5075 5488 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14706 5488 5075 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14705 11019 6497 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14704 11024 6499 11019 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14703 8749 10687 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14702 11024 8748 8749 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14701 7813 9083 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14700 11024 9080 7813 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14699 5040 5321 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14698 11024 5934 5040 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14697 10556 10558 10516 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14696 11024 10561 10516 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14695 10516 10560 10556 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14694 10808 10556 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14693 11024 6545 5565 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14692 11024 8409 5566 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14691 5565 5566 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14690 4410 4617 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14689 11024 4553 4410 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14688 10013 8921 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14687 10013 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14686 11024 8922 10013 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14685 11024 8918 10013 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14684 1865 1862 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14683 1865 7711 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14682 11024 7721 1865 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14681 9411 9972 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14680 11024 9409 9411 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14679 8046 10687 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14678 11024 8407 8046 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14677 7142 8733 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14676 11024 6867 7142 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14675 11024 721 722 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14674 721 1248 652 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14673 651 653 721 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14672 11024 1248 653 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14671 652 5531 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14670 11024 711 651 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14669 722 721 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14668 8709 5898 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14667 8709 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14666 11024 8922 8709 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14665 10170 11075 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14664 11024 11072 10170 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14663 6182 8244 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14662 11024 6574 6182 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14661 2496 2788 2592 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14660 2497 2495 2496 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14659 11024 3079 2497 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14658 8635 7041 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14657 11024 7042 8635 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14656 2974 7426 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14655 11024 1810 2974 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14654 3128 3274 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14653 3126 3273 3267 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14652 11024 8305 3126 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14651 3273 3275 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14650 11024 5083 3275 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14649 11024 3272 3274 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14648 3270 3273 3128 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14647 3127 3275 3270 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14646 11024 3266 3127 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14645 3266 3270 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14644 3267 3275 3266 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14643 11024 3267 8305 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14642 8305 3267 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14641 10184 10542 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14640 10184 10218 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14639 11024 10566 10184 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14638 11024 10541 10184 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14637 9995 10564 9921 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14636 9921 10583 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14635 11024 10565 9995 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14634 9991 9995 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14633 11024 5534 5531 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14632 5534 5736 5532 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14631 5533 5536 5534 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14630 11024 5736 5536 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14629 5532 6449 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14628 11024 10680 5533 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14627 5531 5534 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14626 11024 198 195 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14625 198 1248 196 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14624 197 199 198 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14623 11024 1248 199 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14622 196 3277 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14621 11024 724 197 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14620 195 198 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14619 6123 10269 6122 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14618 6122 10256 6207 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14617 6207 10258 6123 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14616 6123 6210 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14615 11024 6451 6123 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14614 6121 6207 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14613 6230 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14612 6230 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14611 11024 5583 6230 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14610 11024 10268 10259 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14609 11024 10774 10146 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14608 10259 10146 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14607 4998 8921 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14606 4998 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14605 11024 7711 4998 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14604 11024 5293 4998 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14603 5001 9560 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14602 5001 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14601 11024 9309 5001 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14600 11024 8921 5001 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14599 5304 6177 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14598 11024 5926 5304 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14597 4463 5897 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14596 11024 6171 4463 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14595 3696 3695 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14594 11024 7484 3696 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14593 3958 3696 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14592 3883 5153 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14591 11024 5718 3883 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14590 3879 3883 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14589 4313 6811 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14588 11024 4311 4313 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14587 4312 4313 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14586 3663 3928 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14585 11024 4410 3663 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14584 3905 3663 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14583 8431 9418 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14582 11024 9417 8431 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14581 11024 960 963 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14580 960 1284 796 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14579 797 964 960 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14578 11024 1284 964 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14577 796 5707 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14576 11024 959 797 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14575 963 960 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14574 11024 742 743 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14573 742 1284 655 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14572 654 656 742 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14571 11024 1284 656 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14570 655 5732 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14569 11024 729 654 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14568 743 742 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14567 11024 383 377 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14566 383 1284 282 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14565 281 385 383 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14564 11024 1284 385 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14563 282 5531 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14562 11024 708 281 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14561 377 383 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14560 11024 423 419 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14559 423 1284 286 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14558 285 425 423 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14557 11024 1284 425 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14556 286 3277 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14555 11024 726 285 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14554 419 423 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14553 11024 3276 3277 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14552 3276 7042 3130 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14551 3129 3284 3276 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14550 11024 7042 3284 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14549 3130 10995 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14548 11024 8297 3129 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14547 3277 3276 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14546 1537 2741 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14545 1537 6243 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14544 11024 7042 1537 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14543 11024 1881 1537 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14542 6918 10604 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14541 7031 8091 6918 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14540 11024 8930 7031 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14539 4036 3370 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14538 4036 3070 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14537 11024 4029 4036 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14536 1929 2435 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14535 2415 2434 1929 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14534 11024 4325 2415 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14533 9526 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14532 9526 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14531 11024 10031 9526 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14530 11024 8642 9526 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14529 11024 5728 5520 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14528 5520 5727 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14527 11024 10024 5520 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14526 5519 5520 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14525 11024 7459 7456 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14524 7456 7455 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14523 11024 7672 7456 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14522 8095 7456 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14521 11024 6232 6231 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14520 6231 6251 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14519 11024 6230 6231 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14518 8644 6231 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14517 11024 891 892 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14516 891 1248 786 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14515 785 893 891 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14514 11024 1248 893 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14513 786 4910 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14512 11024 902 785 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14511 892 891 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14510 11024 4913 4910 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14509 4913 5736 4912 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14508 4911 4914 4913 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14507 11024 5736 4914 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14506 4912 6401 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14505 11024 10257 4911 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14504 4910 4913 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14503 11024 9514 9503 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14502 11024 10774 9504 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14501 9503 9504 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14500 11024 7721 5794 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14499 5794 6277 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14498 5794 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14497 11024 8122 5794 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14496 6206 5794 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14495 10696 10693 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14494 10695 10694 10696 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14493 11024 10706 10695 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14492 5500 8122 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14491 5500 8885 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14490 11024 7484 5500 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14489 11024 7655 5500 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14488 5769 7045 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14487 11024 6142 5769 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14486 5766 5769 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14485 4321 4323 4244 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14484 11024 6213 4244 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14483 4244 5539 4321 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14482 4322 4321 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14481 11024 8082 7631 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14480 11024 10915 7435 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14479 7631 7435 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14478 9470 9971 9469 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14477 9469 10702 9713 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14476 9713 10694 9470 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14475 9470 10701 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14474 11024 10686 9470 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14473 9710 9713 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14472 7409 7414 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14471 11024 9305 7409 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14470 7408 7409 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14469 4340 4347 4341 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14468 4341 4348 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14467 11024 6503 4340 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14466 4450 4340 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14465 5006 5601 5005 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14464 5003 5008 5006 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14463 5004 5002 5003 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14462 11024 5009 5004 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14461 5024 5005 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14460 1459 7701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14459 11024 1456 1459 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14458 2434 1459 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14457 1406 7701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14456 11024 1403 1406 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14455 2004 1406 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14454 7571 7748 7747 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14453 11024 10027 7748 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14452 7572 8709 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14451 7747 10027 7572 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14450 11024 8708 7571 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14449 11024 10705 9709 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14448 9709 10378 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14447 9709 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14446 11024 11072 9709 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14445 9702 9709 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14444 3055 4014 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14443 3056 10018 3055 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14442 3054 6243 3056 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14441 11024 3714 3054 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14440 3064 3056 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14439 11024 8999 9005 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14438 9002 8995 8803 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14437 8803 8999 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14436 8803 9005 9002 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14435 11024 8998 8803 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14434 8998 8995 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14433 3950 6221 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14432 11024 6220 3950 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14431 5771 3950 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14430 3010 3008 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14429 3011 3009 3010 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14428 11024 6132 3011 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14427 748 10256 749 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14426 749 2472 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14425 11024 8713 748 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14424 752 748 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14423 3778 10596 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14422 3956 10595 3778 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14421 11024 10995 3956 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14420 10106 10269 10105 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14419 10105 10256 10243 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14418 10243 10258 10106 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14417 10106 10896 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14416 11024 10913 10106 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14415 10239 10243 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14414 11024 2133 2134 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14413 2134 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14412 11024 5918 2134 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14411 5736 2134 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14410 2401 3193 2402 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14409 2402 3626 2401 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14408 11024 3632 2402 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14407 5638 6803 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14406 5753 7437 5638 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14405 11024 8937 5753 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14404 7608 7690 7560 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14403 7560 7606 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14402 11024 9275 7608 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14401 7605 7608 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14400 11024 7711 2800 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14399 2800 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14398 2800 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14397 11024 7478 2800 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14396 2801 2800 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14395 11018 10366 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14394 10594 9509 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14393 11024 8746 6897 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14392 6897 8059 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14391 6897 8453 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14390 11024 9433 6897 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14389 6896 6897 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14388 11024 9426 7845 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14387 7845 9433 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14386 11024 9716 7845 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14385 7840 7845 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14384 275 1495 276 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14383 276 1494 346 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14382 346 348 276 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14381 275 338 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14380 11024 1489 275 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14379 276 341 275 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14378 2418 346 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14377 11024 3322 3039 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14376 3039 3311 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14375 3039 3306 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14374 11024 5771 3039 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14373 3285 3039 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14372 5691 6119 5633 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14371 5633 5698 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14370 11024 5703 5691 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14369 6195 5691 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14368 182 183 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14367 178 184 177 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14366 11024 723 178 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14365 184 185 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14364 11024 2446 185 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14363 11024 397 183 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14362 180 184 182 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14361 181 185 180 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14360 11024 179 181 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14359 179 180 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14358 177 185 179 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14357 11024 177 723 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14356 723 177 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14355 6159 6264 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14354 6157 6265 6260 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14353 11024 6261 6157 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14352 6265 6266 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14351 11024 8048 6266 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14350 11024 6538 6264 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14349 6263 6265 6159 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14348 6158 6266 6263 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14347 11024 6262 6158 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14346 6262 6263 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14345 6260 6266 6262 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14344 11024 6260 6261 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14343 6261 6260 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14342 10241 10595 10104 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14341 10104 10596 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14340 11024 10257 10241 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14339 10585 10241 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14338 1933 5557 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14337 2073 2452 1933 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14336 11024 5766 2073 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14335 3922 3941 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14334 11024 3938 3922 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14333 805 1003 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14332 803 1002 992 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14331 11024 1490 803 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14330 1002 1004 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14329 11024 2446 1004 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14328 11024 1265 1003 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14327 997 1002 805 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14326 804 1004 997 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14325 11024 998 804 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14324 998 997 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14323 992 1004 998 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14322 11024 992 1490 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14321 1490 992 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14320 10037 10595 9937 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14319 9937 10596 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14318 11024 11018 10037 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14317 10032 10037 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14316 2081 7027 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14315 11024 2035 2081 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14314 10269 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14313 11024 9560 10269 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14312 5558 5556 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14311 10081 5557 5558 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14310 11024 5776 10081 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14309 8939 9347 8790 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14308 8790 10908 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14307 11024 8938 8939 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14306 8937 8939 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14305 3668 3928 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14304 11024 4410 3668 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14303 10626 10628 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14302 10622 10629 10623 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14301 11024 10909 10622 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14300 10629 10630 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14299 11024 10914 10630 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14298 11024 10995 10628 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14297 10627 10629 10626 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14296 10625 10630 10627 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14295 11024 10624 10625 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14294 10624 10627 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14293 10623 10630 10624 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14292 11024 10623 10909 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14291 10909 10623 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14290 122 124 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14289 118 125 119 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14288 11024 8839 118 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14287 125 126 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14286 11024 2673 126 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14285 11024 4885 124 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14284 123 125 122 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14283 120 126 123 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14282 11024 121 120 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14281 121 123 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14280 119 126 121 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14279 11024 119 8839 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14278 8839 119 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14277 11024 4961 4969 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14276 4961 10915 4963 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14275 4962 4964 4961 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14274 11024 10915 4964 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14273 4963 5191 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14272 11024 6465 4962 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14271 4969 4961 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14270 9471 9760 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14269 9724 10694 9471 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14268 11024 10702 9724 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14267 8771 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14266 8770 10710 8771 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14265 11024 10686 8770 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14264 5073 6586 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14263 5297 5292 5073 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14262 11024 5293 5297 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14261 725 1495 727 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14260 727 1494 728 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14259 728 726 727 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14258 725 723 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14257 11024 1489 725 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14256 727 724 725 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14255 3009 728 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14254 10002 10880 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14253 10002 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14252 11024 10027 10002 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14251 3037 4070 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14250 3037 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14249 11024 6275 3037 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14248 9961 10058 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14247 9959 10060 10053 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14246 11024 10054 9959 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14245 10060 10057 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14244 11024 11051 10057 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14243 11024 10059 10058 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14242 10056 10060 9961 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14241 9960 10057 10056 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14240 11024 10055 9960 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14239 10055 10056 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14238 10053 10057 10055 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14237 11024 10053 10054 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14236 10054 10053 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14235 9269 9271 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14234 9265 9272 9266 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14233 11024 10213 9265 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14232 9272 9273 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14231 11024 10914 9273 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_14230 11024 10177 9271 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14229 9270 9272 9269 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14228 9268 9273 9270 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14227 11024 9267 9268 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14226 9267 9270 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14225 9266 9273 9267 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_14224 11024 9266 10213 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14223 10213 9266 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14222 11024 3023 3272 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14221 3023 10959 3025 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14220 3024 3026 3023 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14219 11024 10959 3026 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14218 3025 3263 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14217 11024 8305 3024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14216 3272 3023 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14215 11024 4269 4496 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14214 4269 10959 4241 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14213 4239 4242 4269 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14212 11024 10959 4242 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14211 4241 4240 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14210 11024 7601 4239 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14209 4496 4269 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14208 11024 4514 4892 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14207 4514 10959 4379 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14206 4378 4518 4514 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14205 11024 10959 4518 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14204 4379 4524 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14203 11024 7418 4378 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14202 4892 4514 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14201 11024 1819 1816 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14200 1819 10959 1817 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14199 1818 1820 1819 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14198 11024 10959 1820 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14197 1817 2003 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14196 11024 7425 1818 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14195 1816 1819 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14194 11024 2066 2062 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14193 2066 10959 1932 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14192 1931 2070 2066 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14191 11024 10959 2070 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14190 1932 2073 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14189 11024 7450 1931 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14188 2062 2066 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14187 11024 2023 2019 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14186 2023 10959 1927 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14185 1926 2028 2023 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14184 11024 10959 2028 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14183 1927 2024 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14182 11024 7611 1926 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14181 2019 2023 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14180 6998 7655 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14179 6998 6992 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14178 11024 8122 6998 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14177 4524 3832 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14176 11024 1409 4524 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14175 1042 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14174 11024 7514 1042 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14173 2661 4617 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14172 11024 4553 2661 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14171 3632 2661 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14170 2627 3817 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14169 11024 4915 2627 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14168 2965 2627 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14167 5176 5181 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14166 11024 6246 5176 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14165 5175 5176 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14164 4916 4959 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14163 4916 5521 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14162 11024 5522 4916 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14161 11024 4954 4916 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14160 3673 3945 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14159 3677 3925 3673 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14158 11024 9987 3677 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14157 11024 2707 2709 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14156 2707 10959 2527 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14155 2526 2718 2707 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14154 11024 10959 2718 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14153 2527 2717 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14152 11024 7466 2526 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14151 2709 2707 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14150 11024 2080 2074 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14149 2080 10959 1935 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14148 1934 2083 2080 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14147 11024 10959 2083 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14146 1935 2081 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14145 11024 7474 1934 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14144 2074 2080 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14143 11024 2699 3019 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14142 2699 10959 2525 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14141 2524 2700 2699 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14140 11024 10959 2700 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14139 2525 3012 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14138 11024 7037 2524 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_14137 3019 2699 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14136 6483 7478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14135 6483 10029 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14134 11024 6275 6483 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14133 11024 8409 6483 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14132 4376 10604 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14131 5665 8091 4376 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14130 11024 8642 5665 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14129 1930 2434 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14128 2035 2435 1930 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14127 11024 10888 2035 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14126 4042 6173 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14125 11024 4183 4042 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14124 2370 3714 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14123 2476 2572 2370 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14122 2369 2728 2476 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14121 11024 4014 2369 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14120 4453 2476 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14119 4981 7514 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14118 4981 5583 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14117 11024 6275 4981 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14116 1542 1055 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14115 1542 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14114 11024 6275 1542 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14113 2114 3703 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14112 2114 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14111 11024 8922 2114 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14110 11024 10002 10001 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14109 10001 10003 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14108 11024 10004 10001 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14107 10000 10001 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14106 11024 5153 4289 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14105 4289 5718 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14104 11024 5131 4289 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14103 4288 4289 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14102 11024 5159 4302 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14101 4302 6127 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14100 11024 5131 4302 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14099 4301 4302 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14098 2466 1871 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14097 2466 1870 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14096 11024 2109 2466 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14095 11024 2114 2466 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14094 3337 3709 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14093 3337 3338 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14092 11024 3331 3337 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14091 11024 3994 3337 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14090 9334 9333 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14089 9332 9609 9334 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14088 11024 9603 9332 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14087 1941 4014 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14086 2153 2578 1941 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14085 1940 2741 2153 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14084 11024 3714 1940 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14083 3063 2153 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14082 3739 5719 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14081 3739 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14080 11024 9309 3739 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14079 11024 5918 3739 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14078 7204 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14077 7204 8746 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14076 11024 8453 7204 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14075 11024 9433 7204 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14074 11024 3084 2545 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14073 2545 3082 2787 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14072 2788 2787 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14071 5936 6905 5648 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14070 5648 6286 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14069 11024 5933 5936 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14068 5934 5936 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14067 8781 8864 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14066 8878 8865 8781 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14065 11024 8866 8878 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14064 9428 9980 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14063 9427 9976 9428 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14062 11024 9426 9427 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14061 3792 4014 4006 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14060 3791 4347 3792 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14059 11024 4348 3791 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14058 4005 4006 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14057 7565 8318 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14056 8084 8316 7565 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14055 11024 8970 8084 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14054 5718 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14053 5718 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14052 11024 5719 5718 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14051 11024 8869 5718 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14050 11024 10078 10077 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14049 10077 10701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14048 11024 10700 10077 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14047 11066 10077 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14046 5045 5093 5092 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14045 5046 10604 5045 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14044 5044 10892 5046 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14043 11024 10888 5044 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_14042 5091 5092 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14041 5677 6762 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14040 11024 6108 5677 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14039 5672 5677 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14038 2112 2121 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14037 11024 4012 2112 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14036 2109 2112 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14035 3359 3379 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14034 11024 6275 3359 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14033 3723 3359 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14032 3048 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14031 11024 6277 3048 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14030 3969 3048 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14029 1399 7701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14028 11024 1396 1399 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14027 2417 1399 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14026 9301 9347 9302 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14025 9302 9955 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14024 11024 9559 9301 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14023 9300 9301 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14022 5551 10608 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14021 5550 10606 5551 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14020 11024 8305 5550 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14019 7413 7690 7412 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14018 7412 7411 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14017 11024 8000 7413 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14016 7410 7413 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14015 7454 7690 7453 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14014 7453 7452 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14013 11024 10239 7454 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14012 7451 7454 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_14011 8159 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14010 11024 11072 8159 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14009 8063 8159 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14008 11024 472 218 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14007 218 1545 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14006 11024 4673 218 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_14005 217 218 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14004 11024 5131 5053 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14003 5053 5523 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14002 5684 5128 5053 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14001 5052 5124 5684 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_14000 5053 5681 5052 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13999 8109 8212 8032 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13998 8032 8113 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13997 11024 8112 8109 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13996 8340 8109 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13995 11024 3355 3080 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13994 3080 3079 3081 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13993 11024 6905 6907 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13992 6907 7217 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13991 6907 7212 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13990 11024 6906 6907 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13989 6904 6907 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13988 9923 10614 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13987 9998 10615 9923 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13986 11024 10312 9998 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13985 3098 3100 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13984 3093 3099 3094 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13983 11024 3092 3093 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13982 3099 3101 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13981 11024 5262 3101 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13980 11024 4370 3100 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13979 3096 3099 3098 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13978 3097 3101 3096 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13977 11024 3095 3097 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13976 3095 3096 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13975 3094 3101 3095 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13974 11024 3094 3092 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13973 3092 3094 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13972 6932 7127 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13971 6930 7126 7119 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13970 11024 7117 6930 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13969 7126 7128 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13968 11024 8048 7128 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13967 11024 7518 7127 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13966 7124 7126 6932 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13965 6931 7128 7124 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13964 11024 7122 6931 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13963 7122 7124 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13962 7119 7128 7122 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13961 11024 7119 7117 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13960 7117 7119 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13959 5928 6286 5646 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13958 5646 7204 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13957 11024 5927 5928 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13956 5926 5928 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13955 11024 8124 2786 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13954 2786 3092 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13953 2786 4066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13952 11024 4070 2786 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13951 3379 2786 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13950 11024 2590 2494 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13949 2494 2589 2782 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13948 11024 6276 1313 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13947 1313 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13946 1313 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13945 11024 5911 1313 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13944 2212 1313 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13943 11024 9309 5013 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13942 5013 5012 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13941 5013 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13940 11024 8643 5013 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13939 5292 5013 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13938 4309 4318 4308 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13937 4308 4925 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13936 11024 4926 4309 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13935 4307 4309 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13934 4491 5496 4375 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13933 4375 4489 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13932 11024 6206 4491 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13931 4488 4491 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13930 205 206 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13929 201 207 200 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13928 11024 726 201 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13927 207 208 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13926 11024 5262 208 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13925 11024 419 206 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13924 203 207 205 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13923 204 208 203 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13922 11024 202 204 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13921 202 203 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13920 200 208 202 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13919 11024 200 726 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13918 726 200 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13917 1287 759 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13916 1287 752 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13915 11024 1041 1287 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13914 2090 2094 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13913 2090 2456 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13912 11024 5727 2090 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13911 2098 2094 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13910 2098 2093 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13909 11024 5727 2098 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13908 4370 4368 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13907 11024 4369 4370 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13906 5553 5552 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13905 5777 10606 5553 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13904 11024 8918 5777 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13903 5490 6978 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13902 11024 1991 5490 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13901 4628 4327 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13900 11024 8713 4628 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13899 6814 7437 6813 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13898 6813 9610 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13897 11024 9346 6814 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13896 6811 6814 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13895 6836 6838 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13894 6832 6839 6833 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13893 11024 7085 6832 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13892 6839 6840 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13891 11024 8048 6840 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13890 11024 7089 6838 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13889 6837 6839 6836 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13888 6834 6840 6837 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13887 11024 6835 6834 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13886 6835 6837 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13885 6833 6840 6835 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13884 11024 6833 7085 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13883 7085 6833 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13882 1910 2016 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13881 1908 2017 2009 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13880 11024 7611 1908 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13879 2017 2018 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13878 11024 2673 2018 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13877 11024 2019 2016 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13876 2014 2017 1910 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13875 1909 2018 2014 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13874 11024 2011 1909 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13873 2011 2014 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13872 2009 2018 2011 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13871 11024 2009 7611 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13870 7611 2009 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13869 6202 6406 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13868 6196 6324 6403 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13867 11024 6992 6196 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13866 6324 6407 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13865 11024 10914 6407 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13864 11024 6404 6406 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13863 6323 6324 6202 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13862 6199 6407 6323 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13861 11024 6320 6199 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13860 6320 6323 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13859 6403 6407 6320 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13858 11024 6403 6992 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13857 6992 6403 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13856 10569 10583 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13855 10566 10564 10569 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13854 11024 10565 10566 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13853 7446 7444 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13852 7445 7463 7446 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13851 11024 7467 7445 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13850 11061 10707 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13849 11024 10704 11061 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13848 10692 10695 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13847 11024 10691 10692 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13846 10074 9427 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13845 11024 9424 10074 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13844 9044 10687 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13843 11024 9033 9044 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13842 5288 5307 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13841 11024 5897 5288 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13840 2999 5726 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13839 3646 2997 2999 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13838 11024 3236 3646 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13837 4267 4498 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13836 4259 4497 4494 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13835 11024 7601 4259 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13834 4497 4499 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13833 11024 5083 4499 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13832 11024 4496 4498 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13831 4407 4497 4267 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13830 4264 4499 4407 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13829 11024 4405 4264 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13828 4405 4407 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13827 4494 4499 4405 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13826 11024 4494 7601 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13825 7601 4494 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13824 9570 9603 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13823 11024 10018 9570 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13822 10014 9570 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13821 9572 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13820 9572 8661 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13819 11024 10031 9572 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13818 11024 8699 9572 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13817 9409 10687 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13816 11024 9395 9409 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13815 7532 8762 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13814 7532 7531 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13813 11024 8765 7532 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13812 2480 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13811 2480 9560 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13810 11024 7721 2480 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13809 9747 10083 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13808 11024 11072 9747 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13807 11024 8692 8989 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13806 8692 9350 8695 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13805 8693 8696 8692 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13804 11024 9350 8696 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13803 8695 8694 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13802 11024 8691 8693 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13801 8989 8692 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13800 11024 8984 8999 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13799 8984 9376 8802 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13798 8801 8993 8984 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13797 11024 9376 8993 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13796 8802 8989 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13795 11024 8985 8801 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13794 8999 8984 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13793 5034 5033 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13792 11024 5606 5034 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13791 11024 8318 6812 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13790 6810 6812 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13789 11024 10018 6810 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13788 6809 6810 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13787 11024 6810 6809 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13786 6807 7041 6808 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13785 11024 10772 6808 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13784 6808 7042 6807 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13783 6806 6807 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13782 3189 4274 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13781 11024 4926 3189 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13780 3188 3189 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13779 4294 4555 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13778 11024 4410 4294 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13777 4932 4294 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13776 5159 10680 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13775 5159 5728 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13774 11024 5727 5159 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13773 11024 148 145 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13772 148 1248 146 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13771 147 149 148 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13770 11024 1248 149 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13769 146 4905 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13768 11024 341 147 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13767 145 148 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13766 9541 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13765 9541 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13764 11024 9560 9541 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13763 11024 10825 9541 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13762 1326 2004 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13761 1401 2006 1326 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13760 11024 10888 1401 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13759 2578 7478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13758 2578 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13757 11024 5918 2578 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13756 8055 10710 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13755 8152 10083 8055 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13754 11024 11072 8152 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13753 7212 8453 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13752 7212 8059 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13751 11024 8746 7212 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13750 11024 9107 7212 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13749 11024 8953 8985 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13748 8953 9350 8795 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13747 8794 8960 8953 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13746 11024 9350 8960 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13745 8795 9335 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13744 11024 8954 8794 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13743 8985 8953 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13742 5307 5593 5070 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13741 5070 5271 5307 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13740 11024 5878 5070 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13739 2485 2741 2486 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13738 2486 4014 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13737 11024 2487 2485 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13736 3068 2485 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13735 3322 4070 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13734 3322 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13733 11024 5898 3322 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13732 2746 8124 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13731 2746 5898 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13730 11024 7514 2746 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13729 10559 10555 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13728 10559 10551 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13727 11024 10546 10559 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13726 11024 10547 10559 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13725 11024 4908 4905 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13724 4908 5736 4907 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13723 4906 4909 4908 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13722 11024 5736 4909 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13721 4907 6106 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13720 11024 10231 4906 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13719 4905 4908 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13718 9306 8921 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13717 9306 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13716 11024 9560 9306 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13715 11024 10854 9306 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13714 4991 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13713 4991 5012 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13712 11024 10031 4991 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13711 11024 8643 4991 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13710 9532 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13709 9532 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13708 11024 9309 9532 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13707 11024 8885 9532 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13706 11024 4981 4647 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13705 4647 7068 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13704 11024 4658 4647 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13703 4983 4647 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13702 2396 3844 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13701 2398 2393 2395 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13700 2395 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13699 11024 2394 2399 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13698 2399 2401 2397 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13697 2397 2396 2398 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13696 2398 3844 2400 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13695 2400 3626 2399 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13694 11024 4929 2394 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13693 3606 2398 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13692 11024 5684 5517 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13691 5693 5518 5516 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13690 5516 5684 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13689 5516 5517 5693 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13688 11024 5515 5516 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13687 5515 5518 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13686 11024 333 329 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13685 333 1248 274 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13684 273 337 333 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13683 11024 1248 337 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13682 274 5510 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13681 11024 692 273 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13680 329 333 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13679 6296 6469 9362 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13678 11024 9987 6469 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13677 6297 6468 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13676 9362 9987 6297 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13675 11024 6465 6296 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13674 7010 7007 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13673 11024 7655 7010 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13672 7006 7010 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13671 8104 8388 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13670 11024 8970 8104 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13669 8030 8104 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13668 8083 8638 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13667 11024 8084 8083 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13666 8012 8083 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13665 10579 10577 10580 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13664 10580 10578 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13663 11024 10800 10579 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13662 10576 10579 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13661 6980 7437 6914 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13660 6914 8893 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13659 11024 7012 6980 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13658 6978 6980 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13657 11024 2630 308 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13656 1796 2385 270 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13655 270 2630 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13654 270 308 1796 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13653 11024 304 270 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13652 304 2385 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13651 11024 8918 5503 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13650 11024 10915 5505 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13649 5503 5505 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13648 858 3152 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13647 11024 4255 858 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13646 3833 858 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13645 3733 3735 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13644 11024 6275 3733 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13643 4030 3733 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13642 2488 2782 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13641 11024 3065 2488 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13640 2492 2488 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13639 11024 8839 5162 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13638 11024 10915 5163 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13637 5162 5163 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13636 8251 8261 8161 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13635 11024 8624 8161 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13634 8161 8613 8251 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13633 8252 8251 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13632 8780 8862 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13631 9293 9295 8780 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13630 11024 9987 9293 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13629 11024 7484 6189 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13628 6189 8122 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13627 11024 7655 6189 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13626 6105 6189 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13625 9052 10698 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13624 11024 10708 9052 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13623 9051 9052 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13622 11024 11076 8156 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13621 8156 10710 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13620 11024 10700 8156 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13619 8059 8156 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13618 7541 10399 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13617 11024 9716 7541 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13616 9424 7541 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13615 11024 5911 1298 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13614 1298 7514 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13613 11024 8124 1298 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13612 1520 1298 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13611 1938 2104 7673 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13610 1937 2105 1938 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13609 11024 2102 1937 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13608 8683 8682 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13607 8680 8690 8683 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13606 8681 8684 8680 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13605 11024 10606 8681 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13604 8679 8680 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13603 7131 7786 6933 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13602 6933 8053 7131 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13601 11024 7129 6933 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13600 10680 10323 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13599 10995 10908 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13598 11024 9020 5249 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13597 5249 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13596 11024 7721 5249 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13595 10606 5249 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13594 11024 4048 3799 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13593 3799 4047 5321 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13592 3727 3722 3724 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13591 3724 3723 3725 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13590 3725 5901 3727 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13589 3727 7523 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13588 11024 6574 3727 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13587 3721 3725 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13586 11024 2099 1551 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13585 1551 1552 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13584 1551 2121 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13583 11024 2480 1551 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13582 1545 1551 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13581 1215 1219 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13580 1212 1218 1213 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13579 11024 1403 1212 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13578 1218 1220 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13577 11024 2673 1220 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13576 11024 1235 1219 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13575 1216 1218 1215 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13574 1217 1220 1216 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13573 11024 1214 1217 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13572 1214 1216 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13571 1213 1220 1214 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13570 11024 1213 1403 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13569 1403 1213 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13568 10041 10606 9941 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13567 9941 10608 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13566 11024 10963 10041 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13565 10043 10041 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13564 9688 10054 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13563 288 466 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13562 438 437 288 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13561 287 449 438 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13560 11024 451 287 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13559 1489 438 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13558 5705 5704 5635 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13557 5635 6201 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13556 11024 5702 5705 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13555 5703 5705 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13554 4332 4676 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13553 4330 4675 4672 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13552 11024 4673 4330 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13551 4675 4677 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13550 11024 5262 4677 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13549 11024 6525 4676 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13548 4438 4675 4332 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13547 4331 4677 4438 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13546 11024 4436 4331 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13545 4436 4438 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13544 4672 4677 4436 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13543 11024 4672 4673 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13542 4673 4672 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13541 7455 8834 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13540 11024 7652 7455 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13539 4318 4323 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13538 11024 5539 4318 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13537 163 165 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13536 159 166 160 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13535 11024 951 159 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13534 166 167 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13533 11024 2673 167 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13532 11024 934 165 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13531 164 166 163 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13530 161 167 164 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13529 11024 162 161 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13528 162 164 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13527 160 167 162 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13526 11024 160 951 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13525 951 160 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13524 1323 1385 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13523 1321 1384 1376 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13522 11024 8617 1321 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13521 1384 1386 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13520 11024 5083 1386 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13519 11024 8312 1385 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13518 1382 1384 1323 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13517 1322 1386 1382 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13516 11024 1380 1322 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13515 1380 1382 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13514 1376 1386 1380 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13513 11024 1376 8617 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13512 8617 1376 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13511 11024 7733 7727 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13510 7733 8708 7552 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13509 7551 7737 7733 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13508 11024 8708 7737 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13507 7552 8297 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13506 11024 8408 7551 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13505 7727 7733 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13504 3012 6440 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13503 11024 3011 3012 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13502 3718 4335 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13501 11024 5293 3718 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13500 4306 5165 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13499 11024 4305 4306 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13498 9970 10068 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13497 9968 10064 10063 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13496 11024 10350 9968 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13495 10064 10065 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13494 11024 11051 10065 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13493 11024 10348 10068 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13492 10067 10064 9970 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13491 9969 10065 10067 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13490 11024 10066 9969 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13489 10066 10067 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13488 10063 10065 10066 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13487 11024 10063 10350 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13486 10350 10063 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13485 1527 4981 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13484 11024 1881 1527 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13483 1868 1527 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13482 11024 5870 5866 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13481 5870 10687 5629 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13480 5630 5872 5870 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13479 11024 10687 5872 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13478 5629 6571 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13477 11024 5863 5630 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13476 5866 5870 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13475 7004 8930 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13474 7004 7007 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13473 11024 7655 7004 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13472 6585 7852 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13471 6585 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13470 11024 10704 6585 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13469 8188 8477 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13468 8474 9974 8188 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13467 8187 9100 8474 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13466 11024 8475 8187 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13465 8472 8474 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13464 5770 8316 5549 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13463 5549 5561 5770 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13462 11024 8318 5549 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13461 5181 4658 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13460 5181 4981 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13459 11024 7068 5181 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13458 7072 7069 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13457 11024 7068 7072 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13456 9347 7072 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13455 9437 9484 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13454 9435 9483 9475 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13453 11024 9922 9435 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13452 9483 9485 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13451 11024 10914 9485 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13450 11024 9916 9484 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13449 9482 9483 9437 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13448 9436 9485 9482 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13447 11024 9479 9436 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13446 9479 9482 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13445 9475 9485 9479 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13444 11024 9475 9922 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13443 9922 9475 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13442 9589 9613 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13441 11024 10018 9589 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13440 10249 9589 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13439 6943 6942 6909 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13438 6909 8831 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13437 11024 10774 6943 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13436 6941 6943 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13435 6908 9433 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13434 11024 9716 6908 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13433 4996 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13432 4996 5253 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13431 11024 10031 4996 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13430 11024 8126 4996 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13429 5580 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13428 5580 5579 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13427 11024 8661 5580 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13426 11024 8643 5580 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13425 11024 2473 502 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13424 501 502 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13423 11024 3413 501 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13422 499 501 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13421 11024 501 499 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13420 3136 4014 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13419 3352 6221 3136 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13418 3135 10018 3352 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13417 11024 3714 3135 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13416 3349 3352 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13415 8176 8318 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13414 8650 8316 8176 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13413 11024 9335 8650 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13412 10207 10206 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13411 11024 10212 10207 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13410 10570 10207 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13409 5522 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13408 5522 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13407 11024 6277 5522 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13406 11024 9287 5522 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13405 11024 2993 2996 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13404 2993 4291 2992 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13403 2991 2994 2993 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13402 11024 4291 2994 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13401 2992 4617 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13400 11024 4553 2991 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13399 2996 2993 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13398 8079 8080 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13397 11024 10018 8079 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13396 8009 8079 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13395 3983 4666 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13394 3983 6221 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13393 11024 4665 3983 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13392 11024 7069 3983 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13391 11024 6279 6273 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13390 6279 10687 6170 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13389 6168 6169 6279 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13388 11024 10687 6169 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13387 6170 9074 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13386 11024 6493 6168 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13385 6273 6279 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13384 7519 9046 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13383 7518 7525 7519 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13382 11024 7517 7518 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13381 11024 3413 493 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13380 491 493 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13379 11024 2473 491 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13378 494 491 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13377 11024 491 494 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13376 4249 4654 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13375 4329 4653 4249 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13374 4248 5911 4329 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13373 11024 7678 4248 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13372 10614 4329 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13371 1300 7041 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13370 1300 5809 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13369 11024 1552 1300 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13368 11024 2099 1300 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13367 11024 9655 10073 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13366 9655 10684 9450 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13365 9449 9658 9655 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13364 11024 10684 9658 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13363 9450 10231 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13362 11024 10289 9449 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13361 10073 9655 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13360 5772 5771 5639 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13359 5639 6455 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13358 11024 5770 5772 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13357 5774 5772 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13356 11024 3306 3302 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13355 3302 3322 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13354 3302 5771 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13353 11024 4012 3302 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13352 7437 3302 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13351 11024 6765 6767 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13350 6767 6766 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13349 11024 7655 6767 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13348 6764 6767 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13347 6286 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13346 6286 7478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13345 11024 7514 6286 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13344 11024 5607 6286 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13343 5910 6176 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13342 11024 5906 5910 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13341 5908 5910 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13340 6219 7430 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13339 11024 6820 6219 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13338 6140 6219 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13337 788 1495 787 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13336 787 1494 911 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13335 911 1423 787 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13334 788 901 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13333 11024 1489 788 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13332 787 902 788 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13331 2006 911 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13330 2988 3860 2987 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13329 2987 2986 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13328 11024 4553 2988 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13327 2985 2988 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13326 2521 2691 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13325 3007 2692 2521 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13324 11024 2688 3007 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13323 11024 4943 4577 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13322 4950 4940 4385 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13321 4385 4943 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13320 4385 4577 4950 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13319 11024 4578 4385 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13318 4578 4940 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13317 11024 8848 8627 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13316 11024 10197 8628 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13315 8627 8628 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13314 7416 7415 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13313 11024 7655 7416 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13312 7421 7416 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13311 11024 9560 1887 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13310 1887 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13309 1887 6275 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13308 11024 7478 1887 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13307 1886 1887 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13306 11024 7711 4678 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13305 4678 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13304 4678 8921 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13303 11024 5293 4678 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13302 4679 4678 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13301 11024 5600 4650 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13300 4650 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13299 11024 5898 4650 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13298 5552 4650 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13297 3767 4080 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13296 3765 4079 4074 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13295 11024 4070 3765 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13294 4079 4081 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13293 11024 5262 4081 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13292 11024 4374 4080 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13291 4078 4079 3767 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13290 3766 4081 4078 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13289 11024 4073 3766 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13288 4073 4078 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13287 4074 4081 4073 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13286 11024 4074 4070 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13285 4070 4074 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13284 11024 10915 661 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13283 660 661 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13282 11024 4254 660 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13281 2609 660 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13280 11024 660 2609 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13279 9328 10595 9327 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13278 9327 10596 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13277 11024 10024 9328 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13276 9329 9328 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13275 11024 6171 4053 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13274 4053 4054 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13273 4053 4057 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13272 11024 4058 4053 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13271 4363 4053 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13270 3713 3712 4000 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13269 3711 3982 3713 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13268 11024 3710 3711 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13267 3788 4005 4344 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13266 3787 4000 3788 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13265 11024 4451 3787 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13264 11024 5017 4366 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13263 4365 4366 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13262 11024 4364 4365 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13261 4368 4365 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13260 11024 4365 4368 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13259 11024 3739 3388 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13258 3388 3738 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13257 3388 3396 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13256 11024 3151 3388 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13255 3382 3388 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13254 9455 9677 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13253 9453 9676 9669 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13252 11024 9667 9453 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13251 9676 9679 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13250 11024 11051 9679 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13249 11024 9682 9677 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13248 9674 9676 9455 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13247 9454 9679 9674 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13246 11024 9673 9454 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13245 9673 9674 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13244 9669 9679 9673 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13243 11024 9669 9667 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13242 9667 9669 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13241 6805 8644 6804 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13240 6804 6803 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13239 11024 7036 6805 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13238 7459 6805 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13237 11024 3337 2531 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13236 2532 3046 2576 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13235 2533 2752 2532 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13234 2531 2575 2533 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13233 3134 3698 3133 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13232 3338 10028 3134 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13231 3134 4654 3338 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13230 3133 5911 3134 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13229 3133 3969 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13228 11024 5918 3133 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13227 9348 9347 9349 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13226 9349 10323 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13225 11024 9613 9348 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13224 9346 9348 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13223 1919 2223 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13222 1917 2222 2217 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13221 11024 2473 1917 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13220 2222 2224 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13219 11024 5262 2224 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13218 11024 4063 2223 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13217 2221 2222 1919 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13216 1918 2224 2221 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13215 11024 2216 1918 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13214 2216 2221 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13213 2217 2224 2216 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13212 11024 2217 2473 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13211 2473 2217 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13210 2445 2444 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13209 2439 2448 2440 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13208 11024 7466 2439 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13207 2448 2447 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13206 11024 2446 2447 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13205 11024 2709 2444 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13204 2442 2448 2445 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13203 2443 2447 2442 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13202 11024 2441 2443 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13201 2441 2442 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13200 2440 2447 2441 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13199 11024 2440 7466 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13198 7466 2440 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13197 3105 3167 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13196 3103 3168 3160 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13195 11024 8642 3103 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13194 3168 3169 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13193 11024 5083 3169 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13192 11024 6370 3167 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13191 3166 3168 3105 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13190 3104 3169 3166 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13189 11024 3164 3104 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13188 3164 3166 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13187 3160 3169 3164 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13186 11024 3160 8642 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13185 8642 3160 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13184 1292 1556 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13183 1292 1061 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13182 11024 2099 1292 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13181 4658 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13180 4658 7711 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13179 11024 7721 4658 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13178 6284 6902 6181 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13177 6181 6286 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13176 11024 6285 6284 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13175 6180 6284 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13174 6214 10594 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13173 6214 5728 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13172 11024 5727 6214 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13171 1268 1504 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13170 11024 1489 1268 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13169 9467 10269 9466 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13168 9466 10256 9627 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13167 9627 10258 9467 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13166 9467 9938 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13165 11024 9939 9467 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13164 9624 9627 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13163 1556 7514 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13162 1556 5898 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13161 11024 7721 1556 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13160 4439 4679 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13159 11024 9002 4439 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13158 11024 4956 4958 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13157 4957 4958 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13156 11024 5177 4957 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13155 4955 4957 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13154 11024 4957 4955 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13153 7431 8869 7429 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13152 7430 9922 7431 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13151 7431 8635 7430 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13150 7429 8636 7431 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13149 7429 9313 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13148 11024 8633 7429 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13147 4891 4893 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13146 4886 4894 4887 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13145 11024 7418 4886 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13144 4894 4895 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13143 11024 5083 4895 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_13142 11024 4892 4893 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13141 4890 4894 4891 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13140 4889 4895 4890 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13139 11024 4888 4889 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13138 4888 4890 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13137 4887 4895 4888 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13136 11024 4887 7418 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13135 7418 4887 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13134 10008 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13133 10008 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13132 11024 10031 10008 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13131 11024 9313 10008 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13130 7675 7673 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13129 11024 7670 7675 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13128 7672 7675 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13127 7824 10700 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13126 7824 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13125 11024 9412 7824 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13124 3370 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13123 3370 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13122 11024 3379 3370 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13121 11024 4048 3139 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13120 3139 4047 3393 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13119 3391 3393 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13118 3032 2728 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13117 3032 3033 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13116 11024 7042 3032 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13115 9992 10564 9919 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13114 9919 10772 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13113 11024 9994 9992 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13112 10182 9992 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_13111 2977 3844 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13110 2979 2974 2976 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13109 2976 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13108 11024 2975 2981 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13107 2981 3179 2978 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13106 2978 2977 2979 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13105 2979 3844 2980 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13104 2980 3183 2981 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13103 11024 4929 2975 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13102 2973 2979 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13101 6854 6861 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13100 6857 10366 6853 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13099 6853 8709 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13098 11024 6852 6858 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13097 6858 7117 6855 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13096 6855 6854 6857 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13095 6857 6861 6856 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13094 6856 9605 6858 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_13093 11024 8709 6852 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_13092 6851 6857 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13091 11024 5511 5510 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13090 5511 5736 5513 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13089 5512 5514 5511 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13088 11024 5736 5514 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13087 5513 7422 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13086 11024 10312 5512 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13085 5510 5511 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13084 9559 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13083 9559 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13082 11024 9560 9559 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13081 11024 10880 9559 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13080 6210 6465 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13079 11024 9987 6210 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13078 5890 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13077 5890 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13076 11024 10029 5890 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13075 11024 7721 5890 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13074 6895 8052 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13073 6895 9057 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13072 11024 9433 6895 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13071 11024 9716 6895 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13070 6579 10704 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13069 6579 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13068 11024 6574 6579 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13067 11024 9747 6579 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13066 11024 5684 5689 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13065 6200 5681 5632 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13064 5632 5684 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13063 5632 5689 6200 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13062 11024 5685 5632 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13061 5685 5681 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13060 3886 5153 3756 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13059 11024 6213 3756 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13058 3756 5718 3886 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13057 3884 3886 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13056 11024 744 1025 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13055 744 1248 658 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13054 657 659 744 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13053 11024 1248 659 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13052 658 5544 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13051 11024 1496 657 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13050 1025 744 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13049 11024 5547 5544 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13048 5547 7042 5545 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13047 5546 5548 5547 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13046 11024 7042 5548 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13045 5545 10024 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13044 11024 8918 5546 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13043 5544 5547 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13042 11024 1246 1244 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13041 1246 1248 1249 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13040 1247 1250 1246 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13039 11024 1248 1250 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13038 1249 5707 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13037 11024 1245 1247 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13036 1244 1246 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13035 11024 5712 5707 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13034 5712 5736 5617 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13033 5616 5715 5712 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13032 11024 5736 5715 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13031 5617 6117 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13030 11024 10594 5616 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13029 5707 5712 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13028 5750 8021 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13027 11024 6131 5750 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13026 5746 5750 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13025 7442 7444 7443 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13024 7440 10604 7442 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13023 7441 10892 7440 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13022 11024 10888 7441 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13021 7439 7443 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13020 9458 9513 9509 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13019 11024 10774 9513 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_13018 9459 9514 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13017 9509 10774 9459 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13016 11024 9505 9458 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13015 2203 9560 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13014 2203 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13013 11024 5600 2203 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13012 11024 9308 2203 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_13011 5020 5286 5022 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13010 5021 5288 5020 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13009 5019 5018 5021 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13008 11024 5024 5019 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13007 5017 5022 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13006 3138 3377 3378 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13005 3137 3375 3138 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13004 11024 3721 3137 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_13003 4064 3378 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13002 10092 10614 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13001 10212 10615 10092 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_13000 11024 10257 10212 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12999 11024 2630 1211 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12998 1210 2967 1209 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12997 1209 2630 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12996 1209 1211 1210 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12995 11024 1208 1209 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12994 1208 2967 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12993 11024 1310 1311 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12992 9314 1311 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12991 11024 1311 9314 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12990 11024 1311 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12989 11024 1311 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12988 11024 1310 1070 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12987 8661 1070 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12986 11024 1070 8661 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12985 11024 1070 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12984 11024 1070 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12983 11024 767 766 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12982 1310 766 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12981 11024 766 1310 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12980 11024 766 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12979 11024 766 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12978 11024 9987 8625 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12977 8626 8625 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12976 11024 8623 8626 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12975 8624 8626 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12974 11024 8626 8624 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12973 1064 3413 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12972 11024 2473 1064 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12971 3734 1064 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12970 6561 6564 6313 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12969 6313 7825 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12968 11024 10027 6561 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12967 6560 6561 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12966 5281 5279 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12965 11024 6579 5281 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12964 5283 5281 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12963 10071 10694 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12962 11024 10702 10071 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12961 9974 10071 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12960 5039 5309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12959 11024 5295 5039 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12958 5038 5039 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12957 7651 8277 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12956 11024 8022 7651 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12955 7648 7651 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12954 11024 10418 9434 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12953 9433 9434 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12952 11024 9434 9433 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12951 11024 9434 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12950 11024 9434 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12949 11024 10418 9108 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12948 9107 9108 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12947 11024 9108 9107 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12946 11024 9108 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12945 11024 9108 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12944 11024 10419 10420 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12943 10418 10420 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12942 11024 10420 10418 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12941 11024 10420 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12940 11024 10420 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12939 11024 10698 9753 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12938 9753 10078 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12937 9753 10701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12936 11024 11072 9753 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12935 10080 9753 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12934 11024 10705 9736 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12933 9736 10414 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12932 9736 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12931 11024 10700 9736 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12930 9732 9736 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12929 11024 5550 3298 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12928 3298 3694 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12927 11024 3292 3298 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12926 3295 3298 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12925 3979 3976 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12924 11024 8092 3979 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12923 3993 3979 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12922 6491 6489 6302 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12921 6302 6819 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12920 11024 6490 6491 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12919 7766 6491 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12918 11024 1035 751 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12917 751 5809 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12916 11024 2578 751 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12915 750 751 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12914 7427 7437 7428 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12913 7428 9305 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12912 11024 8882 7427 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12911 7426 7427 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12910 11024 6278 3371 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12909 3371 3379 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12908 11024 5911 3371 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12907 3726 3371 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12906 9701 10350 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12905 11013 11028 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12904 10332 10999 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12903 7575 9046 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12902 7802 7813 7575 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12901 11024 8046 7802 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12900 10675 10990 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12899 6889 6879 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12898 6358 6261 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12897 4680 5863 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12896 5837 4673 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12895 6864 7516 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12894 11024 2582 2489 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12893 2489 2796 2493 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12892 2983 2986 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12891 2984 3860 2983 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12890 11024 4553 2984 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12889 3242 5535 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12888 11024 3007 3242 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12887 4586 4584 4386 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12886 4386 4925 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12885 11024 4926 4586 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12884 4942 4586 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12883 5055 5142 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12882 5144 5143 5055 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12881 11024 10915 5144 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12880 6113 6194 6404 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12879 11024 9379 6194 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12878 6114 6195 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12877 6404 9379 6114 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12876 11024 6765 6113 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12875 1319 1369 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12874 1317 1372 1363 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12873 11024 1396 1317 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12872 1372 1373 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12871 11024 5083 1373 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12870 11024 1388 1369 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12869 1370 1372 1319 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12868 1318 1373 1370 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12867 11024 1365 1318 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12866 1365 1370 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12865 1363 1373 1365 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12864 11024 1363 1396 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12863 1396 1363 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12862 5067 5264 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12861 5065 5263 5255 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12860 11024 5863 5065 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12859 5263 5265 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12858 11024 5262 5265 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12857 11024 5866 5264 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12856 5261 5263 5067 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12855 5066 5265 5261 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12854 11024 5256 5066 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12853 5256 5261 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12852 5255 5265 5256 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12851 11024 5255 5863 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12850 5863 5255 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12849 10015 10945 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12848 10015 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12847 11024 10027 10015 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12846 7538 10080 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12845 11024 10399 7538 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12844 1862 3413 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12843 10712 10786 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12842 10781 10780 10712 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12841 11024 10777 10781 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12840 1998 2657 1923 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12839 11024 3632 1923 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12838 1923 2984 1998 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12837 2406 1998 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12836 4295 4943 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12835 11024 3890 4295 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12834 2105 1865 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12833 11024 2114 2105 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12832 2104 1302 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12831 11024 6243 2104 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12830 2102 7069 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12829 11024 2099 2102 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12828 7685 10700 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12827 11024 10027 7685 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12826 1290 1287 1289 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12825 1289 1288 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12824 11024 1500 1290 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12823 1501 1290 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12822 11024 8677 8949 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12821 8677 8675 8676 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12820 8674 8678 8677 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12819 11024 8675 8678 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12818 8676 8679 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12817 11024 8954 8674 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12816 8949 8677 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12815 6890 10687 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12814 11024 6889 6890 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12813 6894 7167 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12812 11024 8056 6894 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12811 1374 7408 1320 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12810 1320 6387 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12809 11024 5500 1374 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12808 6394 1374 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12807 10592 10606 10593 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12806 10593 10608 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12805 11024 10825 10592 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12804 10591 10592 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12803 3246 3893 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12802 11024 4410 3246 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12801 8069 8247 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12800 8066 8197 8245 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12799 11024 8623 8066 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12798 8197 8248 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12797 11024 10914 8248 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12796 11024 8252 8247 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12795 8196 8197 8069 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12794 8067 8248 8196 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12793 11024 8192 8067 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12792 8192 8196 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12791 8245 8248 8192 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12790 11024 8245 8623 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12789 8623 8245 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12788 9556 9571 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12787 11024 9927 9556 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12786 10215 9556 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12785 11024 8687 8684 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12784 8687 8709 8688 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12783 8686 8689 8687 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12782 11024 8709 8689 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12781 8688 10680 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12780 11024 8685 8686 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12779 8684 8687 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12778 10608 4981 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12777 11024 7068 10608 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12776 3961 1874 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12775 11024 2109 3961 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12774 3728 3062 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12773 11024 3063 3728 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12772 9546 9559 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12771 11024 10018 9546 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12770 10004 9546 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12769 11024 10774 10563 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12768 10562 10563 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12767 11024 10800 10562 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12766 10561 10562 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12765 11024 10562 10561 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12764 9925 10825 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12763 9925 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12762 11024 10027 9925 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12761 10765 11038 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12760 10763 11040 11030 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12759 11024 11028 10763 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12758 11040 11041 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12757 11024 11051 11041 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12756 11024 11036 11038 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12755 11035 11040 10765 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12754 10764 11041 11035 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12753 11024 11032 10764 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12752 11032 11035 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12751 11030 11041 11032 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12750 11024 11030 11028 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12749 11028 11030 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12748 5615 5662 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12747 5613 5663 5655 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12746 11024 10567 5613 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12745 5663 5664 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12744 11024 10914 5664 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12743 11024 10186 5662 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12742 5660 5663 5615 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12741 5614 5664 5660 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12740 11024 5657 5614 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12739 5657 5660 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12738 5655 5664 5657 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12737 11024 5655 10567 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12736 10567 5655 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12735 7417 7419 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12734 11024 10018 7417 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12733 7585 7417 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12732 811 2472 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12731 1293 10256 811 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12730 11024 8713 1293 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12729 11024 6552 7154 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12728 6552 10687 6312 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12727 6311 6556 6552 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12726 11024 10687 6556 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12725 6312 10080 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12724 11024 7147 6311 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12723 7154 6552 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12722 11024 6542 6543 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12721 6542 10687 6310 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12720 6309 6544 6542 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12719 11024 10687 6544 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12718 6310 7165 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12717 11024 6545 6309 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12716 6543 6542 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12715 6305 6861 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12714 6518 7747 6305 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12713 11024 6862 6518 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12712 10392 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12711 10392 10414 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12710 11024 10705 10392 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12709 11024 10700 10392 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12708 8394 8437 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12707 8394 8395 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12706 11024 8403 8394 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12705 11024 10704 8394 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12704 7414 7655 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12703 7414 7484 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12702 11024 8122 7414 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12701 4256 10604 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12700 4255 8091 4256 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12699 11024 8885 4255 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12698 11024 9636 10078 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12697 9636 10684 9445 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12696 9444 9638 9636 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12695 11024 10684 9638 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12694 9445 9633 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12693 11024 9945 9444 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12692 10078 9636 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12691 11024 10303 10698 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12690 10303 10684 10117 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12689 10116 10304 10303 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12688 11024 10684 10304 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12687 10117 10312 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12686 11024 10662 10116 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12685 10698 10303 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12684 7540 7852 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12683 7540 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12682 11024 9432 7540 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12681 4274 4959 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12680 4274 5123 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12679 11024 5119 4274 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12678 11024 4954 4274 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12677 11024 7594 7596 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12676 8103 8893 7559 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12675 7559 7594 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12674 7559 7596 8103 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12673 11024 7590 7559 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12672 7590 8893 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12671 8121 8124 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12670 8121 8126 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12669 11024 8643 8121 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12668 11024 9987 8121 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12667 2530 5599 2529 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12666 5207 9308 2530 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12665 2530 3040 5207 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12664 2529 2736 2530 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12663 2529 5898 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12662 11024 3379 2529 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12661 11024 10051 10709 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12660 10051 10684 9956 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12659 9954 9957 10051 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12658 11024 10684 9957 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12657 9956 9955 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12656 11024 10302 9954 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12655 10709 10051 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12654 5927 5898 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12653 5927 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12652 11024 8922 5927 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12651 11024 7711 5927 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12650 11024 9547 9538 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12649 9538 9532 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12648 11024 9533 9538 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12647 9996 9538 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12646 8611 8613 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12645 8612 8615 8611 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12644 11024 8610 8612 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12643 7169 7177 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12642 11024 7176 7169 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12641 7167 7169 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12640 9085 11066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12639 11024 9083 9085 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12638 9081 9085 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12637 7083 7476 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12636 11024 9395 7083 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12635 7082 7083 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12634 10528 10772 10603 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12633 10527 10604 10528 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12632 10526 10892 10527 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12631 11024 10888 10526 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12630 10861 10603 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12629 3396 8126 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12628 3396 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12627 11024 7478 3396 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12626 11024 5607 3396 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12625 3151 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12624 3151 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12623 11024 7711 3151 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12622 11024 7478 3151 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12621 6293 9333 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12620 6435 7437 6293 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12619 11024 9321 6435 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12618 8772 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12617 9104 10083 8772 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12616 11024 10708 9104 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12615 11024 6789 6792 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12614 6788 7004 6790 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12613 6790 6789 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12612 6790 6792 6788 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12611 11024 6787 6790 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12610 6787 7004 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12609 2461 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12608 11024 9560 2461 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12607 2736 2461 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12606 1811 2417 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12605 1810 2418 1811 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12604 11024 2688 1810 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12603 10616 10614 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12602 10613 10615 10616 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12601 11024 10680 10613 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12600 11024 7421 7424 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12599 7422 9552 7423 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12598 7423 7421 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12597 7423 7424 7422 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12596 11024 7420 7423 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12595 7420 9552 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12594 4026 7527 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12593 11024 6574 4026 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12592 4023 4026 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12591 3720 4010 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12590 11024 5293 3720 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12589 3719 3720 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12588 11024 3033 1859 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12587 1859 7042 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12586 11024 2728 1859 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12585 1864 1859 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12584 11024 8643 7763 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12583 7763 8126 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12582 7763 8124 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12581 11024 9987 7763 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12580 8403 7763 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12579 11024 10701 8457 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12578 8457 10073 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12577 8457 9405 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12576 11024 10708 8457 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12575 8458 8457 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12574 11024 8126 7479 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12573 7479 7478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12572 7479 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12571 11024 8708 7479 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12570 7476 7479 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12569 11024 8661 5595 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12568 5595 5600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12567 11024 8643 5595 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12566 5593 5595 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12565 11024 3735 1896 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12564 1896 3734 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12563 11024 5293 1896 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12562 2208 1896 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12561 11024 9412 8149 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12560 8149 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12559 8149 10083 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12558 11024 10708 8149 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12557 8051 8149 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12556 11024 5131 3108 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12555 3108 3175 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12554 3607 3188 3108 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12553 3107 5124 3607 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12552 3108 3606 3107 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12551 6846 6848 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12550 6841 6849 6842 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12549 11024 10684 6841 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12548 6849 6850 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12547 11024 8048 6850 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12546 11024 6847 6848 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12545 6845 6849 6846 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12544 6844 6850 6845 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12543 11024 6843 6844 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12542 6843 6845 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12541 6842 6850 6843 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12540 11024 6842 10684 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12539 10684 6842 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12538 11024 8661 1580 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12537 1580 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12536 1580 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12535 11024 5599 1580 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12534 1575 1580 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12533 11024 9412 7528 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12532 7528 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12531 7528 9405 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12530 11024 10700 7528 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12529 7527 7528 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12528 11024 7478 7477 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12527 7477 8126 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12526 11024 10028 7477 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12525 8100 7477 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12524 3355 7041 3150 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_12523 3149 3714 3355 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_12522 11024 6221 3149 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_12521 3150 4014 11024 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_12520 10786 10783 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12519 11024 10915 10786 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12518 3005 3004 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12517 3230 5743 3005 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12516 11024 3219 3230 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12515 4292 4291 4293 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12514 4293 4925 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12513 11024 4926 4292 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12512 4290 4292 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12511 3747 3749 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12510 3743 3750 3744 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12509 11024 4066 3743 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12508 3750 3751 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12507 11024 5262 3751 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12506 11024 4476 3749 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12505 3748 3750 3747 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12504 3746 3751 3748 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12503 11024 3745 3746 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12502 3745 3748 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12501 3744 3751 3745 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12500 11024 3744 4066 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12499 4066 3744 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12498 9387 9389 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12497 9383 9391 9384 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12496 11024 9382 9383 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12495 9391 9390 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12494 11024 11051 9390 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12493 11024 9394 9389 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12492 9388 9391 9387 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12491 9386 9390 9388 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12490 11024 9385 9386 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12489 9385 9388 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12488 9384 9390 9385 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12487 11024 9384 9382 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12486 9382 9384 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12485 2465 2576 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12484 2464 2469 2465 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12483 11024 4327 2464 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12482 11024 8297 8170 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12481 8171 9313 8291 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12480 8169 8699 8171 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12479 8170 8930 8169 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12478 11024 8918 8173 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12477 8174 8885 8290 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12476 8172 8642 8174 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12475 8173 9304 8172 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12474 707 1495 709 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12473 709 1494 710 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12472 710 708 709 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12471 707 706 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12470 11024 1489 707 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12469 709 711 707 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12468 2435 710 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12467 11024 5240 4987 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12466 4987 8409 4988 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12465 4986 4988 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12464 6486 8691 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12463 6486 6487 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12462 11024 6483 6486 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12461 6506 6503 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12460 6506 7498 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12459 11024 10027 6506 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12458 8765 11066 8766 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12457 8766 9977 8765 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12456 11024 8768 8766 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12455 5674 7690 5631 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12454 5631 5671 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12453 11024 6121 5674 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12452 5670 5674 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12451 5640 6867 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12450 8633 5809 5640 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12449 11024 8092 8633 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12448 4486 4488 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12447 11024 6376 4486 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12446 5143 4486 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12445 1850 1852 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12444 1846 1853 1847 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12443 11024 7474 1846 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12442 1853 1854 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12441 11024 2446 1854 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12440 11024 2074 1852 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12439 1851 1853 1850 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12438 1849 1854 1851 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12437 11024 1848 1849 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12436 1848 1851 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12435 1847 1854 1848 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12434 11024 1847 7474 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12433 7474 1847 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12432 777 864 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12431 775 863 859 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12430 11024 8885 775 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12429 863 865 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12428 11024 5083 865 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12427 11024 867 864 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12426 860 863 777 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12425 776 865 860 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12424 11024 861 776 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12423 861 860 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12422 859 865 861 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12421 11024 859 8885 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12420 8885 859 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12419 6571 6569 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12418 6571 8767 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12417 11024 6585 6571 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12416 1841 1504 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12415 11024 7701 1841 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12414 3710 1542 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12413 11024 4981 3710 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12412 3982 4665 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12411 11024 4658 3982 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12410 1330 1420 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12409 1328 1421 1415 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12408 11024 7425 1328 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12407 1421 1422 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12406 11024 2673 1422 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12405 11024 1816 1420 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12404 1418 1421 1330 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12403 1329 1422 1418 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12402 11024 1416 1329 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12401 1416 1418 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12400 1415 1422 1416 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12399 11024 1415 7425 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12398 7425 1415 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12397 10016 10017 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12396 11024 10018 10016 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12395 10009 10016 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12394 8914 8913 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12393 11024 8915 8914 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12392 8912 8914 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12391 3046 4012 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12390 3046 3047 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12389 11024 8709 3046 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12388 3047 3706 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12387 3047 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12386 11024 6277 3047 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12385 2575 2121 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12384 2575 2114 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12383 11024 6243 2575 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12382 1870 3092 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12381 1870 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12380 11024 5911 1870 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12379 8346 10027 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12378 8336 9335 8105 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12377 8105 8340 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12376 11024 8337 8111 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12375 8111 8341 8108 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12374 8108 8346 8336 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12373 8336 10027 8110 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12372 8110 10231 8111 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12371 11024 8340 8337 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_12370 9341 8336 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12369 11058 10699 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12368 11058 11066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12367 11024 10697 11058 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12366 10706 11072 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12365 10706 10705 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12364 11024 11076 10706 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12363 3738 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12362 3738 3719 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12361 11024 3967 3738 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12360 4327 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12359 4327 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12358 11024 6277 4327 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12357 6174 6286 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12356 6175 6902 6174 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12355 11024 6285 6175 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12354 4946 5159 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12353 11024 6127 4946 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12352 4944 4946 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12351 10247 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12350 10247 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12349 11024 9309 10247 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12348 11024 8930 10247 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12347 1350 1520 1521 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12346 1351 7082 1350 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12345 11024 1537 1351 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12344 1519 1521 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12343 9603 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12342 9603 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12341 11024 10029 9603 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12340 11024 10945 9603 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12339 6902 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12338 6902 9080 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12337 11024 9057 6902 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12336 11024 9433 6902 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12335 6282 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12334 6282 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12333 11024 6278 6282 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12332 11024 5911 6282 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12331 6901 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12330 6901 9057 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12329 11024 8746 6901 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12328 11024 9433 6901 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12327 5153 11018 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12326 5153 5728 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12325 11024 5727 5153 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12324 11024 10566 10193 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12323 10193 10218 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12322 10193 10542 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12321 11024 10541 10193 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12320 10547 10193 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12319 6878 10399 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12318 11024 8746 6878 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12317 6877 6878 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12316 9594 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12315 9594 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12314 11024 10029 9594 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12313 11024 10924 9594 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12312 2165 7042 1943 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_12311 1942 3714 2165 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_12310 11024 6220 1942 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_12309 1943 4014 11024 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_12308 2540 2581 2779 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12307 2541 2582 2540 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12306 11024 3716 2541 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12305 4037 2779 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12304 3889 5153 3772 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12303 3772 5718 3889 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12302 11024 6213 3772 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12301 5048 5098 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12300 5100 6195 5048 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12299 11024 10915 5100 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12298 8269 8848 8164 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12297 11024 8267 8164 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12296 8164 8834 8269 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12295 9298 8269 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12294 4632 4983 4392 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12293 4392 6259 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12292 11024 5194 4632 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12291 4631 4632 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12290 11024 1075 1072 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12289 5600 1072 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12288 11024 1072 5600 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12287 11024 1072 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12286 11024 1072 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12285 11024 1075 1076 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12284 6276 1076 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12283 11024 1076 6276 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12282 11024 1076 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12281 11024 1076 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12280 11024 770 771 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12279 1075 771 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12278 11024 771 1075 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12277 11024 771 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12276 11024 771 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12275 11024 4356 3409 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12274 8922 3409 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12273 11024 3409 8922 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12272 11024 3409 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12271 11024 3409 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12270 11024 4356 3742 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12269 9309 3742 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12268 11024 3742 9309 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12267 11024 3742 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12266 11024 3742 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12265 11024 4356 3736 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12264 10031 3736 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12263 11024 3736 10031 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12262 11024 3736 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12261 11024 3736 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12260 11024 4356 4357 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12259 5583 4357 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12258 11024 4357 5583 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12257 11024 4357 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12256 11024 4357 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12255 11024 3410 3412 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12254 4356 3412 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12253 11024 3412 4356 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12252 11024 3412 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12251 11024 3412 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12250 746 4995 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12249 11024 1545 746 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12248 745 746 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12247 1827 7701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12246 11024 1826 1827 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12245 2680 1827 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12244 11024 9087 8761 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12243 8761 9433 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12242 11024 9716 8761 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12241 8760 8761 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12240 3732 3735 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12239 11024 9597 3732 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12238 4031 3732 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12237 8883 9347 8785 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12236 8785 9633 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12235 11024 9306 8883 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12234 8882 8883 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12233 11024 7514 7515 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12232 7515 7721 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12231 7515 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12230 11024 10197 7515 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12229 10697 7515 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12228 4718 4717 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12227 11024 5926 4718 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12226 4720 4718 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12225 11024 9314 3350 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12224 3350 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12223 11024 3703 3350 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12222 3712 3350 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12221 11024 5777 5781 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12220 5781 5782 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12219 11024 5774 5781 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12218 5776 5781 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12217 8129 8392 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12216 8125 8222 8385 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12215 11024 8388 8125 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12214 8222 8393 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12213 11024 10638 8393 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12212 11024 8390 8392 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12211 8221 8222 8129 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12210 8127 8393 8221 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12209 11024 8220 8127 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12208 8220 8221 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12207 8385 8393 8220 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12206 11024 8385 8388 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12205 8388 8385 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12204 11024 7678 1566 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12203 1566 2133 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12202 1566 7514 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12201 11024 5293 1566 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12200 1890 1566 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12199 3703 2473 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12198 3706 8124 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12197 1055 4066 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12196 10302 10662 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12195 9945 10289 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12194 9639 9947 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12193 11024 10378 10377 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12192 10377 11075 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12191 11024 10686 10377 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12190 10704 10377 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12189 11024 7041 4613 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12188 4613 5809 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12187 4613 10018 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12186 11024 7042 4613 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12185 5202 4613 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12184 11024 9560 5559 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12183 5559 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12182 5559 6275 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12181 11024 6867 5559 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12180 8318 5559 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12179 5702 5684 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12178 11024 5518 5702 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12177 1226 1227 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12176 1221 1228 1222 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12175 11024 1813 1221 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12174 1228 1229 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12173 11024 2673 1229 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12172 11024 1230 1227 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12171 1225 1228 1226 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12170 1223 1229 1225 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12169 11024 1224 1223 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12168 1224 1225 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12167 1222 1229 1224 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12166 11024 1222 1813 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12165 1813 1222 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12164 10045 10595 9944 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12163 9944 10596 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12162 11024 10680 10045 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12161 10042 10045 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12160 7719 9395 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12159 5671 7601 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12158 3804 7418 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12157 7411 7425 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12156 11024 3413 290 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12155 290 2473 487 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12154 11024 4066 774 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12153 774 4070 773 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12152 11024 3382 2789 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12151 2789 2597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12150 2789 2592 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12149 11024 2791 2789 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12148 5015 2789 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12147 4919 4555 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12146 11024 4410 4919 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12145 10768 11053 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12144 10766 11052 11044 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12143 11024 11042 10766 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12142 11052 11056 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12141 11024 11051 11056 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12140 11024 11059 11053 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12139 11049 11052 10768 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12138 10767 11056 11049 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12137 11024 11048 10767 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12136 11048 11049 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12135 11044 11056 11048 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12134 11024 11044 11042 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12133 11042 11044 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12132 9586 10924 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12131 9586 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12130 11024 9582 9586 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12129 7053 8644 6921 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12128 6921 9605 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12127 11024 7061 7053 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12126 7447 7053 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12125 11024 3983 2535 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12124 2535 2761 2751 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12123 2752 2751 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12122 11024 3983 2534 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12121 2534 2753 2749 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_12120 2750 2749 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12119 1855 7701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12118 11024 1844 1855 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12117 9920 10772 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12116 10546 10564 9920 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12115 11024 9994 10546 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12114 4584 5159 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12113 11024 6127 4584 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12112 9283 9285 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12111 9279 9286 9280 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12110 11024 9287 9279 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12109 9286 9288 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12108 11024 10914 9288 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12107 11024 9292 9285 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12106 9284 9286 9283 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12105 9282 9288 9284 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12104 11024 9281 9282 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12103 9281 9284 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12102 9280 9288 9281 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12101 11024 9280 9287 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12100 9287 9280 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12099 11024 8320 8670 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12098 8320 8327 8178 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12097 8177 8321 8320 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12096 11024 8327 8321 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12095 8178 8328 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12094 11024 8694 8177 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12093 8670 8320 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12092 11024 8102 8328 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12091 8102 8026 8027 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12090 8025 8028 8102 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12089 11024 8026 8028 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12088 8027 10257 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12087 11024 8642 8025 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12086 8328 8102 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12085 6917 10604 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12084 7023 8091 6917 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12083 11024 8297 7023 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12082 4012 3379 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12081 11024 9597 4012 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12080 1815 8012 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12079 11024 1822 1815 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12078 3043 3698 3042 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12077 3042 3040 3041 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12076 3041 9597 3043 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12075 3043 3967 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12074 11024 5599 3043 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12073 3695 3041 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12072 3664 6811 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12071 11024 4311 3664 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12070 10760 11010 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12069 10758 11009 11001 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12068 11024 10999 10758 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12067 11009 11011 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12066 11024 11051 11011 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12065 11024 11006 11010 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12064 11007 11009 10760 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12063 10759 11011 11007 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12062 11024 11005 10759 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12061 11005 11007 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12060 11001 11011 11005 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12059 11024 11001 10999 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12058 10999 11001 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12057 8273 9296 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12056 11024 9297 8273 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12055 8865 8273 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12054 7438 7445 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12053 11024 7667 7438 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12052 9297 7438 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12051 8929 10700 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12050 11024 10027 8929 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12049 10577 8929 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12048 11024 8706 8977 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12047 8706 8712 8705 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12046 8704 8707 8706 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12045 11024 8712 8707 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12044 8705 8970 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12043 11024 8703 8704 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12042 8977 8706 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12041 11024 8366 8703 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12040 8366 8709 8182 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12039 8181 8373 8366 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12038 11024 8709 8373 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12037 8182 10594 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12036 11024 8697 8181 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_12035 8703 8366 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12034 2741 3379 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12033 11024 5918 2741 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12032 10694 10708 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12031 10694 10414 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12030 11024 10705 10694 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12029 9547 10854 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12028 9547 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12027 11024 10027 9547 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12026 3822 3817 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12025 3822 4959 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12024 11024 4954 3822 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12023 11024 4915 3822 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12022 4320 4323 4319 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12021 4319 5539 4320 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12020 11024 6213 4319 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12019 2508 2624 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12018 2506 2623 2614 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12017 11024 8090 2506 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12016 2623 2622 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12015 11024 5083 2622 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_12014 11024 4881 2624 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12013 2555 2623 2508 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12012 2507 2622 2555 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12011 11024 2554 2507 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12010 2554 2555 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12009 2614 2622 2554 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_12008 11024 2614 8090 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12007 8090 2614 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_12006 9988 9989 9917 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12005 9917 10218 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12004 11024 9987 9988 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12003 10179 9988 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_12002 6387 7655 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12001 6387 7415 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_12000 11024 9304 6387 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11999 11024 8072 7583 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11998 11024 10197 7584 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11997 7583 7584 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11996 4684 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11995 4684 7721 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11994 11024 7514 4684 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11993 11024 6163 4684 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11992 11024 5728 3631 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11991 3631 5727 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11990 11024 10312 3631 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11989 3630 3631 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11988 11024 5554 5555 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11987 8424 5555 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11986 11024 5555 8424 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11985 11024 5555 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11984 11024 5555 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11983 11024 5199 5201 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11982 8145 5201 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11981 11024 5201 8145 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11980 11024 5201 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11979 11024 5201 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11978 11024 8424 8425 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11977 11051 8425 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11976 11024 8425 11051 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11975 11024 8425 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11974 11024 8425 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11973 11024 8424 8422 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11972 10638 8422 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11971 11024 8422 10638 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11970 11024 8422 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11969 11024 8422 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11968 11024 8424 8147 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11967 8048 8147 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11966 11024 8147 8048 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11965 11024 8147 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11964 11024 8147 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11963 11024 8145 8146 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11962 8047 8146 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11961 11024 8146 8047 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11960 11024 8146 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11959 11024 8146 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11958 11024 8424 8289 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11957 10914 8289 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11956 11024 8289 10914 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11955 11024 8289 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11954 11024 8289 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11953 11024 8424 8287 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11952 8286 8287 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11951 11024 8287 8286 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11950 11024 8287 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11949 11024 8287 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11948 11024 1958 1960 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11947 7594 7484 1920 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11946 1920 1958 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11945 1920 1960 7594 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11944 11024 1954 1920 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11943 1954 7484 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11942 11065 11071 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11941 11024 11061 11065 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11940 11063 11065 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11939 11024 6819 5813 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11938 5814 5813 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11937 11024 5811 5814 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11936 6233 5814 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11935 11024 5814 6233 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11934 11024 4070 1082 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11933 1080 1082 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11932 11024 4066 1080 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11931 1079 1080 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11930 11024 1080 1079 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11929 4250 4058 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11928 4250 5295 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11927 11024 4057 4250 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11926 4995 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11925 4995 7721 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11924 11024 7514 4995 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11923 11024 6879 4995 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11922 11024 4508 3629 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11921 3629 4939 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11920 11024 5131 3629 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11919 3628 3629 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11918 5119 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11917 5119 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11916 11024 5719 5119 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11915 11024 8623 5119 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11914 11024 7652 8093 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11913 11024 9987 7654 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11912 8093 7654 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11911 7805 8052 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11910 7805 10399 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11909 11024 9051 7805 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11908 11024 9716 7805 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11907 8808 9046 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11906 9030 9029 8808 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11905 11024 9028 9030 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11904 6382 7410 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11903 11024 6379 6382 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11902 6381 6382 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11901 6799 7460 6802 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11900 6800 10604 6799 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11899 6801 10892 6800 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11898 11024 10888 6801 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11897 6798 6802 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11896 11024 5191 4994 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11895 5012 7484 4993 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11894 4993 5191 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11893 4993 4994 5012 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11892 11024 4992 4993 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11891 4992 7484 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11890 11024 6784 6786 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11889 6789 9605 6785 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11888 6785 6784 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11887 6785 6786 6789 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11886 11024 6783 6785 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11885 6783 9605 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11884 10108 10269 10107 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11883 10107 10256 10263 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11882 10263 10258 10108 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11881 10108 10621 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11880 11024 10259 10108 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11879 10255 10263 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11878 7030 7033 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11877 11024 7439 7030 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11876 7027 7030 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11875 4982 4981 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11874 11024 7068 4982 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11873 5214 4982 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11872 2455 5809 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11871 11024 7041 2455 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11870 2454 2455 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11869 769 4066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11868 11024 4070 769 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11867 767 769 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11866 3365 3735 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11865 11024 3734 3365 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11864 3722 3365 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11863 8168 8617 8167 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11862 8652 10838 8168 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11861 8168 8635 8652 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11860 8167 8636 8168 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11859 8167 8885 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11858 11024 8633 8167 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11857 4533 5525 4380 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11856 4380 5519 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11855 11024 4553 4533 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11854 4530 4533 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11853 5537 7437 5538 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11852 5538 9605 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11851 11024 9323 5537 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11850 5535 5537 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11849 11024 3956 3291 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11848 3291 3295 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11847 11024 3285 3291 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11846 3288 3291 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11845 9356 9358 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11844 9351 9360 9352 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11843 11024 9350 9351 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11842 9360 9359 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11841 11024 10638 9359 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11840 11024 9355 9358 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11839 9357 9360 9356 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11838 9353 9359 9357 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11837 11024 9354 9353 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11836 9354 9357 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11835 9352 9359 9354 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11834 11024 9352 9350 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11833 9350 9352 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11832 9400 9402 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11831 9396 9404 9397 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11830 11024 9395 9396 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11829 9404 9403 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11828 11024 11051 9403 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11827 11024 9411 9402 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11826 9401 9404 9400 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11825 9399 9403 9401 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11824 11024 9398 9399 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11823 9398 9401 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11822 9397 9403 9398 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11821 11024 9397 9395 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11820 9395 9397 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11819 6300 6477 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11818 6478 10027 6300 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11817 11024 6499 6478 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11816 11024 11076 7524 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11815 7524 9412 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11814 11024 10700 7524 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11813 7523 7524 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11812 10082 10083 9981 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11811 9981 10698 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11810 11024 10708 10082 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11809 9980 10082 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11808 4310 4955 4243 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11807 11024 4952 4243 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11806 4243 4631 4310 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11805 4925 4310 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11804 3002 3000 3001 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11803 3001 5753 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11802 11024 3236 3002 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11801 2998 3002 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11800 784 889 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11799 782 888 884 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11798 11024 902 782 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11797 888 890 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11796 11024 2673 890 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11795 11024 892 889 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11794 885 888 784 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11793 783 890 885 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11792 11024 886 783 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11791 886 885 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11790 884 890 886 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11789 11024 884 902 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11788 902 884 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11787 10586 10591 10836 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11786 10587 10584 10586 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11785 11024 10585 10587 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11784 1327 2417 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11783 1409 2418 1327 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11782 11024 10888 1409 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11781 11024 5901 2195 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11780 2195 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11779 2195 5898 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11778 11024 7711 2195 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11777 2589 2195 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11776 6591 7848 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11775 11024 7852 6591 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11774 10545 10555 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11773 11024 10547 10545 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11772 11024 7484 3155 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11771 11024 9987 1791 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11770 3155 1791 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11769 8742 8743 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11768 8737 8745 8738 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11767 11024 8748 8737 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11766 8745 8744 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11765 11024 11051 8744 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11764 11024 8751 8743 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11763 8740 8745 8742 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11762 8739 8744 8740 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11761 11024 8741 8739 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11760 8741 8740 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11759 8738 8744 8741 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11758 11024 8738 8748 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11757 8748 8738 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11756 9098 10083 8815 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11755 8815 10701 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11754 11024 10708 9098 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11753 9426 9098 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11752 2520 3009 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11751 3003 3008 2520 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11750 11024 4325 3003 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11749 4929 5181 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11748 11024 5842 4929 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11747 3871 4617 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11746 3871 5521 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11745 11024 5522 3871 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11744 3017 3020 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11743 3013 3021 3014 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11742 11024 7037 3013 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11741 3021 3022 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11740 11024 5083 3022 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11739 11024 3019 3020 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11738 3018 3021 3017 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11737 3016 3022 3018 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11736 11024 3015 3016 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11735 3015 3018 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11734 3014 3022 3015 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11733 11024 3014 7037 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11732 7037 3014 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11731 1248 1504 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11730 11024 1495 1248 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11729 5002 4997 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11728 11024 4453 5002 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11727 10560 10571 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11726 11024 10559 10560 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11725 5521 10024 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11724 5521 5728 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11723 11024 5727 5521 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11722 4266 4265 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11721 4257 4260 4258 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11720 11024 9304 4257 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11719 4260 4268 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11718 11024 5083 4268 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11717 11024 5494 4265 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11716 4262 4260 4266 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11715 4263 4268 4262 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11714 11024 4261 4263 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11713 4261 4262 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11712 4258 4268 4261 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11711 11024 4258 9304 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11710 9304 4258 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11709 8649 8648 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11708 11024 10018 8649 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11707 8647 8649 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11706 7533 10399 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11705 7533 8155 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11704 11024 9421 7533 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11703 1284 1504 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11702 11024 1494 1284 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11701 3709 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11700 3709 8661 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11699 11024 5600 3709 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11698 7161 9080 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11697 11024 8453 7161 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11696 2407 5490 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11695 2409 3688 2405 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11694 2405 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11693 11024 2404 2411 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11692 2411 2406 2408 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11691 2408 2407 2409 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11690 2409 5490 2410 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11689 2410 2985 2411 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11688 11024 4929 2404 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11687 2403 2409 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11686 2650 5490 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11685 2642 4142 2514 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11684 2514 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11683 11024 2645 2517 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11682 2517 2646 2515 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11681 2515 2650 2642 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11680 2642 5490 2516 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11679 2516 2984 2517 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11678 11024 4929 2645 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11677 2962 2642 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11676 4282 5521 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11675 11024 5522 4282 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11674 4281 4282 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11673 1916 2059 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11672 1914 2060 2053 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11671 11024 7450 1914 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11670 2060 2061 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11669 11024 2446 2061 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11668 11024 2062 2059 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11667 2057 2060 1916 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11666 1915 2061 2057 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11665 11024 2054 1915 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11664 2054 2057 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11663 2053 2061 2054 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11662 11024 2053 7450 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11661 7450 2053 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11660 9993 8824 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11659 9993 8831 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11658 11024 8833 9993 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11657 11024 8817 9993 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11656 4253 8817 4252 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11655 4252 8824 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11654 11024 10915 4253 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11653 8313 4253 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11652 7828 9716 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11651 7828 8458 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11650 11024 9433 7828 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11649 11024 10652 9939 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11648 11024 10774 9940 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11647 9939 9940 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11646 6285 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11645 6285 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11644 11024 6278 6285 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11643 11024 5918 6285 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11642 8813 10073 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11641 9080 10701 8813 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11640 11024 10708 9080 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11639 1828 2692 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11638 2426 2691 1828 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11637 11024 4325 2426 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11636 11024 5728 2768 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11635 2768 5727 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11634 11024 10257 2768 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11633 2986 2768 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11632 2388 2974 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11631 2390 5490 2387 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11630 2387 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11629 11024 2386 2391 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11628 2391 2632 2389 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11627 2389 2388 2390 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11626 2390 2974 2392 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11625 2392 3621 2391 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11624 11024 4929 2386 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11623 2385 2390 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11622 1988 2974 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11621 1985 1993 1904 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11620 1904 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11619 11024 1977 1907 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11618 1907 2640 1905 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11617 1905 1988 1985 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11616 1985 2974 1906 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11615 1906 3625 1907 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11614 11024 4929 1977 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_11613 2967 1985 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11612 10017 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11611 10017 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11610 11024 10029 10017 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11609 11024 10641 10017 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11608 4015 4012 3794 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11607 3794 4014 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11606 11024 4013 4015 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11605 4701 4015 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11604 11024 9925 9531 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11603 9531 9526 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11602 11024 9540 9531 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11601 10206 9531 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11600 11024 2470 2471 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11599 2471 2578 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11598 11024 8713 2471 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11597 5818 2471 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11596 2372 3714 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11595 2479 4012 2372 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11594 2371 2480 2479 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11593 11024 4014 2371 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11592 3062 2479 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11591 4397 4451 4681 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11590 4398 4452 4397 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11589 11024 4450 4398 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11588 4708 4681 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11587 8023 8318 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11586 8022 8316 8023 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11585 11024 8694 8022 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11584 11024 4277 4270 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11583 5098 4272 4273 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11582 4273 4277 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11581 4273 4270 5098 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11580 11024 4271 4273 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11579 4271 4272 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11578 11024 5608 5291 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11577 9560 5291 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11576 11024 5291 9560 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11575 11024 5291 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11574 11024 5291 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11573 11024 5608 5609 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11572 9020 5609 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11571 11024 5609 9020 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11570 11024 5609 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11569 11024 5609 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11568 11024 5608 5597 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11567 10029 5597 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11566 11024 5597 10029 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11565 11024 5597 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11564 11024 5597 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11563 11024 5035 5036 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11562 5608 5036 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11561 11024 5036 5608 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11560 11024 5036 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11559 11024 5036 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11558 11024 762 761 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11557 5898 761 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11556 11024 761 5898 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11555 11024 761 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11554 11024 761 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11553 11024 762 763 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11552 5911 763 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11551 11024 763 5911 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11550 11024 763 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11549 11024 763 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11548 11024 762 760 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11547 6275 760 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11546 11024 760 6275 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11545 11024 760 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11544 11024 760 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11543 11024 494 496 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11542 762 496 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11541 11024 496 762 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11540 11024 496 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11539 11024 496 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11538 7568 7719 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11537 8106 7701 7568 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11536 11024 7702 8106 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11535 7820 8054 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11534 11024 7835 7820 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11533 8151 7820 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11532 11024 10073 9422 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11531 9422 10701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11530 11024 10700 9422 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11529 9421 9422 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11528 10102 10568 10233 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11527 10101 10604 10102 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11526 10100 10892 10101 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11525 11024 10888 10100 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11524 10279 10233 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11523 6138 8654 6218 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11522 6139 10604 6138 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11521 6136 10892 6139 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11520 11024 10888 6136 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11519 6137 6218 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11518 10553 10780 10552 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11517 10552 10551 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11516 11024 10774 10553 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11515 10550 10553 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11514 11024 1067 765 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11513 5918 765 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11512 11024 765 5918 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11511 11024 765 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11510 11024 765 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11509 11024 1067 764 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11508 5599 764 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11507 11024 764 5599 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11506 11024 764 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11505 11024 764 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11504 11024 1067 1069 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11503 7678 1069 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11502 11024 1069 7678 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11501 11024 1069 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11500 11024 1069 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11499 11024 499 498 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11498 1067 498 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11497 11024 498 1067 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11496 11024 498 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11495 11024 498 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11494 11024 1610 1612 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11493 6277 1612 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11492 11024 1612 6277 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11491 11024 1612 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11490 11024 1612 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11489 11024 1610 1316 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11488 7711 1316 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11487 11024 1316 7711 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11486 11024 1316 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11485 11024 1316 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11484 11024 1610 1312 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11483 5719 1312 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11482 11024 1312 5719 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11481 11024 1312 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11480 11024 1312 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11479 11024 1079 1078 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11478 1610 1078 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11477 11024 1078 1610 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11476 11024 1078 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11475 11024 1078 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11474 8655 8654 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11473 8831 10564 8655 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11472 11024 8912 8831 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11471 11024 10709 9060 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11470 9060 10083 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11469 11024 10700 9060 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11468 9083 9060 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11467 3061 3062 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11466 11024 3063 3061 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11465 3070 3061 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11464 3383 3379 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11463 11024 5918 3383 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11462 4038 3383 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11461 3740 3738 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11460 11024 3739 3740 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11459 4717 3740 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11458 11024 5581 5250 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11457 5901 5250 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11456 11024 5250 5901 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11455 11024 5250 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11454 11024 5250 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11453 11024 5581 5582 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11452 6278 5582 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11451 11024 5582 6278 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11450 11024 5582 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11449 11024 5582 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11448 11024 5577 5578 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11447 5581 5578 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11446 11024 5578 5581 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11445 11024 5578 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11444 11024 5578 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11443 9463 9610 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11442 10044 9609 9463 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11441 11024 9613 10044 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11440 2539 4014 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11439 2769 3033 2539 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11438 2538 3057 2769 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11437 11024 3714 2538 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11436 3065 2769 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11435 8158 10710 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11434 11024 11072 8158 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11433 8062 8158 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11432 3342 5600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11431 11024 6277 3342 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11430 3704 3342 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11429 11024 3735 1895 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11428 1895 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11427 11024 5293 1895 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11426 1898 1895 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11425 11024 472 456 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11424 456 1545 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11423 11024 6261 456 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11422 451 456 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11421 11024 10771 10777 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11420 11024 10915 8818 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11419 10777 8818 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11418 1338 1454 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11417 1336 1453 1445 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11416 11024 2432 1336 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11415 1453 1455 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11414 11024 2446 1455 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11413 11024 1461 1454 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11412 1451 1453 1338 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11411 1337 1455 1451 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11410 11024 1449 1337 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11409 1449 1451 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11408 1445 1455 1449 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11407 11024 1445 2432 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11406 2432 1445 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11405 7574 9033 7770 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11404 7573 8748 7574 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11403 11024 8407 7573 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11402 7570 8388 7740 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11401 7569 7739 7570 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11400 11024 8409 7569 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11399 6244 6518 6153 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11398 6153 6851 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11397 11024 6243 6244 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11396 6152 6244 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11395 11024 10378 9420 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11394 9420 9419 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11393 9420 11075 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11392 11024 11072 9420 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11391 9418 9420 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11390 7691 7690 7564 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11389 7564 7689 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11388 11024 10255 7691 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11387 8096 7691 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11386 7019 7450 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11385 7606 7611 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11384 7689 7466 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11383 3624 3837 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11382 3625 4567 3624 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11381 11024 4553 3625 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11380 3873 4539 3770 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11379 3770 3875 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11378 11024 3872 3873 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11377 6201 3873 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11376 8045 8141 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11375 8043 8142 8136 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11374 11024 8409 8043 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11373 8142 8144 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11372 11024 10638 8144 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11371 11024 8734 8141 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11370 8139 8142 8045 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11369 8044 8144 8139 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11368 11024 8138 8044 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11367 8138 8139 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11366 8136 8144 8138 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11365 11024 8136 8409 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11364 8409 8136 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11363 2468 3337 2469 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11362 2467 2466 2468 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11361 11024 2750 2467 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11360 1291 4981 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11359 11024 1881 1291 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11358 7475 7474 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11357 7452 7037 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11356 10575 10800 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11355 10839 10838 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11354 10772 10771 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11353 10619 4254 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11352 11024 5898 1902 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11351 1902 5600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11350 1902 6277 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11349 11024 5607 1902 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11348 2211 1902 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11347 11024 9309 3085 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11346 3085 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11345 3085 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11344 11024 8126 3085 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11343 3084 3085 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11342 5140 6214 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11341 11024 6215 5140 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11340 1343 1479 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11339 1341 1480 1472 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11338 11024 1844 1341 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11337 1480 1481 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11336 11024 2446 1481 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11335 11024 1839 1479 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11334 1477 1480 1343 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11333 1342 1481 1477 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11332 11024 1474 1342 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11331 1474 1477 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11330 1472 1481 1474 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11329 11024 1472 1844 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11328 1844 1472 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11327 6162 6269 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11326 6160 6270 6267 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11325 11024 6493 6160 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11324 6270 6272 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11323 11024 8048 6272 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11322 11024 6273 6269 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11321 6268 6270 6162 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11320 6161 6272 6268 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11319 11024 6271 6161 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11318 6271 6268 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11317 6267 6272 6271 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11316 11024 6267 6493 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11315 6493 6267 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11314 6232 4653 4396 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_11313 4395 7678 6232 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_11312 11024 5911 4395 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_11311 4396 4654 11024 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_11310 6827 6240 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11309 11024 6486 6827 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11308 6537 8733 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11307 11024 6358 6537 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11306 6489 5811 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11305 5059 5552 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11304 5757 10606 5059 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11303 11024 9304 5757 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11302 11024 2958 2956 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11301 2958 9379 2960 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11300 2959 2961 2958 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11299 11024 9379 2961 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11298 2960 2964 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11297 11024 2957 2959 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11296 2956 2958 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11295 4936 6431 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11294 11024 3213 4936 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11293 10011 10641 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11292 10011 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11291 11024 10027 10011 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11290 11024 8701 8697 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11289 8701 8708 8700 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11288 8698 8702 8701 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11287 11024 8708 8702 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11286 8700 8699 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11285 11024 8983 8698 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11284 8697 8701 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11283 4029 7527 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11282 11024 6574 4029 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11281 2427 6140 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11280 11024 2426 2427 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11279 3652 3651 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11278 11024 4314 3652 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11277 1799 3611 1797 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11276 1797 1796 1798 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11275 1798 2637 1799 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11274 1799 1964 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11273 11024 2962 1799 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11272 1805 1798 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11271 8779 8858 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11270 8777 8859 8850 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11269 11024 8848 8777 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11268 8859 8860 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11267 11024 10914 8860 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11266 11024 8856 8858 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11265 8855 8859 8779 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11264 8778 8860 8855 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11263 11024 8852 8778 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11262 8852 8855 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11261 8850 8860 8852 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11260 11024 8850 8848 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11259 8848 8850 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11258 5641 5816 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11257 6240 6150 5641 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11256 11024 7480 6240 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11255 11024 8727 8724 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11254 8727 8733 8730 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11253 8726 8729 8727 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11252 11024 8733 8729 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11251 8730 8728 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11250 11024 8725 8726 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11249 8724 8727 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11248 6906 9747 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11247 6906 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11246 11024 10704 6906 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11245 6793 7648 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11244 11024 6791 6793 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11243 3029 5809 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11242 11024 7041 3029 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11241 5194 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11240 5194 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11239 11024 10029 5194 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11238 11024 5191 5194 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11237 10755 10986 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11236 10753 10985 10979 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11235 11024 10990 10753 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11234 10985 10987 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11233 11024 11051 10987 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11232 11024 10989 10986 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11231 10984 10985 10755 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11230 10754 10987 10984 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11229 11024 10980 10754 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11228 10980 10984 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11227 10979 10987 10980 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11226 11024 10979 10990 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11225 10990 10979 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11224 10612 10611 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11223 11024 10613 10612 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11222 10610 10612 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11221 7562 7633 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11220 7634 9297 7562 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11219 11024 7631 7634 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11218 8112 8126 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11217 8112 8038 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11216 11024 7721 8112 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11215 11024 9308 8112 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11214 11024 7512 7509 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11213 7512 10687 7511 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11212 7510 7513 7512 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11211 11024 10687 7513 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11210 7511 7817 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11209 11024 7739 7510 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11208 7509 7512 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11207 11024 5846 5841 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11206 5846 10687 5625 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11205 5624 5850 5846 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11204 11024 10687 5850 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11203 5625 6877 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11202 11024 5842 5624 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11201 5841 5846 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11200 11024 6528 6530 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11199 6528 10687 6308 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11198 6307 6531 6528 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11197 11024 10687 6531 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11196 6308 7526 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11195 11024 6527 6307 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11194 6530 6528 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11193 11024 9729 7829 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11192 7827 7829 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11191 11024 8152 7827 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11190 7825 7827 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11189 11024 7827 7825 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11188 11024 4631 4594 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11187 4594 4954 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11186 11024 4955 4594 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11185 5131 4594 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11184 11024 7107 7108 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11183 7107 10687 6929 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11182 6928 7116 7107 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11181 11024 10687 7116 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11180 6929 8429 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11179 11024 7109 6928 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11178 7108 7107 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11177 9460 9552 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11176 10599 9609 9460 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11175 11024 9559 10599 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11174 11024 1890 1892 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11173 1892 1893 1891 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11172 3079 1891 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11171 11024 1574 1357 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11170 1357 1575 1572 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11169 2167 1572 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11168 1939 2140 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11167 4348 2138 1939 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11166 11024 10258 4348 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11165 9729 10395 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11164 9729 10701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11163 11024 10705 9729 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11162 11024 11072 9729 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11161 6179 7852 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11160 6179 7848 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11159 11024 6574 6179 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11158 5809 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11157 5809 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11156 11024 9020 5809 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11155 2537 3050 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11154 2763 2761 2537 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11153 11024 11042 2763 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11152 8163 9298 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11151 8629 8865 8163 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11150 11024 10197 8629 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11149 8710 8714 8712 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11148 11024 8713 8714 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11147 8711 9016 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11146 8712 8713 8711 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11145 11024 8709 8710 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11144 11024 8862 8254 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11143 8254 8262 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11142 8254 9298 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11141 11024 8865 8254 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11140 8817 8254 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11139 11024 3941 3947 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11138 3945 3938 3777 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11137 3777 3941 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11136 3777 3947 3945 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11135 11024 3942 3777 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11134 3942 3938 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_11133 11024 10709 10412 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11132 10412 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11131 11024 10708 10412 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11130 10408 10412 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11129 3975 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11128 11024 10031 3975 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11127 3974 3975 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11126 2171 4453 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11125 11024 2168 2171 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11124 2490 2171 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11123 1353 5599 1352 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11122 1352 1862 1533 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11121 1533 1529 1353 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11120 1353 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11119 11024 3967 1353 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11118 1528 1533 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11117 7020 7690 6919 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11116 6919 7019 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11115 11024 8903 7020 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11114 7046 7020 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11113 11024 10414 10404 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11112 10404 10705 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11111 11024 10708 10404 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11110 10399 10404 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11109 11024 4465 4362 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11108 4362 5297 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11107 11024 4361 4362 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11106 4369 4362 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11105 11024 5811 5560 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11104 5560 6241 5561 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11103 4381 5519 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11102 4535 5525 4381 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11101 11024 4553 4535 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11100 9325 9347 9326 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11099 9326 10366 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11098 11024 10017 9325 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11097 9323 9325 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_11096 738 739 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11095 733 740 734 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11094 11024 1005 733 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11093 740 741 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11092 11024 5262 741 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11091 11024 1008 739 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11090 736 740 738 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11089 737 741 736 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11088 11024 735 737 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11087 735 736 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11086 734 741 735 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11085 11024 734 1005 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11084 1005 734 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11083 8759 9421 8757 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11082 8758 9424 8759 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11081 8759 8756 8758 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11080 8757 9724 8759 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11079 8757 8760 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11078 11024 9073 8757 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11077 11024 10395 9721 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11076 9721 10710 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11075 11024 11072 9721 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11074 9716 9721 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11073 3790 4005 5009 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11072 3789 4003 3790 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11071 11024 4451 3789 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11070 11024 2213 2210 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11069 2210 2203 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11068 11024 3349 2210 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11067 5302 2210 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11066 9369 9372 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11065 9366 9373 9367 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11064 11024 9376 9366 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11063 9373 9374 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11062 11024 10638 9374 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11061 11024 9375 9372 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11060 9370 9373 9369 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11059 9371 9374 9370 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11058 11024 9368 9371 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11057 9368 9370 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11056 9367 9374 9368 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11055 11024 9367 9376 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11054 9376 9367 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11053 6226 6454 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11052 6223 6345 6452 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11051 11024 6468 6223 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11050 6345 6456 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11049 11024 10914 6456 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11048 11024 10257 6454 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11047 6344 6345 6226 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11046 6225 6456 6344 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11045 11024 6341 6225 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11044 6341 6344 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11043 6452 6456 6341 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11042 11024 6452 6468 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11041 6468 6452 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11040 10097 10228 10589 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11039 10096 10139 10097 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11038 11024 10232 10096 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11037 140 142 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11036 136 143 137 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11035 11024 341 136 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11034 143 144 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11033 11024 2673 144 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11032 11024 145 142 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11031 141 143 140 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11030 138 144 141 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11029 11024 139 138 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11028 139 141 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11027 137 144 139 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11026 11024 137 341 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11025 341 137 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11024 7557 7779 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11023 7555 7780 7773 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11022 11024 8407 7555 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11021 7780 7781 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11020 11024 8048 7781 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_11019 11024 7802 7779 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11018 7777 7780 7557 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11017 7556 7781 7777 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11016 11024 7774 7556 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11015 7774 7777 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11014 7773 7781 7774 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_11013 11024 7773 8407 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11012 8407 7773 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11011 7561 9552 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11010 8007 8644 7561 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11009 11024 8009 8007 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11008 8107 8713 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11007 8107 8709 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11006 11024 8092 8107 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11005 11024 8411 8179 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11004 8179 9033 8357 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_11003 8358 8357 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_11002 10847 10836 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11001 11024 10832 10847 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_11000 8184 10698 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10999 8453 10083 8184 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10998 11024 10708 8453 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10997 4970 4972 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10996 4965 4974 4966 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10995 11024 5191 4965 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10994 4974 4973 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10993 11024 5262 4973 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10992 11024 4969 4972 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10991 4971 4974 4970 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10990 4967 4973 4971 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10989 11024 4968 4967 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10988 4968 4971 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10987 4966 4973 4968 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10986 11024 4966 5191 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10985 5191 4966 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10984 4901 4902 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10983 4897 4904 4896 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10982 11024 8918 4897 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10981 4904 4903 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10980 11024 5083 4903 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10979 11024 5097 4902 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10978 4900 4904 4901 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10977 4898 4903 4900 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10976 11024 4899 4898 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10975 4899 4900 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10974 4896 4903 4899 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10973 11024 4896 8918 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10972 8918 4896 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10971 10544 10541 10543 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10970 10543 10542 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10969 11024 10774 10544 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10968 10540 10544 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10967 8029 8358 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10966 8341 8103 8029 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10965 11024 8206 8341 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10964 10769 11057 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10963 11059 11058 10769 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10962 11024 11054 11059 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10961 3976 3706 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10960 3976 6277 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10959 11024 5918 3976 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10958 220 4673 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10957 220 472 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10956 11024 1545 220 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10955 3690 4976 3692 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10954 3691 3958 3690 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10953 3689 3959 3691 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10952 11024 4979 3689 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10951 3688 3692 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10950 3045 3047 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10949 11024 7068 3045 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10948 3044 3045 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10947 3653 3893 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10946 11024 4410 3653 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10945 3658 3653 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10944 11024 9586 9577 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10943 9577 9572 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10942 11024 9579 9577 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10941 9571 9577 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10940 8657 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10939 8657 8661 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10938 11024 8922 8657 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10937 11024 8297 8657 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10936 8690 8708 8180 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10935 8180 8709 8690 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10934 11024 10606 8180 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10933 7079 7476 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10932 11024 7084 7079 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10931 7702 7079 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10930 8402 10704 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10929 8402 8403 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10928 11024 8437 8402 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10927 2728 7711 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10926 2728 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10925 11024 5898 2728 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10924 6592 10399 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10923 11024 9716 6592 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10922 452 219 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10921 452 482 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10920 11024 747 452 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10919 464 5837 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10918 464 472 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10917 11024 1545 464 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10916 3239 5181 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10915 11024 5842 3239 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10914 3236 3239 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10913 11024 5123 3619 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10912 3619 5119 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10911 11024 5131 3619 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10910 3617 3619 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10909 9613 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10908 9613 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10907 11024 9020 9613 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10906 11024 10963 9613 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10905 1881 8126 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10904 1881 5599 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10903 11024 7478 1881 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10902 11024 5809 1512 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10901 1512 4981 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10900 1512 7041 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10899 11024 1881 1512 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10898 2462 1512 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10897 815 10256 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10896 1044 1042 815 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10895 814 2472 1044 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10894 11024 2474 814 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10893 1041 1044 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10892 9926 10614 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10891 10006 10615 9926 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10890 11024 10024 10006 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10889 7048 7046 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10888 11024 7050 7048 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10887 7045 7048 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10886 6442 7022 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10885 11024 6798 6442 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10884 6440 6442 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10883 3783 3962 3963 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10882 3784 10596 3783 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10881 3782 3961 3784 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10880 11024 10595 3782 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10879 5168 3963 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10878 2548 2602 2797 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10877 2549 2801 2548 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10876 11024 2601 2549 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10875 2799 2797 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10874 11024 9421 8769 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10873 8769 9057 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10872 11024 9433 8769 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10871 8768 8769 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10870 818 4070 1059 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10869 819 8124 818 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10868 817 3092 819 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10867 11024 4066 817 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10866 1061 1059 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10865 2794 2792 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10864 11024 2791 2794 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10863 3403 2794 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10862 11024 3607 3609 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10861 3814 3606 3608 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10860 3608 3607 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10859 3608 3609 3814 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10858 11024 3605 3608 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10857 3605 3606 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10856 4883 6941 4882 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10855 11024 4880 4882 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10854 4882 9993 4883 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10853 4881 4883 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10852 11024 10073 8440 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10851 8440 10698 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10850 11024 11072 8440 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10849 8437 8440 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10848 9431 9433 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10847 11024 9716 9431 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10846 9750 9431 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10845 1880 4014 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10844 1879 6220 1880 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10843 1878 1881 1879 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10842 11024 3714 1878 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10841 2147 1879 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10840 8078 8623 8008 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10839 11024 8007 8008 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10838 8008 8834 8078 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10837 8262 8078 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10836 11024 7711 2504 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10835 2504 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10834 2504 7478 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10833 11024 9597 2504 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10832 2602 2504 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10831 11024 5583 5584 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10830 5584 6275 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10829 11024 7514 5584 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10828 6861 5584 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10827 1333 1433 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10826 1331 1435 1424 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10825 11024 1423 1331 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10824 1435 1434 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10823 11024 2673 1434 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10822 11024 1431 1433 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10821 1430 1435 1333 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10820 1332 1434 1430 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10819 11024 1427 1332 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10818 1427 1430 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10817 1424 1434 1427 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10816 11024 1424 1423 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10815 1423 1424 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10814 8035 8116 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10813 8033 8117 8114 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10812 11024 8122 8033 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10811 8117 8119 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10810 11024 10638 8119 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10809 11024 8120 8116 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10808 8115 8117 8035 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10807 8034 8119 8115 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10806 11024 8118 8034 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10805 8118 8115 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10804 8114 8119 8118 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10803 11024 8114 8122 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10802 8122 8114 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10801 10090 10568 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10800 10542 10564 10090 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10799 11024 10610 10542 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10798 6487 6506 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10797 11024 6496 6487 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10796 5063 7484 5579 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10795 5062 11042 5063 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10794 11024 6493 5062 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10793 5562 7749 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10792 6259 6246 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10791 8654 8090 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10790 10568 10567 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10789 10583 9922 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10788 10890 10213 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10787 5783 7041 5620 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10786 11024 10619 5620 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10785 5620 7042 5783 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10784 5782 5783 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10783 1255 1257 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10782 1251 1259 1252 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10781 11024 1826 1251 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10780 1259 1258 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10779 11024 2446 1258 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10778 11024 1437 1257 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10777 1256 1259 1255 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10776 1254 1258 1256 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10775 11024 1253 1254 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10774 1253 1256 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10773 1252 1258 1253 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10772 11024 1252 1826 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10771 1826 1252 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10770 11024 6859 5836 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10769 10687 5836 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10768 11024 5836 10687 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10767 11024 5836 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10766 11024 5836 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10765 11024 6859 6860 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10764 8733 6860 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10763 11024 6860 8733 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10762 11024 6860 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10761 11024 6860 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10760 11024 6255 6256 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10759 6859 6256 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10758 11024 6256 6859 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10757 11024 6256 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10756 11024 6256 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10755 11024 7667 7563 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10754 7563 9379 7669 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10753 8094 7669 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10752 10230 10606 10098 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10751 10098 10608 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10750 11024 10854 10230 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10749 10228 10230 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10748 3768 10604 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10747 6379 8091 3768 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10746 11024 9304 6379 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10745 2138 3413 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10744 11024 2473 2138 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10743 5541 8623 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10742 6116 8617 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10741 5093 8839 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10740 4975 7085 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10739 6797 7652 6795 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10738 6796 8090 6797 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10737 6797 8635 6796 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10736 6795 8636 6797 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10735 6795 8297 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10734 11024 8633 6795 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10733 1821 2412 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10732 5748 2413 1821 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10731 11024 4325 5748 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10730 4500 4277 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10729 11024 4272 4500 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10728 1806 1804 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10727 1806 2998 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10726 11024 1805 1806 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10725 6940 7158 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10724 6938 7157 7149 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10723 11024 7147 6938 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10722 7157 7160 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10721 11024 8048 7160 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10720 11024 7154 7158 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10719 7156 7157 6940 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10718 6939 7160 7156 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10717 11024 7153 6939 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10716 7153 7156 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10715 7149 7160 7153 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10714 11024 7149 7147 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10713 7147 7149 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10712 8767 9429 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10711 11024 9732 8767 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10710 11054 10687 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10709 11024 11042 11054 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10708 8752 9046 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10707 8751 8750 8752 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10706 11024 8749 8751 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10705 10258 3379 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10704 11024 6275 10258 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10703 2416 8014 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10702 11024 2415 2416 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10701 3006 5535 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10700 11024 3007 3006 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10699 3654 3006 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10698 3219 2996 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10697 11024 4410 3219 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10696 8784 8880 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10695 8782 8879 8870 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10694 11024 8869 8782 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10693 8879 8881 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10692 11024 10914 8881 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10691 11024 8878 8880 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10690 8876 8879 8784 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10689 8783 8881 8876 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10688 11024 8873 8783 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10687 8873 8876 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10686 8870 8881 8873 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10685 11024 8870 8869 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10684 8869 8870 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10683 10248 10963 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10682 10248 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10681 11024 10027 10248 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10680 7619 7618 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10679 11024 7615 7619 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10678 8081 7619 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10677 11024 9987 4014 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10676 11024 2481 1888 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10675 4014 1888 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10674 730 1495 732 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10673 732 1494 731 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10672 731 729 732 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10671 730 984 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10670 11024 1489 730 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10669 732 1005 730 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10668 2692 731 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10667 8017 8651 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10666 11024 8089 8017 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10665 4291 5153 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10664 11024 5718 4291 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10663 7688 7684 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10662 11024 7685 7688 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10661 10564 7688 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10660 7695 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10659 7695 7711 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10658 11024 7721 7695 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10657 11024 8725 7695 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10656 9680 9433 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10655 9680 9421 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10654 11024 10697 9680 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10653 11024 9716 9680 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10652 9073 10073 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10651 11024 10708 9073 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10650 8024 8318 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10649 8101 8316 8024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10648 11024 8954 8101 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10647 8816 5755 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10646 11024 5748 8816 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10645 2383 2962 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10644 2384 5124 2383 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10643 11024 3615 2384 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10642 3830 4959 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10641 3830 4508 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10640 11024 4939 3830 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10639 11024 4954 3830 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10638 3915 4306 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10637 3914 4312 3759 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10636 3759 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10635 11024 3906 3762 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10634 3762 3905 3760 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10633 3760 3915 3914 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10632 3914 4306 3761 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10631 3761 4322 3762 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10630 11024 4929 3906 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10629 3917 3914 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10628 3666 4306 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10627 3670 3664 3665 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10626 3665 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10625 11024 3667 3671 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10624 3671 3668 3669 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10623 3669 3666 3670 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10622 3670 4306 3672 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10621 3672 4320 3671 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10620 11024 4929 3667 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_10619 3938 3670 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10618 11024 8659 8660 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10617 8660 8657 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10616 11024 8658 8660 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10615 8913 8660 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10614 6299 8713 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10613 6475 6473 6299 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10612 6298 10018 6475 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10611 11024 6476 6298 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10610 7468 6475 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10609 11024 9663 10701 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10608 9663 10684 9452 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10607 9451 9666 9663 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10606 11024 10684 9666 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10605 9452 10257 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10604 11024 9947 9451 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10603 10701 9663 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10602 11024 7670 7462 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10601 7462 7673 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10600 7667 7459 7462 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10599 7461 7460 7667 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10598 7462 7463 7461 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10597 1936 7678 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10596 2093 5898 1936 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10595 11024 2736 2093 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10594 8154 8155 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10593 11024 11066 8154 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10592 8460 8154 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10591 5840 10687 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10590 11024 5837 5840 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10589 6524 5840 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10588 7534 8453 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10587 7534 9421 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10586 11024 10399 7534 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10585 11024 9716 7534 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10584 10518 10575 10574 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10583 10519 10604 10518 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10582 10517 10892 10519 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10581 11024 10888 10517 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10580 10832 10574 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10579 3716 6251 3717 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_10578 3715 3714 3716 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_10577 11024 7465 3715 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_10576 3717 3718 11024 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_10575 7999 8065 9633 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10574 11024 9987 8065 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10573 7998 8072 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10572 9633 9987 7998 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10571 11024 8064 7999 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10570 4956 10018 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10569 4956 5809 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10568 11024 6221 4956 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10567 11024 6220 4956 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10566 11024 7711 4565 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10565 4565 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10564 4565 8921 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10563 11024 8617 4565 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10562 4567 4565 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10561 6120 6778 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10560 6119 6205 6120 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10559 11024 6206 6119 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10558 8454 9421 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10557 11024 8453 8454 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10556 8756 8454 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10555 6763 7605 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10554 11024 6959 6763 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10553 6762 6763 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10552 211 217 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10551 210 213 211 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10550 209 449 210 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10549 11024 451 209 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10548 1495 210 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10547 11024 6241 5801 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10546 11024 6476 5800 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10545 5801 5800 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10544 7537 7824 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10543 11024 10027 7537 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10542 7536 7537 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10541 4334 4333 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10540 11024 4439 4334 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10539 4342 4334 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10538 1349 1501 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10537 1503 2090 1349 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10536 1348 2098 1503 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10535 11024 1500 1348 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10534 2459 1503 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10533 8837 8839 8774 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10532 11024 8835 8774 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10531 8774 8834 8837 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10530 8833 8837 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10529 8615 8617 8614 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10528 8614 8834 8615 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10527 11024 8616 8614 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10526 11024 10701 9094 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10525 9094 10709 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10524 9094 9405 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10523 11024 10708 9094 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10522 9087 9094 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10521 11024 7484 6958 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10520 7415 8122 6910 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10519 6910 7484 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10518 6910 6958 7415 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10517 11024 6954 6910 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10516 6954 8122 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10515 11024 8047 5576 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10514 5576 10915 5577 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10513 11024 9309 3737 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10512 3737 9314 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10511 3737 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10510 11024 5293 3737 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10509 4048 3737 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10508 4304 5159 4303 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10507 4303 6127 4304 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10506 11024 6213 4303 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10505 716 718 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10504 713 719 712 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10503 11024 711 713 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10502 719 720 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10501 11024 2446 720 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10500 11024 722 718 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10499 717 719 716 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10498 715 720 717 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10497 11024 714 715 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10496 714 717 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10495 712 720 714 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10494 11024 712 711 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10493 711 712 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10492 8719 8721 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10491 8715 8722 8716 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10490 11024 9007 8715 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10489 8722 8723 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10488 11024 10638 8723 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10487 11024 9006 8721 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10486 8720 8722 8719 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10485 8718 8723 8720 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10484 11024 8717 8718 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10483 8717 8720 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10482 8716 8723 8717 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10481 11024 8716 9007 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10480 9007 8716 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10479 8006 8075 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10478 8004 8076 8071 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10477 11024 8072 8004 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10476 8076 8077 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10475 11024 10914 8077 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10474 11024 10231 8075 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10473 8074 8076 8006 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10472 8005 8077 8074 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10471 11024 8073 8005 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10470 8073 8074 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10469 8071 8077 8073 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10468 11024 8071 8072 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10467 8072 8071 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10466 10602 10605 10865 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10465 10601 10599 10602 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10464 11024 10600 10601 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10463 11024 6175 5602 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10462 5604 5603 5606 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10461 5605 5931 5604 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10460 5602 5601 5605 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10459 132 133 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10458 128 134 127 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10457 11024 692 128 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10456 134 135 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10455 11024 2673 135 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10454 11024 329 133 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10453 130 134 132 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10452 131 135 130 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10451 11024 129 131 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10450 129 130 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10449 127 135 129 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10448 11024 127 692 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10447 692 127 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10446 9331 9932 10142 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10445 9330 9332 9331 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10444 11024 9329 9330 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10443 1812 2413 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10442 2000 2412 1812 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10441 11024 10888 2000 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10440 11024 5610 5028 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10439 5030 5040 5032 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10438 5031 5029 5030 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10437 5028 5286 5031 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10436 5060 5214 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10435 5216 5565 5060 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10434 11024 5220 5216 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10433 6871 6874 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10432 6868 6875 6869 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10431 11024 6867 6868 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10430 6875 6876 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10429 11024 8048 6876 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10428 11024 7144 6874 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10427 6872 6875 6871 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10426 6873 6876 6872 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10425 11024 6870 6873 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10424 6870 6872 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10423 6869 6876 6870 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10422 11024 6869 6867 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10421 6867 6869 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10420 2379 2380 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10419 2374 2381 2375 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10418 11024 7484 2374 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10417 2381 2382 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10416 11024 5083 2382 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10415 11024 3158 2380 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10414 2378 2381 2379 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10413 2377 2382 2378 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10412 11024 2376 2377 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10411 2376 2378 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10410 2375 2382 2376 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10409 11024 2375 7484 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10408 7484 2375 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10407 9985 9984 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10406 11024 9987 9985 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10405 10877 10589 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10404 11024 10590 10877 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10403 8475 8059 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10402 11024 9107 8475 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10401 10137 9996 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10400 11024 9997 10137 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10399 4926 4955 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10398 4926 4631 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10397 11024 4954 4926 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10396 1973 4915 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10395 1973 5131 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10394 11024 3817 1973 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10393 2414 2413 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10392 2989 2412 2414 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10391 11024 2688 2989 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10390 7550 7665 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10389 7548 7664 7657 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10388 11024 7655 7548 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10387 7664 7666 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10386 11024 10914 7666 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10385 11024 8030 7665 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10384 7662 7664 7550 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10383 7549 7666 7662 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10382 11024 7661 7549 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10381 7661 7662 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10380 7657 7666 7661 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10379 11024 7657 7655 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10378 7655 7657 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10377 7059 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10376 7059 5801 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10375 11024 5919 7059 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10374 11024 9308 7059 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10373 8443 9057 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10372 8443 9702 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10371 11024 9080 8443 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10370 8092 7721 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10369 8092 9020 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10368 11024 5911 8092 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10367 5286 5283 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10366 11024 5891 5286 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10365 3053 3704 3051 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10364 3051 3967 3052 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10363 3052 9308 3053 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10362 3053 3969 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10361 11024 5599 3053 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10360 3050 3052 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10359 3193 4617 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10358 3193 5123 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10357 11024 5119 3193 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10356 3676 3677 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10355 3684 3675 3676 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10354 11024 3952 3684 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10353 6754 6757 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10352 6750 6756 6751 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10351 11024 8699 6750 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10350 6756 6758 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10349 11024 10914 6758 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10348 11024 6963 6757 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10347 6755 6756 6754 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10346 6753 6758 6755 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10345 11024 6752 6753 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10344 6752 6755 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10343 6751 6758 6752 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10342 11024 6751 8699 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10341 8699 6751 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10340 10223 10222 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10339 11024 10225 10223 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10338 10565 10223 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10337 6862 6863 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10336 6862 6861 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10335 11024 6864 6862 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10334 7817 7835 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10333 7817 8754 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10332 11024 8054 7817 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10331 8754 10704 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10330 8754 9066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10329 11024 9095 8754 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10328 5000 4998 4999 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10327 4999 9002 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10326 11024 5001 5000 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10325 4997 5000 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10324 11024 5194 5190 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10323 5190 5202 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10322 11024 5771 5190 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10321 5185 5190 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10320 3620 4508 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10319 11024 4939 3620 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10318 3618 3620 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10317 5123 10312 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10316 5123 5728 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10315 11024 5727 5123 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10314 11024 866 867 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10313 866 9379 779 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10312 778 868 866 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10311 11024 9379 868 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10310 779 4489 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10309 11024 8885 778 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10308 867 866 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10307 11024 6369 6370 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10306 6369 9379 6288 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10305 6287 6371 6369 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10304 11024 9379 6371 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10303 6288 6376 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10302 11024 8642 6287 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10301 6370 6369 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10300 11024 5492 5487 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10299 5492 9379 5491 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10298 5489 5493 5492 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10297 11024 9379 5493 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10296 5491 5490 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10295 11024 5488 5489 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10294 5487 5492 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10293 11024 4991 4669 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10292 4669 4665 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10291 11024 4666 4669 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10290 7457 4669 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10289 7529 8052 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10288 7529 8155 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10287 11024 10399 7529 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10286 2475 2474 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10285 4347 2472 2475 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10284 11024 4327 4347 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10283 460 6261 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10282 460 472 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10281 11024 1545 460 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10280 11024 5498 5494 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10279 5498 9379 5497 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10278 5495 5499 5498 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10277 11024 9379 5499 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10276 5497 5496 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10275 11024 9304 5495 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10274 5494 5498 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10273 8938 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10272 8938 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10271 11024 9560 8938 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10270 11024 8305 8938 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10269 10111 10273 10323 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10268 11024 10774 10273 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10267 10110 10652 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10266 10323 10774 10110 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10265 11024 10789 10111 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10264 7404 8064 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10263 11024 10197 7404 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10262 10525 10839 10588 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10261 10524 10604 10525 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10260 10523 10892 10524 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10259 11024 10888 10523 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10258 10590 10588 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10257 6911 10604 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10256 6959 8091 6911 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10255 11024 8699 6959 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10254 5069 6493 5267 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10253 5068 7484 5069 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10252 11024 11042 5068 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10251 5269 5267 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10250 8620 8840 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10249 11024 10197 8620 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10248 6216 6796 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10247 11024 6817 6216 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10246 6130 6216 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10245 11024 10698 10069 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10244 10069 10083 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10243 11024 10700 10069 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10242 10689 10069 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10241 5089 5667 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10240 11024 5091 5089 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10239 5086 5089 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10238 5051 6116 5104 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10237 5049 10604 5051 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10236 5050 10892 5049 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10235 11024 10888 5050 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10234 5103 5104 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10233 9464 9620 10366 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10232 11024 10774 9620 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10231 9465 10268 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10230 10366 10774 9465 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10229 11024 10620 9464 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10228 5180 7041 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10227 11024 7042 5180 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10226 5177 5180 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10225 216 482 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10224 11024 219 216 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10223 215 216 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10222 2518 5753 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10221 2679 3000 2518 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10220 11024 3236 2679 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10219 11024 10073 9070 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10218 9070 10709 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10217 11024 10686 9070 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10216 9066 9070 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10215 11024 6760 6761 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10214 6761 6766 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10213 11024 7655 6761 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10212 6759 6761 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10211 11024 3735 2502 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10210 2502 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10209 11024 5293 2502 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10208 2500 2502 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10207 11024 10698 8755 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10206 8755 9405 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10205 11024 10708 8755 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10204 9057 8755 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10203 156 155 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10202 151 157 150 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10201 11024 348 151 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10200 157 158 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10199 11024 2673 158 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10198 11024 347 155 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10197 154 157 156 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10196 152 158 154 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10195 11024 153 152 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10194 153 154 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10193 150 158 153 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10192 11024 150 348 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10191 348 150 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10190 11024 9922 9986 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10189 11024 10774 9274 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10188 9986 9274 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10187 11024 5600 5234 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10186 5234 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10185 11024 6277 5234 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10184 5229 5234 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10183 11024 9314 1303 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10182 1303 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10181 1303 5600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10180 11024 9308 1303 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10179 1573 1303 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10178 7448 8869 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10177 6109 8848 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10176 6455 9287 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10175 1928 2680 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10174 3213 2681 1928 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10173 11024 2688 3213 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10172 3877 4290 3771 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10171 3771 4288 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10170 11024 4285 3877 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10169 3875 3877 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10168 7504 7506 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10167 7500 7508 7501 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10166 11024 7739 7500 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10165 7508 7507 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10164 11024 8048 7507 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10163 11024 7509 7506 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10162 7505 7508 7504 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10161 7502 7507 7505 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10160 11024 7503 7502 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10159 7503 7505 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10158 7501 7507 7503 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10157 11024 7501 7739 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10156 7739 7501 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10155 8080 7425 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10154 8080 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10153 11024 10027 8080 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10152 6995 6997 6916 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10151 6916 7004 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10150 11024 6994 6995 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10149 6993 6995 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_10148 4452 4996 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10147 11024 5580 4452 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10146 6863 7117 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10145 8995 9007 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10144 5851 7147 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10143 5564 6527 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10142 7460 7652 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10141 7444 8082 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10140 1913 2049 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10139 1911 2048 2039 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10138 11024 2038 1911 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10137 2048 2050 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10136 11024 2446 2050 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10135 11024 2047 2049 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10134 2046 2048 1913 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10133 1912 2050 2046 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10132 11024 2043 1912 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10131 2043 2046 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10130 2039 2050 2043 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10129 11024 2039 2038 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10128 2038 2039 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10127 5628 5861 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10126 5626 5860 5853 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10125 11024 6545 5626 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10124 5860 5862 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10123 11024 8048 5862 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10122 11024 6543 5861 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10121 5858 5860 5628 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10120 5627 5862 5858 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10119 11024 5857 5627 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10118 5857 5858 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10117 5853 5862 5857 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10116 11024 5853 6545 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10115 6545 5853 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10114 10731 10875 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10113 10729 10874 10868 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10112 11024 10880 10729 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10111 10874 10876 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10110 11024 10914 10876 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10109 11024 10879 10875 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10108 10873 10874 10731 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10107 10730 10876 10873 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10106 11024 10869 10730 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10105 10869 10873 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10104 10868 10876 10869 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10103 11024 10868 10880 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10102 10880 10868 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10101 8648 7450 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10100 8648 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10099 11024 10027 8648 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10098 2472 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10097 11024 8126 2472 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10096 8893 8642 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10095 11024 2209 1897 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10094 1900 1898 2791 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10093 1901 1899 1900 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10092 1897 2208 1901 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10091 3425 6130 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10090 11024 3003 3425 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10089 9918 9993 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10088 9984 10200 9918 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10087 11024 9991 9984 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10086 1301 4981 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10085 11024 1302 1301 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10084 1296 1292 1297 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10083 1294 1293 1296 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10082 1295 1528 1294 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10081 11024 1291 1295 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_10080 1500 1297 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10079 7165 7533 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10078 11024 7828 7165 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10077 8390 8128 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10076 11024 8402 8390 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10075 8128 8121 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10074 11024 8388 8128 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10073 10699 10698 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10072 11024 10708 10699 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10071 10128 10414 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10070 10419 11075 10128 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10069 11024 10686 10419 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10068 11024 4070 820 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10067 821 8124 3735 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10066 822 3092 821 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10065 820 4066 822 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10064 4953 5181 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10063 11024 7109 4953 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10062 4952 4953 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10061 7544 7629 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10060 7542 7628 7622 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10059 11024 8082 7542 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10058 7628 7630 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10057 11024 10914 7630 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_10056 11024 7634 7629 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10055 7627 7628 7544 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10054 7543 7630 7627 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10053 11024 7623 7543 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10052 7623 7627 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10051 7622 7630 7623 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_10050 11024 7622 8082 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10049 8082 7622 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10048 8659 8305 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10047 8659 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10046 11024 10027 8659 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10045 7499 7770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10044 11024 7740 7499 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_10043 7498 7499 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10042 11024 10046 9946 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10041 10046 11019 9949 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10040 9948 9950 10046 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10039 11024 11019 9950 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10038 9949 10257 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10037 11024 9947 9948 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10036 9946 10046 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10035 11024 10050 10292 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10034 10050 11019 9952 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10033 9951 9953 10050 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10032 11024 11019 9953 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10031 9952 10231 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10030 11024 10289 9951 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10029 10292 10050 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10028 11024 10294 10668 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10027 10294 11019 10115 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10026 10114 10296 10294 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10025 11024 11019 10296 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10024 10115 10312 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10023 11024 10662 10114 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10022 10668 10294 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10021 11024 10061 10059 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10020 10061 11019 9963 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10019 9962 9964 10061 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10018 11024 11019 9964 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10017 9963 10024 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10016 11024 10054 9962 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10015 10059 10061 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10014 11024 10347 10348 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10013 10347 11019 10123 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10012 10122 10354 10347 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10011 11024 11019 10354 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10010 10123 10594 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10009 11024 10350 10122 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10008 10348 10347 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10007 11024 9364 9419 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10006 9364 10684 9363 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10005 9361 9365 9364 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10004 11024 10684 9365 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10003 9363 9362 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10002 11024 9639 9361 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_10001 9419 9364 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_10000 4915 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09999 4915 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09998 11024 6277 4915 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09997 11024 8839 4915 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09996 11024 11014 11036 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09995 11014 11019 10762 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09994 10761 11023 11014 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09993 11024 11019 11023 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09992 10762 11018 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09991 11024 11028 10761 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09990 11036 11014 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09989 11024 10679 11006 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09988 10679 11019 10537 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09987 10536 10678 10679 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09986 11024 11019 10678 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09985 10537 10680 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09984 11024 10999 10536 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09983 11006 10679 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09982 7522 9046 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09981 7521 8050 7522 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09980 11024 7520 7521 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09979 5933 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09978 5933 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09977 11024 6278 5933 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09976 11024 7514 5933 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09975 9924 10614 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09974 9997 10615 9924 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09973 11024 10231 9997 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09972 2646 2657 1924 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09971 1924 2984 2646 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09970 11024 3632 1924 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09969 4939 8921 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09968 4939 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09967 11024 5719 4939 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09966 11024 8617 4939 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09965 11024 7615 6460 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09964 6460 7465 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09963 11024 8713 6460 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09962 6457 6460 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09961 11024 3033 3034 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09960 3034 10018 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09959 3034 7042 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09958 11024 6251 3034 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09957 5727 3034 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09956 11024 7756 7752 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09955 7756 8733 7553 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09954 7554 7758 7756 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09953 11024 8733 7758 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09952 7553 8042 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09951 11024 7749 7554 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09950 7752 7756 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09949 11024 10334 10414 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09948 10334 10684 10121 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09947 10120 10340 10334 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09946 11024 10684 10340 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09945 10121 10680 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09944 11024 10999 10120 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09943 10414 10334 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09942 11024 2462 2463 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09941 2463 3044 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09940 2463 2727 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09939 11024 3036 2463 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09938 5728 2463 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09937 8634 9296 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09936 8864 9297 8634 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09935 11024 10197 8864 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09934 9474 9979 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09933 10075 9750 9474 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09932 11024 9747 10075 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09931 8429 8426 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09930 8429 8431 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09929 11024 8430 8429 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09928 11024 8443 8429 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09927 11024 7006 6444 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09926 6449 9610 6295 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09925 6295 7006 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09924 6295 6444 6449 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09923 11024 6445 6295 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09922 6445 9610 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09921 9278 10269 9277 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09920 9277 10256 9276 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09919 9276 10258 9278 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09918 9278 9486 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09917 11024 9503 9278 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09916 9275 9276 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09915 6112 6109 6193 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09914 6110 10604 6112 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09913 6111 10892 6110 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09912 11024 10888 6111 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09911 6108 6193 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09910 1825 2680 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09909 1824 2681 1825 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09908 11024 10888 1824 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09907 3377 2491 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09906 3377 2492 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09905 11024 2493 3377 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09904 11024 2490 3377 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09903 1823 2681 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09902 1822 2680 1823 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09901 11024 4325 1822 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09900 11024 1210 1205 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09899 4489 3611 1204 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09898 1204 1210 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09897 1204 1205 4489 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09896 11024 1203 1204 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09895 1203 3611 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09894 10094 10890 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09893 10218 10564 10094 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09892 11024 10215 10218 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09891 10257 9362 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09890 5598 6896 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09889 11024 6574 5598 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09888 5601 5598 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09887 1838 7701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09886 11024 1844 1838 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09885 1837 1838 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09884 5637 9605 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09883 5743 7437 5637 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09882 11024 9323 5743 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09881 9294 9293 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09880 9292 9290 9294 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09879 11024 9291 9292 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09878 11024 10698 8153 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09877 8153 11076 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09876 11024 10700 8153 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09875 8155 8153 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09874 1045 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09873 11024 7514 1045 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09872 1529 1045 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09871 11024 3064 3067 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09870 3067 3065 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09869 11024 3066 3067 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09868 3076 3067 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09867 8031 8725 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09866 8675 8106 8031 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09865 11024 8107 8675 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09864 11024 6592 6596 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09863 6596 6591 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09862 11024 6908 6596 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09861 6590 6596 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09860 2430 2692 2431 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09859 2431 2691 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09858 11024 2688 2430 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09857 3004 2430 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09856 2522 3008 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09855 4305 3009 2522 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09854 11024 2688 4305 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09853 191 192 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09852 186 193 187 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09851 11024 724 186 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09850 193 194 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09849 11024 2446 194 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09848 11024 195 192 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09847 190 193 191 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09846 189 194 190 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09845 11024 188 189 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09844 188 190 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09843 187 194 188 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09842 11024 187 724 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09841 724 187 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09840 11024 753 473 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09839 473 750 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09838 473 1871 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09837 11024 8713 473 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09836 472 473 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09835 794 1495 795 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09834 795 1494 958 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09833 958 959 795 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09832 794 951 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09831 11024 1489 794 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09830 795 1245 794 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09829 2681 958 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09828 1347 1496 1346 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09827 1857 1493 1347 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09826 1347 1494 1857 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09825 1346 1495 1347 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09824 1346 1490 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09823 11024 1489 1346 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09822 2638 3611 2512 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09821 2512 2968 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09820 11024 2637 2638 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09819 2636 2638 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09818 249 251 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09817 245 252 246 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09816 11024 244 245 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09815 252 253 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09814 11024 5262 253 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09813 11024 2373 251 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09812 250 252 249 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09811 248 253 250 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09810 11024 247 248 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09809 247 250 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09808 246 253 247 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09807 11024 246 244 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09806 244 246 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09805 9440 9497 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09804 9438 9499 9491 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09803 11024 9489 9438 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09802 9499 9500 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09801 11024 10914 9500 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09800 11024 10312 9497 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09799 9498 9499 9440 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09798 9439 9500 9498 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09797 11024 9493 9439 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09796 9493 9498 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09795 9491 9500 9493 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09794 11024 9491 9489 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09793 9489 9491 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09792 10738 10899 10918 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09791 10737 10900 10738 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09790 11024 10897 10737 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09789 9462 9605 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09788 10034 9609 9462 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09787 11024 10017 10034 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09786 11024 5901 1894 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09785 1894 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09784 1894 5719 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09783 11024 7678 1894 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09782 1893 1894 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09781 4985 5564 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09780 4984 4983 4985 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09779 11024 4986 4984 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09778 810 1027 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09777 808 1026 1020 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09776 11024 1496 808 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09775 1026 1028 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09774 11024 5262 1028 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09773 11024 1025 1027 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09772 1022 1026 810 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09771 809 1028 1022 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09770 11024 1023 809 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09769 1023 1022 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09768 1020 1028 1023 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09767 11024 1020 1496 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09766 1496 1020 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09765 8811 9043 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09764 8809 9042 9035 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09763 11024 9033 8809 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09762 9042 9045 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09761 11024 11051 9045 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09760 11024 9047 9043 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09759 9041 9042 8811 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09758 8810 9045 9041 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09757 11024 9039 8810 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09756 9039 9041 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09755 9035 9045 9039 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09754 11024 9035 9033 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09753 9033 9035 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09752 5623 5831 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09751 5621 5833 5824 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09750 11024 6819 5621 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09749 5833 5834 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09748 11024 8048 5834 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09747 11024 5829 5831 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09746 5832 5833 5623 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09745 5622 5834 5832 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09744 11024 5826 5622 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09743 5826 5832 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09742 5824 5834 5826 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09741 11024 5824 6819 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09740 6819 5824 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09739 269 5488 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09738 11024 5488 300 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09737 293 2957 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09736 11024 293 269 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09735 269 300 297 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09734 297 2957 269 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09733 1958 297 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09732 11024 297 1958 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09731 11024 9433 8764 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09730 8764 9746 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09729 8762 9750 8764 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09728 8763 9081 8762 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09727 8764 9087 8763 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09726 10917 10865 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09725 11024 10861 10917 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09724 10265 10606 10109 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09723 10109 10608 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09722 11024 10924 10265 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09721 10899 10265 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09720 3154 7690 3102 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09719 3102 3804 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09718 11024 7403 3154 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09717 3152 3154 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09716 6281 7176 6172 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09715 6172 6286 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09714 11024 6280 6281 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09713 6171 6281 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09712 4960 5771 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09711 4960 5194 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09710 11024 5202 4960 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09709 5124 4955 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09708 5124 4631 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09707 11024 4952 5124 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09706 11024 5131 2966 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09705 2966 2965 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09704 2964 3615 2966 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09703 2963 2962 2964 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09702 2966 5124 2963 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09701 1199 1200 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09700 1194 1201 1195 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09699 11024 2957 1194 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09698 1201 1202 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09697 11024 5083 1202 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09696 11024 2956 1200 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09695 1198 1201 1199 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09694 1197 1202 1198 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09693 11024 1196 1197 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09692 1196 1198 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09691 1195 1202 1196 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09690 11024 1195 2957 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09689 2957 1195 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09688 9743 11072 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09687 9743 10078 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09686 11024 10701 9743 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09685 10951 10142 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09684 11024 10618 10951 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09683 5610 6177 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09682 11024 6180 5610 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09681 3072 2782 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09680 3072 3349 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09679 11024 3081 3072 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09678 6828 6829 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09677 6823 6831 6822 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09676 11024 8691 6823 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09675 6831 6830 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09674 11024 10638 6830 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09673 11024 6827 6829 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09672 6826 6831 6828 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09671 6825 6830 6826 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09670 11024 6824 6825 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09669 6824 6826 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09668 6822 6830 6824 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09667 11024 6822 8691 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09666 8691 6822 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09665 6772 6774 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09664 6768 6775 6769 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09663 11024 9313 6768 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09662 6775 6776 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09661 11024 10914 6776 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09660 11024 6777 6774 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09659 6773 6775 6772 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09658 6771 6776 6773 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09657 11024 6770 6771 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09656 6770 6773 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09655 6769 6776 6770 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09654 11024 6769 9313 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09653 9313 6769 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09652 7558 9305 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09651 8616 8644 7558 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09650 11024 7585 8616 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09649 7064 7059 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09648 11024 7058 7064 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09647 7061 7064 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09646 2460 2464 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09645 10959 2459 2460 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09644 11024 9987 10959 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09643 8822 10547 8773 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09642 8773 10555 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09641 11024 10915 8822 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09640 8821 8822 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09639 4977 4984 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09638 11024 8691 4977 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09637 4976 4977 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09636 1809 2004 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09635 1991 2006 1809 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09634 11024 2688 1991 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09633 7014 7063 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09632 11024 9541 7014 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09631 7012 7014 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09630 11024 6781 6777 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09629 6781 9379 6779 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09628 6780 6782 6781 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09627 11024 9379 6782 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09626 6779 6778 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09625 11024 9313 6780 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09624 6777 6781 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09623 11024 6962 6963 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09622 6962 9379 6913 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09621 6912 6973 6962 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09620 11024 9379 6973 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09619 6913 6967 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09618 11024 8699 6912 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09617 6963 6962 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09616 8613 9298 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09615 8613 8262 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09614 11024 8862 8613 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09613 11024 8865 8613 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09612 8054 8152 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09611 8054 9421 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09610 11024 9433 8054 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09609 1035 1862 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09608 1035 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09607 11024 7514 1035 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09606 11024 3032 2368 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09605 2368 3029 2449 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09604 2450 2449 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09603 11024 6212 6427 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09602 6212 9379 6124 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09601 6125 6126 6212 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09600 11024 9379 6126 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09599 6124 6205 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09598 11024 8930 6125 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09597 6427 6212 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09596 11024 10248 10254 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09595 10254 10247 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09594 11024 10249 10254 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09593 10611 10254 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09592 11024 8833 5653 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09591 5653 8824 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09590 11024 8817 5653 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09589 6942 5653 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09588 11024 9298 8631 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09587 8631 8862 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09586 8631 9296 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09585 11024 9297 8631 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09584 9290 8631 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09583 11024 9033 8685 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09582 11024 8930 8209 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09581 8685 8209 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09580 10070 9975 9973 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09579 11024 10687 9973 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09578 9973 10692 10070 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09577 9972 10070 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09576 9105 9104 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09575 11024 10080 9105 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09574 9103 9105 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09573 7835 9433 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09572 7835 8458 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09571 11024 8059 7835 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09570 11024 2481 1356 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09569 1356 10915 1560 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09568 3714 1560 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09567 11024 11042 3793 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09566 3793 7484 4011 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09565 4010 4011 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09564 11024 8124 3091 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09563 3090 3091 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09562 11024 3092 3090 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09561 3410 3090 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09560 11024 3090 3410 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09559 8906 9316 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09558 11024 10197 8906 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09557 2729 10269 2528 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09556 2528 10256 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09555 11024 2728 2729 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09554 3035 2729 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09553 1922 5124 1921 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09552 1921 2962 1967 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09551 1967 3615 1922 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09550 1922 2965 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09549 11024 5131 1922 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09548 1964 1967 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09547 11024 5719 5110 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09546 5110 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09545 5110 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09544 11024 8623 5110 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09543 5105 5110 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09542 8789 10614 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09541 8915 10615 8789 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09540 11024 10995 8915 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09539 8150 8758 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09538 11024 8151 8150 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09537 8053 8150 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09536 10736 10890 10893 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09535 10734 10891 10736 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09534 10735 10892 10734 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09533 11024 10888 10735 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09532 10919 10893 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09531 6173 6574 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09530 6173 8770 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09529 11024 9107 6173 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09528 11024 7852 6173 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09527 9486 9505 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09526 11024 10774 9486 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09525 11024 8709 2739 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09524 2739 2572 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09523 2739 4012 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09522 11024 2578 2739 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09521 3036 2739 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09520 9307 9305 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09519 10139 9609 9307 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09518 11024 9306 10139 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09517 8098 8096 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09516 11024 8097 8098 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09515 8021 8098 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09514 10621 10620 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09513 11024 10774 10621 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09512 8157 10083 8061 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09511 8061 10710 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09510 11024 11072 8157 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09509 8060 8157 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09508 6588 6898 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09507 11024 6590 6588 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09506 6586 6588 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09505 5323 5321 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09504 11024 5934 5323 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09503 5320 5323 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09502 3038 10018 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09501 11024 3057 3038 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09500 3306 3038 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09499 6128 6214 6129 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09498 6129 6215 6128 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09497 11024 6213 6129 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09496 11024 10701 9423 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09495 9423 10078 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09494 9423 10083 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09493 11024 11072 9423 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09492 9429 9423 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09491 1814 7701 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09490 11024 1813 1814 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09489 2413 1814 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09488 3184 5105 3110 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09487 3110 3630 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09486 11024 4553 3184 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09485 3183 3184 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09484 10178 10179 10085 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09483 11024 10176 10085 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09482 10085 10184 10178 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09481 10177 10178 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09480 11024 8661 4695 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09479 4695 6276 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09478 11024 5898 4695 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09477 5275 4695 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09476 11024 4465 4722 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09475 4722 5032 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09474 4722 5297 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09473 11024 4467 4722 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09472 4723 4722 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09471 11024 5202 4326 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09470 4326 5771 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09469 11024 8092 4326 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09468 4325 4326 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09467 11024 9987 1963 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09466 1961 1963 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09465 11024 8617 1961 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09464 8310 1961 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09463 11024 1961 8310 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09462 8807 9382 9016 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09461 8806 9667 8807 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09460 11024 9033 8806 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09459 11024 9020 4990 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09458 4990 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09457 11024 7478 4990 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09456 5226 4990 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09455 11024 4720 4358 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09454 4358 4359 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09453 11024 4710 4358 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09452 4364 4358 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09451 11024 5898 3089 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09450 3089 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09449 3089 7711 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09448 11024 7721 3089 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09447 3088 3089 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09446 11024 7204 7196 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09445 7196 7536 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09444 7196 7837 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09443 11024 7201 7196 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09442 7190 7196 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09441 11024 8472 6899 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09440 6899 6904 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09439 6899 7190 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09438 11024 6900 6899 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09437 6898 6899 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09436 791 926 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09435 789 928 915 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09434 11024 916 789 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09433 928 929 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09432 11024 2673 929 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09431 11024 925 926 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09430 917 928 791 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09429 790 929 917 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09428 11024 920 790 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09427 920 917 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09426 915 929 920 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09425 11024 915 916 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09424 916 915 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09423 5572 5573 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09422 5567 5574 5568 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09421 11024 5842 5567 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09420 5574 5575 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09419 11024 8048 5575 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09418 11024 5841 5573 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09417 5571 5574 5572 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09416 5570 5575 5571 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09415 11024 5569 5570 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09414 5569 5571 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09413 5568 5575 5569 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09412 11024 5568 5842 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09411 5842 5568 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09410 9305 8885 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09409 6760 7484 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09408 9552 9304 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09407 9333 8918 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09406 9566 8699 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09405 9605 9313 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09404 11024 3084 3083 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09403 3083 3082 4361 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09402 11024 6435 5057 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09401 5057 5528 5151 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09400 5150 5151 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09399 4296 4948 4297 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09398 4297 4298 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09397 11024 4295 4296 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09396 4539 4296 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09395 800 978 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09394 798 980 969 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09393 11024 1456 798 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09392 980 981 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09391 11024 2446 981 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09390 11024 1260 978 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09389 970 980 800 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09388 799 981 970 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09387 11024 974 799 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09386 974 970 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09385 969 981 974 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09384 11024 969 1456 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09383 1456 969 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09382 7618 7611 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09381 7618 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09380 11024 9582 7618 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09379 6146 6241 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09378 6473 6233 6146 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09377 11024 7474 6473 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09376 8026 8092 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09375 11024 8713 8026 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09374 10235 10595 10099 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09373 10099 10596 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09372 11024 10231 10235 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09371 10232 10235 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09370 3071 3066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09369 3071 3064 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09368 11024 3065 3071 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09367 11024 1575 1359 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09366 1360 1583 3077 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09365 1358 1573 1360 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09364 1359 1574 1358 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09363 4451 3993 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09362 11024 3994 4451 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09361 6765 6992 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09360 6766 8122 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09359 9610 8930 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09358 6803 8297 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09357 11024 3079 2543 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09356 2544 2590 3402 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09355 2542 3355 2544 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09354 2543 2589 2542 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09353 3610 3607 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09352 11024 2973 3610 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09351 10745 10941 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09350 10743 10940 10935 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09349 11024 10945 10743 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09348 10940 10942 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09347 11024 11051 10942 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09346 11024 10944 10941 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09345 10939 10940 10745 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09344 10744 10942 10939 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09343 11024 10934 10744 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09342 10934 10939 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09341 10935 10942 10934 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09340 11024 10935 10945 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09339 10945 10935 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09338 11024 1861 1863 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09337 1863 1862 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09336 2094 3040 1863 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09335 1860 7678 2094 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09334 1863 5898 1860 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09333 8120 8394 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09332 11024 8123 8120 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09331 6228 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09330 6228 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09329 11024 10029 6228 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09328 6243 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09327 6243 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09326 11024 8661 6243 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09325 2140 5600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09324 11024 6277 2140 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09323 3705 5898 3701 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09322 3701 5599 3702 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09321 3702 4653 3705 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09320 3705 3703 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09319 11024 3704 3705 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09318 10595 3702 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09317 2670 6431 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09316 11024 3213 2670 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09315 3198 2670 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09314 7547 7645 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09313 7545 7644 7638 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09312 11024 7652 7545 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09311 7644 7646 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09310 11024 10914 7646 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09309 11024 8019 7645 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09308 7643 7644 7547 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09307 7546 7646 7643 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09306 11024 7639 7546 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09305 7639 7643 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09304 7638 7646 7639 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09303 11024 7638 7652 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09302 7652 7638 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09301 8298 8938 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09300 11024 10018 8298 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09299 8658 8298 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09298 7599 7600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09297 11024 10018 7599 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09296 8070 7599 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09295 11024 10988 10989 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09294 10988 11019 10757 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09293 10756 10998 10988 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09292 11024 11019 10998 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09291 10757 10995 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09290 11024 10990 10756 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09289 10989 10988 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09288 8123 8121 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09287 11024 8122 8123 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09286 3033 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09285 3033 2133 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09284 11024 9020 3033 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09283 3057 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09282 3057 2133 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09281 11024 9314 3057 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09280 2419 2418 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09279 8089 2417 2419 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09278 11024 4325 8089 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09277 3178 5123 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09276 11024 5119 3178 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09275 3175 3178 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09274 11024 7086 7089 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09273 7086 10687 6923 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09272 6924 7094 7086 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09271 11024 10687 7094 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09270 6923 7784 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09269 11024 7085 6924 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09268 7089 7086 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09267 6255 10028 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09266 6255 7721 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09265 11024 7514 6255 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09264 11024 10197 6255 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09263 11024 10020 9315 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09262 11024 10774 9317 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09261 9315 9317 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09260 11024 2481 1307 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09259 1306 1307 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09258 11024 9987 1306 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09257 1308 1306 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09256 11024 1306 1308 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09255 11024 10673 10705 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09254 10673 10684 10533 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09253 10532 10674 10673 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09252 11024 10684 10674 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09251 10533 10908 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09250 11024 10675 10532 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09249 10705 10673 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09248 11024 10676 11075 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09247 10676 10684 10535 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09246 10534 10677 10676 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09245 11024 10684 10677 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09244 10535 10995 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09243 11024 10990 10534 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09242 11075 10676 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09241 11024 10318 10378 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09240 10318 10684 10119 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09239 10118 10324 10318 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09238 11024 10684 10324 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09237 10119 10323 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09236 11024 10332 10118 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09235 10378 10318 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09234 11024 2753 2536 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09233 2536 3723 2759 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09232 2761 2759 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09231 11024 5240 1869 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09230 1869 1867 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09229 11024 1868 1869 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09228 1866 1869 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09227 3627 3630 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09226 3626 5105 3627 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09225 11024 4553 3626 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09224 11024 5131 4278 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09223 4278 4281 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09222 4277 4279 4278 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09221 4276 5124 4277 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09220 4278 4275 4276 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09219 3656 3664 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_09218 3662 3654 3655 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09217 3655 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09216 11024 3657 3660 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09215 3660 3658 3659 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09214 3659 3656 3662 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09213 3662 3664 3661 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09212 3661 4587 3660 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09211 11024 4929 3657 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_09210 4940 3662 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09209 11024 9489 8621 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09208 11024 10197 8622 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09207 8621 8622 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09206 11024 10358 10395 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09205 10358 10684 10125 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09204 10124 10367 10358 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09203 11024 10684 10367 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09202 10125 10366 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09201 11024 11013 10124 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09200 10395 10358 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09199 11024 10682 11076 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09198 10682 10684 10539 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09197 10538 10683 10682 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09196 11024 10684 10683 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09195 10539 11018 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09194 11024 11028 10538 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09193 11076 10682 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09192 11024 6277 5526 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09191 5526 10031 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09190 5526 8643 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09189 11024 9287 5526 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09188 5525 5526 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09187 3637 3871 3111 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09186 3111 4535 3637 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09185 11024 3632 3111 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09184 3251 3664 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_09183 3255 3242 3122 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09182 3122 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09181 11024 3243 3125 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09180 3125 3246 3123 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09179 3123 3251 3255 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09178 3255 3664 3124 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09177 3124 4304 3125 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09176 11024 4929 3243 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_09175 3890 3255 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09174 4884 6749 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09173 4885 6942 4884 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09172 11024 5162 4885 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09171 11024 11063 10072 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09170 10072 10074 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09169 11024 10075 10072 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09168 9975 10072 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09167 11024 3032 2453 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09166 2451 2453 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09165 11024 2454 2451 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09164 2452 2451 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09163 11024 2451 2452 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09162 10521 10583 10581 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09161 10522 10604 10521 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09160 10520 10892 10522 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09159 11024 10888 10520 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09158 10582 10581 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09157 8639 8848 8637 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09156 8638 10213 8639 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09155 8639 8635 8638 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09154 8637 8636 8639 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09153 8637 8699 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09152 11024 8633 8637 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09151 10198 10559 10088 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09150 10088 10571 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09149 11024 10197 10198 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09148 10558 10198 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09147 3121 3884 3120 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09146 3120 3242 3232 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09145 3232 3230 3121 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09144 3121 5842 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09143 11024 5181 3121 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09142 3647 3232 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09141 11024 3814 3816 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09140 5496 4501 3769 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09139 3769 3814 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09138 3769 3816 5496 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09137 11024 3810 3769 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09136 3810 4501 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09135 11024 8869 8866 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09134 11024 10774 8632 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09133 8866 8632 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09132 3836 3833 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09131 11024 5103 3836 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09130 3832 3836 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09129 1858 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09128 11024 9560 1858 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09127 3040 1858 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09126 6503 6493 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09125 7084 7739 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09124 9379 10774 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09123 6499 8047 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09122 8983 9382 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09121 5274 5269 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09120 11024 5607 5274 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09119 5271 5274 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09118 11024 2962 1207 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09117 1207 1964 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09116 1801 2637 1207 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09115 1206 1796 1801 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09114 1207 3611 1206 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09113 8311 8313 8175 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09112 11024 8310 8175 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09111 8175 8309 8311 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_09110 8312 8311 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09109 8646 9333 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09108 8645 8644 8646 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09107 11024 8647 8645 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09106 3060 4014 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09105 3058 7042 3060 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09104 3059 6220 3058 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09103 11024 3714 3059 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09102 3066 3058 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09101 4360 4359 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09100 11024 4710 4360 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09099 4467 4360 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09098 6477 6476 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09097 6490 6241 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09096 8408 8407 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09095 8708 9033 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09094 8731 8409 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09093 11024 215 212 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09092 212 220 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09091 212 745 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09090 11024 460 212 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09089 1494 212 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09088 8166 8839 8165 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09087 8277 10800 8166 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09086 8166 8635 8277 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09085 8165 8636 8166 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09084 8165 8642 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09083 11024 8633 8165 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09082 10557 10619 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09081 10555 10564 10557 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09080 11024 10554 10555 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09079 11024 10915 3805 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09078 3803 3805 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09077 11024 8090 3803 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09076 4880 3803 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09075 11024 3803 4880 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09074 2457 10269 2458 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09073 2458 10256 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09072 11024 2578 2457 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09071 2456 2457 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_09070 3700 3967 3697 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09069 3697 3974 3699 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09068 3699 5599 3700 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09067 3700 3698 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09066 11024 9308 3700 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09065 10596 3699 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09064 11024 9314 2178 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09063 2178 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09062 2178 8922 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09061 11024 7678 2178 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09060 2177 2178 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09059 11024 11042 5064 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09058 5064 7484 5253 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09057 11024 8922 5879 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09056 5879 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09055 5879 8126 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09054 11024 9597 5879 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09053 5878 5879 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09052 5142 1806 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09051 11024 1807 5142 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_09050 226 228 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09049 222 229 223 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09048 11024 6241 222 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09047 229 230 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09046 11024 5262 230 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09045 11024 231 228 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09044 227 229 226 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09043 225 230 227 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09042 11024 224 225 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09041 224 227 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09040 223 230 224 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09039 11024 223 6241 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09038 6241 223 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09037 9931 10023 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09036 9929 10025 10019 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09035 11024 10020 9929 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09034 10025 10026 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09033 11024 10914 10026 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09032 11024 10024 10023 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09031 10022 10025 9931 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09030 9930 10026 10022 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09029 11024 10021 9930 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09028 10021 10022 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09027 10019 10026 10021 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09026 11024 10019 10020 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09025 10020 10019 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09024 8610 8839 8160 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09023 8160 8834 8610 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09022 11024 8835 8160 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09021 9935 10033 10147 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09020 9934 10034 9935 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09019 11024 10032 9934 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09018 11024 4344 4345 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09017 4343 4345 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09016 11024 4342 4343 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09015 4465 4343 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09014 11024 4343 4465 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09013 11024 10137 10091 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09012 10091 10214 10205 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_09011 10551 10205 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_09010 702 703 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09009 697 704 699 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09008 11024 1245 697 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09007 704 705 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09006 11024 2673 705 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_09005 11024 1244 703 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09004 701 704 702 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09003 698 705 701 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09002 11024 700 698 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09001 700 701 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_09000 699 705 700 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08999 11024 699 1245 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08998 1245 699 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08997 10171 10542 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08996 11024 10541 10171 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08995 8020 8094 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08994 8019 8095 8020 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08993 11024 8093 8019 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08992 10548 10550 10515 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08991 11024 10773 10515 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08990 10515 10559 10548 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08989 10796 10548 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08988 9342 9343 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08987 9337 9345 9336 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08986 11024 9335 9337 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08985 9345 9344 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08984 11024 10914 9344 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08983 11024 9341 9343 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08982 9339 9345 9342 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08981 9340 9344 9339 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08980 11024 9338 9340 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08979 9338 9339 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08978 9336 9344 9338 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08977 11024 9336 9335 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08976 9335 9336 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08975 10718 10810 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08974 10716 10811 10803 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08973 11024 10800 10716 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08972 10811 10812 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08971 11024 10914 10812 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08970 11024 10808 10810 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08969 10807 10811 10718 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08968 10717 10812 10807 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08967 11024 10804 10717 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08966 10804 10807 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08965 10803 10812 10804 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08964 11024 10803 10800 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08963 10800 10803 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08962 10977 10918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08961 11024 10919 10977 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08960 9943 10043 10158 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08959 9942 10044 9943 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08958 11024 10042 9942 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08957 9061 9080 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08956 11024 9057 9061 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08955 2487 5911 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08954 2487 3735 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08953 11024 6278 2487 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08952 7067 7069 6922 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08951 11024 9362 6922 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08950 6922 7068 7067 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08949 7063 7067 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08948 2657 4617 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08947 2657 3817 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08946 11024 4915 2657 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08945 3182 3193 3109 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08944 11024 3632 3109 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08943 3109 3626 3182 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08942 3179 3182 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08941 8793 8951 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08940 8791 8950 8943 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08939 11024 8954 8791 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08938 8950 8952 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08937 11024 10914 8952 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08936 11024 8949 8951 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08935 8948 8950 8793 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08934 8792 8952 8948 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08933 11024 8942 8792 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08932 8942 8948 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08931 8943 8952 8942 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08930 11024 8943 8954 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08929 8954 8943 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08928 6242 6506 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08927 11024 6496 6242 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08926 6150 6242 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08925 8292 8291 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08924 11024 8290 8292 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08923 8682 8292 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08922 9976 10700 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08921 9976 10073 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08920 11024 10701 9976 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08919 9692 10700 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08918 9692 10698 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08917 11024 10083 9692 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08916 8788 10269 8787 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08915 8787 10256 8908 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08914 8908 10258 8788 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08913 8788 8906 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08912 11024 9315 8788 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08911 8903 8908 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08910 4700 3734 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08909 4700 3735 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08908 11024 6278 4700 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08907 4013 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08906 4013 3735 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08905 11024 6278 4013 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08904 10007 10005 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08903 11024 10006 10007 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08902 10554 10007 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08901 2982 4617 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08900 2982 4508 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08899 11024 4939 2982 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08898 11024 6214 5137 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08897 5137 6215 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08896 11024 5131 5137 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08895 5132 5137 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08894 11024 3934 3928 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08893 3934 4318 3764 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08892 3763 3937 3934 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08891 11024 4318 3937 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08890 3764 4617 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08889 11024 4553 3763 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08888 3928 3934 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08887 6211 6429 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08886 6208 6333 6425 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08885 11024 8930 6208 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08884 6333 6430 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08883 11024 10914 6430 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08882 11024 6427 6429 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08881 6332 6333 6211 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08880 6209 6430 6332 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08879 11024 6331 6209 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08878 6331 6332 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08877 6425 6430 6331 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08876 11024 6425 8930 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08875 8930 6425 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08874 10201 10564 10089 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08873 10089 10568 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08872 11024 10610 10201 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08871 10200 10201 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08870 7684 6251 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08869 7684 6457 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08868 11024 6232 7684 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08867 11024 6230 7684 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08866 9746 9743 9473 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_08865 9472 9980 9746 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_08864 11024 9976 9472 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_08863 9473 9760 11024 11024 sg13_lv_pmos L=0.13U W=3.47U AS=0.8328P AD=0.8328P PS=7.42U PD=7.42U 
Mtr_08862 9760 10708 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08861 9760 10709 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08860 11024 11076 9760 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08859 9468 9692 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08858 9682 9680 9468 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08857 11024 9678 9682 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08856 10702 10686 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08855 10702 10378 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08854 11024 11075 10702 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08853 7201 9747 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08852 7201 10704 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08851 11024 9716 7201 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08850 5556 8092 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08849 5556 5202 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08848 11024 5771 5556 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08847 4508 10231 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08846 4508 5728 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08845 11024 5727 4508 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08844 5539 8921 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08843 5539 9309 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08842 11024 7711 5539 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08841 11024 7652 5539 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08840 9971 10686 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08839 9971 10073 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08838 11024 10709 9971 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08837 10892 5214 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08836 10892 5207 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08835 11024 9609 10892 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08834 11024 8092 10892 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08833 4183 6277 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08832 4183 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08831 11024 10031 4183 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08830 11024 8643 4183 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08829 11024 10909 10913 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08828 11024 10915 10916 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08827 10913 10916 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08826 11024 6201 6197 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08825 6967 6200 6115 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08824 6115 6201 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08823 6115 6197 6967 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08822 11024 6198 6115 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08821 6198 6200 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08820 6135 7448 6217 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08819 6133 10604 6135 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08818 6134 10892 6133 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08817 11024 6132 6134 11024 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_08816 6131 6217 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08815 7176 8052 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08814 7176 8453 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08813 11024 9433 7176 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08812 11024 9716 7176 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08811 6280 6275 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08810 6280 6278 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08809 11024 6276 6280 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08808 11024 6277 6280 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08807 9938 10789 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08806 11024 10774 9938 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08805 6821 8318 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08804 6820 8316 6821 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08803 11024 6819 6820 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08802 11024 6992 6420 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08801 6420 8122 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08800 11024 7655 6420 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08799 6784 6420 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08798 8018 10604 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08797 8097 8091 8018 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08796 11024 9313 8097 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08795 4399 4708 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08794 4710 6560 4399 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08793 11024 5293 4710 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08792 10896 10901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08791 11024 10915 10896 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08790 3999 4666 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08789 11024 6243 3999 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08788 4003 3999 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08787 11024 4543 4538 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08786 6778 4539 4382 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08785 4382 4543 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08784 4382 4538 6778 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08783 11024 4540 4382 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08782 4540 4539 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08781 11024 11026 10685 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08780 10708 10685 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08779 11024 10685 10708 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08778 11024 10685 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08777 11024 10685 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08776 11024 11026 10681 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08775 10700 10681 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08774 11024 10681 10700 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08773 11024 10681 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08772 11024 10681 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08771 11024 11026 11027 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08770 11072 11027 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08769 11024 11027 11072 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08768 11024 11027 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08767 11024 11027 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08766 11024 11026 10688 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08765 10686 10688 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08764 11024 10688 10686 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08763 11024 10688 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08762 11024 10688 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08761 11024 7766 7768 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08760 11026 7768 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08759 11024 7768 11026 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08758 11024 7768 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08757 11024 7768 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08756 11024 4701 4704 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08755 4704 5873 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08754 11024 4700 4704 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08753 5014 4704 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08752 11024 5293 3796 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08751 3796 4038 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08750 4354 6278 3796 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08749 3795 4030 4354 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08748 3796 4031 3795 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08747 758 1881 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08746 11024 1556 758 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08745 759 758 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08744 2682 2681 2519 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08743 2519 2680 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08742 11024 2688 2682 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08741 2997 2682 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08740 11024 1314 768 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08739 7514 768 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08738 11024 768 7514 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08737 11024 768 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08736 11024 768 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08735 11024 1314 1315 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08734 8126 1315 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08733 11024 1315 8126 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08732 11024 1315 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08731 11024 1315 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08730 11024 773 772 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08729 1314 772 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08728 11024 772 1314 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08727 11024 772 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08726 11024 772 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08725 11024 508 504 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08724 7721 504 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08723 11024 504 7721 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08722 11024 504 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08721 11024 504 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08720 11024 508 506 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08719 7478 506 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08718 11024 506 7478 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08717 11024 506 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08716 11024 506 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08715 11024 510 509 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08714 508 509 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08713 11024 509 508 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08712 11024 509 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08711 11024 509 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08710 11024 8662 8663 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08709 10027 8663 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08708 11024 8663 10027 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08707 11024 8663 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08706 11024 8663 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08705 11024 8662 8656 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08704 9582 8656 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08703 11024 8656 9582 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08702 11024 8656 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08701 11024 8656 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08700 11024 8100 8099 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08699 8662 8099 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08698 11024 8099 8662 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08697 11024 8099 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08696 11024 8099 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08695 7472 7690 7473 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08694 7473 7475 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08693 11024 9624 7472 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08692 7471 7472 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08691 11024 9609 4978 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08690 4978 5214 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08689 11024 8092 4978 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08688 7690 4978 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08687 11024 1884 1885 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08686 1885 1886 2168 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08685 11024 7540 6903 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08684 6903 6901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08683 11024 6902 6903 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08682 6900 6903 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08681 11024 2158 2152 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08680 2152 2776 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08679 11024 2147 2152 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08678 4333 2152 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08677 11024 5757 5762 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08676 5762 5756 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08675 11024 6141 5762 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08674 5755 5762 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08673 11024 8297 3952 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08672 11024 10915 3954 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08671 3952 3954 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08670 11024 6402 6396 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08669 6401 6394 6290 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08668 6290 6402 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08667 6290 6396 6401 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08666 11024 6397 6290 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08665 6397 6394 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08664 11024 5600 1304 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08663 1304 8661 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08662 1304 6275 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08661 11024 5293 1304 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08660 1884 1304 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08659 1275 1277 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08658 1271 1278 1272 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08657 11024 1493 1271 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08656 1278 1279 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08655 11024 5262 1279 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08654 11024 1280 1277 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08653 1276 1278 1275 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08652 1273 1279 1276 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08651 11024 1274 1273 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08650 1274 1276 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08649 1272 1279 1274 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08648 11024 1272 1493 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08647 1493 1272 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08646 8037 8388 8038 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08645 8036 8411 8037 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08644 11024 9033 8036 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08643 10607 10606 10609 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08642 10609 10608 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08641 11024 10880 10607 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08640 10605 10607 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08639 11024 5600 1607 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08638 1607 5901 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08637 1607 7711 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08636 11024 5599 1607 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08635 1899 1607 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08634 11024 2212 1951 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08633 1951 2211 2213 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08632 4401 5023 4478 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08631 4400 5037 4401 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08630 11024 4476 4400 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08629 6257 6522 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08628 6253 6357 6520 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08627 11024 6527 6253 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08626 6357 6523 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08625 11024 8048 6523 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08624 11024 6530 6522 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08623 6356 6357 6257 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08622 6254 6523 6356 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08621 11024 6353 6254 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08620 6353 6356 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08619 6520 6523 6353 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08618 11024 6520 6527 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08617 6527 6520 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08616 6303 6493 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08615 6496 8713 6303 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08614 11024 8709 6496 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08613 5829 6152 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08612 11024 6151 5829 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08611 8430 10399 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08610 11024 8746 8430 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08609 8426 10399 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08608 11024 9080 8426 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08607 10636 10637 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08606 10632 10639 10631 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08605 11024 10924 10632 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08604 10639 10640 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08603 11024 10638 10640 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08602 11024 10923 10637 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08601 10635 10639 10636 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08600 10633 10640 10635 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08599 11024 10634 10633 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08598 10634 10635 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08597 10631 10640 10634 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08596 11024 10631 10924 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08595 10924 10631 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08594 10095 10614 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08593 10225 10615 10095 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08592 11024 11018 10225 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08591 7058 7466 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08590 7058 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08589 11024 10027 7058 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08588 6151 6518 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08587 11024 6819 6151 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08586 9029 11066 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08585 11024 10689 9029 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08584 7042 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08583 7042 2133 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08582 11024 9020 7042 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08581 6220 5918 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08580 6220 2133 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08579 11024 9314 6220 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08578 11024 3726 3730 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08577 3731 3728 4058 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08576 3729 4037 3731 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08575 3730 4023 3729 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08574 449 4995 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08573 11024 1545 449 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08572 213 482 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08571 11024 219 213 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08570 11024 4324 4553 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08569 4324 5181 4245 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08568 4246 4247 4324 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08567 11024 5181 4247 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08566 4245 4628 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08565 11024 4975 4246 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08564 4553 4324 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08563 11024 4634 6213 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08562 4634 5181 4394 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08561 4393 4635 4634 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08560 11024 5181 4635 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08559 4394 4640 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08558 11024 7085 4393 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08557 6213 4634 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08556 11024 4615 4617 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08555 4615 5181 4391 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08554 4390 4621 4615 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08553 11024 5181 4621 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08552 4391 4628 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08551 11024 5562 4390 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08550 4617 4615 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08549 7600 7601 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08548 7600 10036 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08547 11024 9582 7600 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08546 7526 7529 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08545 11024 7805 7526 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08544 2099 9308 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08543 2099 5600 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08542 11024 9020 2099 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08541 1995 6978 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08540 11024 1991 1995 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08539 1993 1995 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08538 3616 4926 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08537 11024 3822 3616 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08536 3615 3616 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08535 4920 4936 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08534 4922 5150 4918 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08533 4918 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08532 11024 4917 4923 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08531 4923 4919 4921 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08530 4921 4920 4922 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08529 4922 4936 4924 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08528 4924 6128 4923 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08527 11024 4929 4917 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08526 5518 4922 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08525 4933 4936 11024 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08524 4934 5527 4931 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08523 4931 4929 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08522 11024 4930 4937 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08521 4937 4932 4935 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08520 4935 4933 4934 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08519 4934 4936 4938 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08518 4938 5148 4937 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08517 11024 4929 4930 11024 sg13_lv_pmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08516 5681 4934 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08515 10721 10819 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08514 10719 10822 10813 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08513 11024 10825 10719 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08512 10822 10823 11024 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08511 11024 10914 10823 11024 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08510 11024 10824 10819 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08509 10820 10822 10721 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08508 10720 10823 10820 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08507 11024 10815 10720 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08506 10815 10820 11024 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08505 10813 10823 10815 11024 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08504 11024 10813 10825 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08503 10825 10813 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08502 7449 7448 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08501 9296 7463 7449 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08500 11024 7447 9296 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08499 3049 3057 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08498 11024 6220 3049 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08497 3331 3049 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08496 10076 10408 9978 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08495 9978 11067 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08494 11024 10399 10076 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08493 9977 10076 11024 11024 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_08492 11024 8962 9355 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08491 8962 9379 8797 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08490 8796 8969 8962 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08489 11024 9379 8969 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08488 8797 9095 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08487 11024 9350 8796 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08486 9355 8962 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08485 11024 9377 9375 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08484 9377 9379 9380 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08483 9378 9381 9377 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08482 11024 9379 9381 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08481 9380 9958 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08480 11024 9376 9378 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08479 9375 9377 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08478 11024 9004 9006 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08477 9004 9379 8805 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08476 8804 9015 9004 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08475 11024 9379 9015 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08474 8805 9051 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08473 11024 9007 8804 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08472 9006 9004 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08471 11024 233 231 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08470 233 6241 234 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08469 232 235 233 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08468 11024 6241 235 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08467 234 241 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08466 11024 6243 232 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08465 231 233 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08464 11024 9413 9412 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08463 9413 10684 9415 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08462 9414 9416 9413 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08461 11024 10684 9416 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08460 9415 9509 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08459 11024 9701 9414 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08458 9412 9413 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08457 11024 10062 10710 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08456 10062 10684 9965 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08455 9966 9967 10062 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08454 11024 10684 9967 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08453 9965 10594 11024 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08452 11024 10350 9966 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08451 10710 10062 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08450 6221 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08449 6221 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08448 11024 7711 6221 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08447 7041 9597 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08446 7041 5919 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08445 11024 7514 7041 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08444 9303 9306 11024 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08443 11024 10018 9303 11024 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08442 9533 9303 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08441 2640 2982 2513 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08440 2513 3625 2640 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08439 11024 3632 2513 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08438 3633 3871 3634 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08437 11024 3632 3634 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08436 3634 4535 3633 11024 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08435 3849 3633 11024 11024 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_08434 9892 10008 9891 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08433 9894 10011 10010 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08432 11074 10009 9893 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08431 10222 10010 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08430 878 1268 877 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08429 11074 875 876 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08428 11074 1268 883 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08427 881 4910 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08426 882 880 881 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08425 879 901 878 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08424 876 875 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08423 323 1268 321 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08422 11074 325 320 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08421 11074 1268 326 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08420 327 4905 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08419 322 328 327 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08418 324 338 323 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08417 320 325 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08416 4663 5898 4664 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08415 4662 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08414 4665 7711 4663 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08413 9212 10684 9211 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08412 11074 9408 9405 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08411 11074 10684 9216 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08410 9214 9612 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08409 9215 9410 9214 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08408 9213 9688 9212 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08407 9405 9408 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08406 9694 10684 9693 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08405 11074 9698 10083 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08404 11074 10684 9699 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08403 9696 10024 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08402 9697 9700 9696 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08401 9695 10054 9694 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_08400 10083 9698 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08399 2160 7721 2159 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08398 2161 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08397 2156 8126 2155 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08396 2158 9597 2157 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08395 1626 2384 1625 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08394 1627 1973 1800 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08393 11074 2403 1628 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08392 1802 1800 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08391 5097 5100 5096 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08390 5096 5094 5097 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08389 11074 5503 5095 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08388 11074 9743 9078 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08387 9076 9732 9077 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08386 9074 9077 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08385 8384 9419 8383 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08384 8383 10036 8384 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08383 11074 8970 8383 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08382 8395 8384 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08381 11074 10689 10490 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08380 10491 11066 10690 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08379 10691 10690 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08378 5509 5541 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08377 11074 10604 5509 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08376 5509 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08375 11074 10888 5509 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08374 5504 5509 5346 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08373 3862 6277 3867 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08372 3863 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08371 3865 10028 3864 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08370 3860 3866 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08369 3866 3861 3865 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08368 11074 7031 7034 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08367 7032 7471 7035 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08366 7033 7035 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08365 2 116 6376 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08364 11074 2636 3 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08363 5 1793 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08362 6376 115 4 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08361 6 1793 116 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08360 115 2636 1 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08359 10175 10540 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08358 10174 10171 10173 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08357 11074 10172 10174 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08356 10186 10174 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08355 11074 8126 3343 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08354 3344 10031 3345 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08353 3967 3345 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08352 11074 7721 1125 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08351 1126 9020 1286 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08350 1861 1286 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08349 6439 9333 6438 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08348 6438 7437 6439 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08347 11074 9321 6438 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08346 6437 6439 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08345 1040 756 606 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08344 606 1042 1040 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08343 11074 1873 605 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08342 6500 6497 6501 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08341 6501 6498 6500 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08340 11074 6499 6501 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08339 6847 6500 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08338 7788 8430 7792 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08337 7793 8431 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08336 7790 8443 7789 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08335 7786 7791 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08334 7791 7787 7790 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08333 7050 10891 7052 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08332 7052 8091 7050 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08331 11074 8918 7051 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08330 11074 4183 4044 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08329 4045 6173 4046 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08328 4043 4046 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08327 6646 9560 6645 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08326 6647 9309 6794 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08325 11074 8921 6648 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08324 8091 6794 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08323 11074 10700 7851 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08322 7853 10083 7854 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08321 7852 7854 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08320 4221 4701 4220 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08319 4224 4354 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08318 4223 5873 4222 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08317 5313 4355 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08316 4355 4219 4223 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08315 2756 6277 2755 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08314 2758 5600 2757 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08313 11074 3413 2754 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08312 2753 2757 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08311 91 753 90 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08310 92 750 221 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08309 11074 1871 93 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08308 219 221 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08307 6009 6236 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08306 6008 6237 6235 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08305 6006 6239 6234 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08304 11074 6476 6006 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08303 11074 8048 6239 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08302 6237 6239 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08301 11074 6478 6236 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08300 6235 6239 6009 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08299 6007 6235 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08298 11074 6238 6010 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08297 6234 6237 6238 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08296 6476 6234 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08295 11074 6234 6476 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08294 7679 10031 7681 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08293 7682 9314 7683 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08292 11074 7678 7680 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08291 10615 7683 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08290 1563 2741 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08289 11074 3714 1563 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08288 1563 2578 1561 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08287 1562 4014 1563 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08286 8570 9419 8569 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08285 8571 10073 8747 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08284 11074 10708 8572 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08283 8746 8747 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08282 2942 7721 2941 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08281 2943 5898 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08280 2940 7514 2939 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08279 3086 3087 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08278 3087 2938 2940 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08277 4458 5583 4457 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08276 4461 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08275 4460 9560 4459 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08274 5008 4690 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_08273 4690 4456 4460 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08272 3170 3617 3171 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08271 3171 3188 3170 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08270 11074 3606 3171 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08269 3612 3170 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08268 11074 8424 8088 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08267 8016 8088 7884 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08266 11074 8088 8016 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08265 11074 8088 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08264 11024 8088 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08263 11074 8145 8087 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08262 8015 8087 7883 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08261 11074 8087 8015 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08260 11074 8087 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08259 11024 8087 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08258 11074 8424 2775 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08257 5262 2775 2774 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08256 11074 2775 5262 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08255 11074 2775 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08254 11024 2775 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08253 11074 8424 2771 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08252 2773 2771 2772 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08251 11074 2771 2773 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08250 11074 2771 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08249 11024 2771 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08248 11074 8424 2484 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08247 2483 2484 2308 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08246 11074 2484 2483 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08245 11074 2484 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08244 11024 2484 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08243 11074 8145 2482 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08242 2481 2482 2307 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08241 11074 2482 2481 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08240 11074 2482 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08239 11024 2482 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08238 11074 8424 2676 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08237 5083 2676 2675 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08236 11074 2676 5083 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08235 11074 2676 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08234 11024 2676 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08233 11074 8424 2674 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08232 2673 2674 2672 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08231 11074 2674 2673 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08230 11074 2674 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08229 11024 2674 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08228 11074 8424 2422 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08227 2446 2422 2268 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08226 11074 2422 2446 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08225 11074 2422 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08224 11024 2422 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08223 11074 8145 2421 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08222 2420 2421 2267 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08221 11074 2421 2420 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08220 11074 2421 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08219 11024 2421 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08218 8463 9750 8462 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08217 8464 9107 8463 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08216 8465 9087 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08215 8459 8463 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08214 11074 9103 8461 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08213 8464 8460 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08212 11074 244 243 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08211 108 243 242 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08210 11074 2373 108 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08209 241 242 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08208 11074 242 241 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08207 4359 2796 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08206 11074 2799 4359 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08205 523 678 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08204 522 677 676 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08203 520 679 672 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08202 11074 901 520 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08201 11074 2673 679 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08200 677 679 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08199 11074 876 678 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08198 676 679 523 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08197 521 676 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08196 11074 673 524 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08195 672 677 673 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08194 901 672 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08193 11074 672 901 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08192 9522 9524 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08191 9517 9523 9521 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08190 9515 9525 9516 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08189 11074 9514 9515 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08188 11074 10914 9525 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08187 9523 9525 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08186 11074 10594 9524 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08185 9521 9525 9522 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08184 9518 9521 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08183 11074 9520 9519 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08182 9516 9523 9520 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08181 9514 9516 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08180 11074 9516 9514 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08179 2001 5501 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08178 2003 2000 2002 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08177 1485 1495 1488 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08176 1488 1494 1486 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08175 1487 1493 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08174 1483 1490 1488 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08173 11074 1489 1482 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08172 11074 1496 1484 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08171 1834 1488 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08170 10783 10184 10185 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08169 10185 10194 10783 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08168 11074 10182 10183 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08167 3194 5727 3195 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08166 3196 5728 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08165 3817 10257 3194 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08164 9645 9649 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08163 9644 9648 9647 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08162 9640 9650 9643 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08161 11074 9947 9640 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08160 11074 10638 9650 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08159 9648 9650 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08158 11074 9946 9649 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08157 9647 9650 9645 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08156 9641 9647 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08155 11074 9642 9646 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08154 9643 9648 9642 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08153 9947 9643 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08152 11074 9643 9947 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08151 10598 10596 10449 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08150 10449 10595 10598 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08149 11074 10594 10449 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08148 10897 10598 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08147 10148 10147 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08146 11012 10582 10149 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08145 4233 4363 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08144 4476 4364 4234 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08143 11074 1556 1558 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_08142 1558 3714 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_08141 2776 1557 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08140 1558 3057 1557 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_08139 1557 4014 1558 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_08138 6817 8318 6661 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08137 6661 8316 6817 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08136 11074 8691 6662 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08135 10794 10798 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08134 10793 10797 10795 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08133 10788 10799 10787 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08132 11074 10838 10788 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08131 11074 10914 10799 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08130 10797 10799 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08129 11074 10796 10798 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08128 10795 10799 10794 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08127 10790 10795 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08126 11074 10792 10791 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08125 10787 10797 10792 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08124 10838 10787 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08123 11074 10787 10838 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08122 7386 7539 7385 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08121 7387 7538 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08120 7383 7534 7382 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08119 7535 10697 7384 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08118 9685 10083 9684 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08117 9687 10709 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08116 9686 10700 9685 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08115 1151 3735 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08114 1302 9597 1152 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08113 2597 2167 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08112 11074 2165 2597 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08111 2597 2581 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08110 11074 2166 2597 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08109 2491 2211 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08108 11074 2212 2491 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08107 2491 2208 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08106 11074 2209 2491 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08105 11074 4926 4108 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08104 4109 4916 4280 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08103 4279 4280 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08102 8541 8671 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08101 8539 8672 8668 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08100 8537 8673 8664 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08099 11074 8694 8537 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08098 11074 10914 8673 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08097 8672 8673 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08096 11074 8670 8671 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08095 8668 8673 8541 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08094 8538 8668 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08093 11074 8667 8540 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08092 8664 8672 8667 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08091 8694 8664 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08090 11074 8664 8694 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08089 3522 3685 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08088 3521 3686 3683 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08087 3519 3687 3679 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08086 11074 8297 3519 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08085 11074 5083 3687 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08084 3686 3687 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_08083 11074 3684 3685 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_08082 3683 3687 3522 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08081 3520 3683 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08080 11074 3680 3523 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08079 3679 3686 3680 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08078 8297 3679 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08077 11074 3679 8297 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08076 8264 8262 8263 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08075 8263 9290 8264 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08074 11074 9987 8263 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08073 8261 8264 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08072 11074 7457 7277 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08071 7278 7685 7458 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08070 7670 7458 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08069 7697 7695 7699 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08068 7698 7702 7697 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08067 7700 7704 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08066 8327 7697 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08065 11074 7719 7696 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08064 7698 7701 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_08063 7393 9057 7392 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08062 7397 9421 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08061 7395 9433 7394 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08060 7539 9716 7396 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08059 7373 9433 7371 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08058 7372 10697 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08057 9046 9716 7373 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08056 10159 10158 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08055 11039 10279 10160 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_08054 10398 10710 10396 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08053 10397 10395 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08052 10693 11072 10398 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08051 4205 4952 4204 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08050 4207 4631 4315 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08049 11074 4955 4206 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08048 4314 4315 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_08047 1633 2384 1631 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08046 1632 1973 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08045 1804 2403 1633 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08044 11074 1810 1639 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08043 1640 7426 1808 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08042 2393 1808 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08041 5149 6214 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08040 5147 6215 5146 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08039 11074 6213 5147 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08038 5148 5147 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08037 4590 5159 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08036 4589 6127 4588 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08035 11074 6213 4589 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08034 4587 4589 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08033 6892 8459 6704 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08032 6704 7535 6892 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08031 11074 6890 6704 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08030 6891 6892 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08029 7179 9083 7178 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08028 7180 11066 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08027 7182 10399 7181 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08026 7177 9716 7183 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08025 7783 8429 7782 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08024 7785 8049 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08023 7784 8426 7783 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08022 8579 9073 8577 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08021 8578 9418 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08020 8753 9051 8579 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08019 2915 3068 2916 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08018 2917 3069 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08017 3375 4349 2915 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08016 11074 10697 7374 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08015 7375 7534 7530 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08014 7531 7530 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08013 9227 10698 9225 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08012 9226 10073 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08011 9417 11072 9227 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08010 6410 6408 6413 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08009 11074 9566 6411 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08008 6414 6764 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08007 6413 6409 6412 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08006 6326 6764 6408 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08005 6409 9566 6325 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08004 11074 5610 5027 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08003 11074 5024 5027 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08002 5027 5286 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_08001 5023 5027 4870 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_08000 4188 4250 4371 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07999 4371 5023 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07998 4374 4371 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07997 11074 10702 10504 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07996 10505 10706 10703 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07995 11057 10703 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07994 8446 9080 8449 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07993 8448 9702 8450 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07992 11074 9057 8447 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07991 8728 8450 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07990 10217 10578 10216 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07989 10216 10577 10217 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07988 11074 10838 10216 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07987 10214 10217 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07986 4774 4951 6205 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07985 11074 4948 4772 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07984 4775 4950 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07983 6205 4947 4776 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07982 4777 4950 4951 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07981 4947 4948 4773 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07980 11074 4352 4008 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07979 10028 4008 4007 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07978 11074 4008 10028 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07977 11074 4008 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07976 11024 4008 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07975 11074 4352 1066 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07974 9597 1066 1065 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07973 11074 1066 9597 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07972 11074 1066 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07971 11024 1066 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07970 11074 4352 4353 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07969 8643 4353 4182 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07968 11074 4353 8643 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07967 11074 4353 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07966 11024 4353 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07965 11074 4352 3361 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07964 9308 3361 3362 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07963 11074 3361 9308 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07962 11074 3361 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07961 11024 3361 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07960 11074 4352 4346 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07959 8921 4346 4181 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07958 11074 4346 8921 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07957 11074 4346 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07956 11024 4346 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07955 11074 487 486 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07954 4352 486 485 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07953 11074 486 4352 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07952 11074 486 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07951 11024 486 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07950 4217 5275 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07949 4349 5901 4218 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07948 4216 4694 4349 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07947 11074 4347 4216 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07946 4216 4348 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07945 11074 5897 5311 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07944 5308 5307 5310 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07943 5309 5310 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07942 11074 1601 1599 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07941 5293 1599 1598 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07940 11074 1599 5293 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07939 11074 1599 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07938 11024 1599 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07937 11074 1601 1602 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07936 5607 1602 1600 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07935 11074 1602 5607 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07934 11074 1602 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07933 11024 1602 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07932 11074 1308 1309 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07931 1601 1309 1183 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07930 11074 1309 1601 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07929 11074 1309 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07928 11024 1309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07927 9291 9287 9125 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07926 11074 10197 9289 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07925 9126 9289 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07924 76 747 75 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07923 77 482 214 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07922 11074 219 74 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07921 437 214 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07920 2861 9560 2860 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07919 2862 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07918 2859 10028 2863 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07917 3028 3027 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07916 3027 2858 2859 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07915 3970 3969 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07914 9609 5599 3971 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07913 3968 9308 9609 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07912 11074 3974 3968 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07911 3968 3967 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07910 3404 3402 3407 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07909 3405 3403 3406 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07908 11074 4043 3401 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07907 4054 3406 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07906 6432 9566 6433 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07905 6433 7437 6432 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07904 11074 9310 6433 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07903 6431 6432 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07902 7931 8133 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07901 7930 8134 8132 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07900 7927 8135 8130 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07899 11074 8725 7927 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07898 11074 10638 8135 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07897 8134 8135 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07896 11074 8724 8133 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07895 8132 8135 7931 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07894 7928 8132 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07893 11074 8131 7929 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07892 8130 8134 8131 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07891 8725 8130 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07890 11074 8130 8725 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07889 7144 7161 7145 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07888 7145 9046 7144 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07887 11074 7142 7146 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07886 6390 6388 6402 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07885 11074 8893 6391 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07884 6393 6759 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07883 6402 6389 6392 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07882 6315 6759 6388 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07881 6389 8893 6314 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07880 1757 9560 1760 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07879 1761 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07878 1759 7678 1758 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07877 2172 1889 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07876 1889 1787 1759 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07875 1594 5600 1597 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07874 1595 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07873 1592 5918 1596 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07872 3082 1593 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07871 1593 1591 1592 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07870 4783 5185 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07869 4959 5183 4784 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07868 4603 5181 4606 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07867 4604 4952 4603 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07866 4607 5842 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07865 4602 4603 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07864 11074 4960 4605 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07863 4604 5175 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07862 391 395 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07861 390 394 393 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07860 386 396 388 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07859 11074 959 386 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07858 11074 2446 396 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07857 394 396 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07856 11074 963 395 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07855 393 396 391 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07854 387 393 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07853 11074 389 392 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07852 388 394 389 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07851 959 388 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07850 11074 388 959 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07849 7103 7104 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07848 7100 7106 7101 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07847 7097 7105 7096 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07846 11074 7109 7097 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07845 11074 8048 7105 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07844 7106 7105 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07843 11074 7108 7104 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07842 7101 7105 7103 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07841 7095 7101 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07840 11074 7099 7102 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07839 7096 7106 7099 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07838 7109 7096 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07837 11074 7096 7109 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07836 7470 9610 7289 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07835 7289 8644 7470 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07834 11074 7468 7289 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07833 7467 7470 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07832 8204 8885 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07831 8206 9033 8205 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07830 8230 8733 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07829 9028 8411 8231 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07828 6283 6286 6071 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07827 6071 6901 6283 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07826 11074 6282 6071 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07825 6177 6283 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07824 5931 6286 5932 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07823 5932 6905 5931 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07822 11074 5933 5929 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07821 4475 4723 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07820 4726 4472 4473 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07819 5184 5181 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07818 5183 6246 5182 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07817 2828 7432 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07816 3844 2989 2829 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07815 4299 4301 4122 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07814 4122 4942 4299 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07813 11074 4940 4122 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07812 4298 4299 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07811 7977 10689 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07810 8050 8746 7978 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07809 7346 8733 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07808 7520 7516 7347 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07807 7356 9083 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07806 7525 8746 7357 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07805 6686 8733 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07804 7517 7117 6687 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07803 7850 10704 7849 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07802 7849 8063 7850 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07801 11074 8062 7849 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07800 7848 7850 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07799 4874 5312 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07798 5037 5038 4875 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07797 4236 4478 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07796 4472 4369 4235 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07795 629 1545 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07794 747 8713 630 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07793 7878 10567 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07792 8086 8635 7876 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07791 7877 8636 8086 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07790 11074 8082 7877 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07789 7874 8930 8086 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07788 11074 8633 7875 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07787 13 2630 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07786 2637 2385 12 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07785 10474 10649 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07784 10471 10650 10648 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07783 10470 10651 10643 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07782 11074 10641 10470 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07781 11074 11051 10651 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07780 10650 10651 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07779 11074 10646 10649 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07778 10648 10651 10474 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07777 10472 10648 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07776 11074 10644 10473 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07775 10643 10650 10644 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07774 10641 10643 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07773 11074 10643 10641 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07772 7238 10027 7237 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07771 7239 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07770 7419 7418 7238 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07769 11074 1300 1038 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07768 11074 1301 1038 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07767 1038 1040 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07766 1288 1038 1039 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07765 10900 9566 9567 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07764 9567 9609 10900 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07763 11074 9594 9565 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07762 1732 6276 1730 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07761 1731 8661 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07760 2121 5599 1732 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07759 7985 10701 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07758 8052 11072 7986 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07757 5892 6286 5893 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07756 5893 6895 5892 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07755 11074 5890 5893 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07754 5891 5892 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07753 11074 9998 9779 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07752 9780 10000 9999 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07751 9994 9999 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07750 11074 5539 4129 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07749 4130 4323 4317 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07748 4316 4317 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07747 10848 10849 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07746 10844 10850 10846 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07745 10842 10851 10841 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07744 11074 10854 10842 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07743 11074 10914 10851 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07742 10850 10851 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07741 11074 10853 10849 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07740 10846 10851 10848 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07739 10840 10846 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07738 11074 10843 10845 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07737 10841 10850 10843 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07736 10854 10841 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07735 11074 10841 10854 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07734 11074 8709 7313 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07733 7311 10995 7312 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07732 7483 7740 7320 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_07731 7312 7481 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07730 7310 8709 7481 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_07729 7480 7486 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_07728 7321 7727 7314 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07727 7316 7740 7315 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07726 7318 7483 7317 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07725 7319 7484 7321 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07724 531 1268 530 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07723 11074 689 690 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07722 11074 1268 533 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07721 534 5510 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07720 535 647 534 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07719 532 691 531 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07718 690 689 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07717 995 1268 993 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07716 11074 1266 1265 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07715 11074 1268 999 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07714 1000 5544 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07713 994 1270 1000 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07712 996 1490 995 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07711 1265 1266 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07710 942 1268 940 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07709 11074 931 934 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07708 11074 1268 943 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07707 944 5707 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07706 941 937 944 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07705 938 951 942 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07704 934 931 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07703 987 1268 986 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07702 11074 982 983 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07701 11074 1268 990 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07700 991 5732 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07699 989 988 991 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07698 985 984 987 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07697 983 982 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07696 370 1268 369 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07695 11074 374 368 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07694 11074 1268 375 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07693 372 5531 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07692 373 376 372 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07691 371 706 370 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07690 368 374 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07689 3964 6276 3965 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07688 3966 8661 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07687 7068 5898 3964 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07686 1736 2763 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07685 1877 4325 1737 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07684 9136 9309 9140 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07683 9141 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07682 9138 9308 9137 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07681 10003 9304 9139 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07680 11074 4410 2832 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07679 2833 2996 2995 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07678 3202 2995 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07677 9927 10614 9793 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07676 9793 10615 9927 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07675 11074 10594 9792 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07674 7283 7685 7282 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07673 7284 7684 7464 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07672 11074 7465 7285 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07671 7463 7464 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07670 400 1268 398 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07669 11074 402 397 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07668 11074 1268 403 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07667 404 3277 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07666 399 405 404 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07665 401 723 400 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07664 397 402 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07663 918 1841 924 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07662 11074 1237 1235 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07661 11074 1841 927 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07660 921 4910 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07659 922 1239 921 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07658 919 1403 918 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07657 1235 1237 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07656 1393 1841 1390 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07655 11074 1387 1388 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07654 11074 1841 1394 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07653 1391 4905 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07652 1392 1395 1391 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07651 1389 1396 1393 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07650 1388 1387 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07649 909 1841 908 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07648 11074 1232 1230 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07647 11074 1841 914 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07646 912 5510 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07645 913 1234 912 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07644 910 1813 909 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07643 1230 1232 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07642 6976 6992 6975 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07641 6977 9313 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07640 6971 8122 6974 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07639 6994 7655 6972 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07638 4167 5719 4165 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07637 4166 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07636 4666 7678 4167 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07635 8478 9100 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07634 11074 8475 8478 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07633 8478 9974 8476 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07632 8479 8477 8478 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07631 11074 4036 3073 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07630 11074 3072 3073 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07629 3073 3071 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07628 5029 3073 2921 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07627 5222 7478 5221 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07626 5223 5719 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07625 5218 9597 5217 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07624 5220 7739 5219 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07623 3839 5727 3838 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07622 3840 5728 3842 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07621 11074 10231 3841 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07620 3837 3842 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07619 2631 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07618 2630 3618 2629 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07617 2628 2971 2630 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07616 11074 5124 2628 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07615 2628 2967 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07614 2305 8709 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07613 11074 3714 2305 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07612 2305 2572 2303 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07611 2304 4014 2305 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07610 9160 10197 9612 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07609 9164 10197 9320 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07608 9161 10020 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07607 9163 9320 9162 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07606 11074 9316 9159 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07605 11074 4036 4041 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07604 11074 4042 4041 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07603 4041 4037 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07602 5018 4041 4035 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07601 11074 4929 3222 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07600 3217 4936 3218 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07599 3223 3242 3146 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_07598 3218 3216 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07597 3145 4929 3216 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_07596 3651 3228 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_07595 3229 3219 3220 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07594 3221 3242 3224 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07593 3226 3223 3225 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07592 3227 3889 3229 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07591 11074 4929 3204 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07590 3200 3198 3201 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07589 3209 3242 3144 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_07588 3201 3199 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07587 3143 4929 3199 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_07586 4285 3203 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_07585 3211 3202 3205 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07584 3207 3242 3206 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07583 3208 3209 3212 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07582 3210 3884 3211 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_07581 11074 5764 5765 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07580 10891 5765 5763 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07579 11074 5765 10891 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07578 11074 5765 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07577 11024 5765 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07576 11074 5168 5170 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07575 5764 5170 5169 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07574 11074 5170 5764 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07573 11074 5170 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07572 11024 5170 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07571 7713 7721 7718 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07570 7714 7711 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07569 7716 9308 7715 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07568 8113 7717 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07567 7717 7712 7716 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07566 8842 10197 9955 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07565 8847 10197 8846 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07564 8843 9489 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07563 8845 8846 8844 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07562 11074 8840 8841 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07561 11077 11075 11078 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07560 11078 11076 11077 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07559 11074 11072 11073 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07558 484 4680 483 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07557 483 1545 484 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07556 11074 4684 483 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07555 482 484 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07554 11074 8101 7881 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07553 7882 8086 8085 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07552 8014 8085 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07551 11074 1855 1696 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07550 1695 1857 1856 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07549 5557 1856 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07548 11074 5764 5540 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07547 10604 5540 5396 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07546 11074 5540 10604 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07545 11074 5540 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07544 11024 5540 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07543 6984 6988 7007 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07542 11074 8122 6981 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07541 6985 6992 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07540 7007 6983 6986 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07539 6987 6992 6988 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07538 6983 8122 6982 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07537 8068 8620 7953 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07536 7954 10258 8068 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07535 7955 8621 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07534 8000 8068 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07533 11074 10256 7956 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07532 7954 10269 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07531 538 1495 694 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07530 694 1494 539 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07529 541 916 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07528 536 691 694 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07527 11074 1489 537 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07526 11074 692 540 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07525 2412 694 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07524 9322 9612 9165 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07523 9165 9347 9322 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07522 11074 9603 9165 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07521 9321 9322 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07520 3476 3647 3649 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07519 3649 3879 3477 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07518 3478 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07517 3473 3652 3649 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07516 11074 4290 3474 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07515 11074 3646 3475 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07514 3872 3649 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07513 1616 1795 1793 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07512 11074 2962 1617 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07511 1618 2964 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07510 1793 1792 1619 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07509 1620 2964 1795 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07508 1792 2962 1615 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07507 11074 6815 6463 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07506 10018 6463 6464 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07505 11074 6463 10018 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07504 11074 6463 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07503 11024 6463 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07502 11074 6815 6816 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07501 7615 6816 6660 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07500 11074 6816 7615 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07499 11074 6816 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07498 11024 6816 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07497 11074 6228 6229 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07496 6815 6229 6003 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07495 11074 6229 6815 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07494 11074 6229 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07493 11024 6229 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07492 7974 8430 7973 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07491 7976 8753 8148 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07490 11074 8443 7975 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07489 8049 8148 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07488 11074 10708 9841 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07487 9842 10073 10052 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07486 9958 10052 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07485 3622 3837 3443 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07484 3443 4567 3622 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07483 11074 4553 3443 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07482 3621 3622 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07481 4927 4925 4758 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07480 4758 5140 4927 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07479 11074 4926 4758 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07478 5128 4927 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07477 5228 5229 5227 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07476 5227 5226 5228 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07475 11074 9987 5227 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07474 6497 5228 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07473 10584 8893 8894 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07472 8894 9609 10584 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07471 11074 9541 8892 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07470 7405 7404 7225 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07469 7224 10258 7405 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07468 7226 7583 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07467 7403 7405 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07466 11074 10256 7223 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07465 7224 10269 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_07464 1876 2140 1733 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07463 1733 2138 1876 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07462 11074 1873 1733 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07461 1874 1876 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07460 770 8124 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07459 11074 3092 770 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07458 5129 5132 5130 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07457 5130 5128 5129 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07456 11074 5681 5130 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07455 5704 5129 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07454 2428 3008 2275 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07453 2275 3009 2428 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07452 11074 2688 2275 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07451 3000 2428 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07450 4503 5098 4502 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07449 4502 6195 4503 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07448 11074 4500 4502 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07447 4501 4503 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07446 413 415 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07445 408 414 412 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07444 406 416 407 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07443 11074 984 406 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07442 11074 2446 416 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07441 414 416 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07440 11074 983 415 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07439 412 416 413 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07438 409 412 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07437 11074 411 410 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07436 407 414 411 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07435 984 407 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07434 11074 407 984 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07433 6700 6887 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07432 6699 6886 6884 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07431 6697 6888 6881 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07430 11074 6879 6697 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07429 11074 8048 6888 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07428 6886 6888 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07427 11074 6891 6887 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07426 6884 6888 6700 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07425 6698 6884 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07424 11074 6882 6701 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07423 6881 6886 6882 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07422 6879 6881 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07421 11074 6881 6879 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07420 9047 9061 9049 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07419 9049 9046 9047 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07418 11074 9044 9048 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07417 10036 6819 6482 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07416 6482 6489 10036 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07415 11074 6490 6481 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07414 1782 3734 1781 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07413 1785 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07412 1784 5600 1783 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07411 2209 1903 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07410 1903 1790 1784 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07409 4865 5014 4864 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07408 4866 5015 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07407 4868 5908 4867 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07406 5033 5016 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07405 5016 4863 4868 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07404 637 7042 636 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07403 638 3033 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07402 640 1881 639 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07401 753 754 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07400 754 635 640 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07399 314 318 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07398 313 317 316 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07397 309 319 311 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07396 11074 338 309 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07395 11074 2673 319 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07394 317 319 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07393 11074 320 318 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07392 316 319 314 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07391 310 316 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07390 11074 312 315 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07389 311 317 312 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07388 338 311 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07387 11074 311 338 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07386 11074 9987 9983 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07385 9763 9983 9982 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07384 11074 10213 9763 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07383 10176 9982 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07382 11074 9982 10176 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07381 10035 10608 9818 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07380 9818 10606 10035 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07379 11074 10641 9818 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07378 10033 10035 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07377 11074 3032 3292 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07376 3292 3028 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07375 2864 3029 3292 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07374 4142 3958 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07373 11074 3959 4142 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07372 4142 4979 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07371 11074 4976 4142 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07370 2970 3628 2805 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07369 2805 2971 2970 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07368 11074 2967 2805 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07367 2968 2970 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07366 10270 10272 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07365 10154 10156 10155 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07364 10150 10271 10267 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07363 11074 10268 10150 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07362 11074 10638 10271 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07361 10156 10271 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07360 11074 11018 10272 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07359 10155 10271 10270 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07358 10151 10155 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07357 11074 10153 10152 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07356 10267 10156 10153 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07355 10268 10267 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07354 11074 10267 10268 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07353 6607 8612 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07352 6749 10915 6608 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07351 9394 9686 9205 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07350 9205 9680 9394 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07349 11074 9392 9204 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07348 1663 5672 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07347 2024 1824 1664 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07346 10290 10293 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07345 10165 10167 10166 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07344 10161 10291 10288 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07343 11074 10289 10161 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07342 11074 11051 10291 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07341 10167 10291 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07340 11074 10292 10293 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07339 10166 10291 10290 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07338 10162 10166 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07337 11074 10164 10163 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07336 10288 10167 10164 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07335 10289 10288 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07334 11074 10288 10289 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07333 5941 6186 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07332 5938 6187 6185 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07331 5937 6188 6183 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07330 11074 10771 5937 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07329 11074 10914 6188 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07328 6187 6188 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07327 11074 10781 6186 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07326 6185 6188 5941 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07325 5939 6185 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07324 11074 6184 5940 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07323 6183 6187 6184 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07322 10771 6183 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07321 11074 6183 10771 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07320 11070 11066 11068 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07319 11069 11067 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07318 11071 11077 11070 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07317 10503 10701 10501 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07316 10502 10709 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07315 10707 10700 10503 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07314 1162 3735 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07313 1552 3734 1163 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07312 854 3735 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07311 1873 5599 855 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07310 11074 8713 4145 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07309 4144 4327 4328 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07308 4640 4328 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07307 5726 9566 5725 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07306 5725 7437 5726 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07305 11074 9310 5724 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07304 11074 6195 4504 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07303 4506 5098 4505 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07302 5094 4505 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07301 8978 8980 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07300 8974 8981 8979 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07299 8972 8982 8971 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07298 11074 8970 8972 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07297 11074 10638 8982 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07296 8981 8982 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07295 11074 8977 8980 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07294 8979 8982 8978 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07293 8975 8979 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07292 11074 8973 8976 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07291 8971 8981 8973 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07290 8970 8971 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07289 11074 8971 8970 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07288 6041 10687 6042 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07287 11074 6274 6164 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07286 11074 10687 6043 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07285 6039 6894 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07284 6040 6167 6039 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07283 6038 6163 6041 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07282 6164 6274 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07281 8554 8733 8734 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07280 8556 8733 8735 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07279 8557 10382 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07278 8559 8735 8558 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07277 11074 8731 8555 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07276 3261 3288 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07275 3263 6137 3262 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07274 10425 10555 10424 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07273 10426 10546 10549 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07272 11074 10547 10427 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07271 10780 10549 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07270 11074 10018 9539 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07269 9542 9541 9543 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07268 9540 9543 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07267 11074 10576 10573 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07266 10440 10573 10572 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07265 11074 10570 10440 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07264 10571 10572 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07263 11074 10572 10571 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07262 11074 5564 4799 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07261 4800 5216 4980 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07260 4979 4980 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07259 3894 4584 3896 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07258 11074 3899 3893 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07257 11074 4584 3900 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07256 3897 4617 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07255 3898 3901 3897 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07254 3895 4553 3894 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_07253 3893 3899 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07252 9916 9985 9765 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07251 9765 9989 9916 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07250 11074 9986 9764 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07249 11074 10170 9876 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07248 9877 10080 10079 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07247 9979 10079 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07246 2693 2691 2694 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07245 2694 2692 2693 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07244 11074 6132 2695 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07243 2600 3086 2790 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07242 2790 3088 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07241 2796 2790 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07240 11074 4066 4069 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07239 4067 4069 4068 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07238 11074 4070 4067 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07237 5035 4068 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07236 11074 4068 5035 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07235 4856 5008 5010 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07234 5010 5009 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07233 5603 5010 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07232 3308 3322 3313 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07231 3312 3311 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07230 3310 3306 3309 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07229 3962 5771 3307 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07228 10196 10619 10195 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07227 10195 10564 10196 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07226 11074 10554 10195 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07225 10194 10196 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07224 5982 6277 5981 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07223 5983 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07222 5985 9597 5984 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07221 6127 8082 5986 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07220 7993 9087 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07219 8056 9750 7991 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07218 7992 9107 8056 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07217 11074 9103 7992 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07216 7992 8460 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_07215 4161 8126 4159 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07214 4160 7478 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07213 8713 10028 4161 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07212 7838 9729 7839 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07211 7839 8060 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07210 7837 7839 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07209 6791 2006 2007 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07208 2007 2004 6791 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07207 11074 4325 2005 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07206 2123 2121 2122 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07205 2124 2470 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07204 2118 2480 2125 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07203 2119 2120 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07202 2120 2117 2118 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07201 2564 7069 2563 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07200 2565 6221 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07199 2567 3057 2566 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07198 2727 2726 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07197 2726 2562 2567 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07196 4112 4283 4543 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07195 11074 4285 4113 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07194 4115 4286 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07193 4543 4284 4116 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07192 4117 4286 4283 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07191 4284 4285 4114 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07190 8856 8629 8492 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07189 8492 9295 8856 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07188 11074 8627 8493 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07187 11074 5504 5342 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07186 5343 6381 5502 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07185 5501 5502 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07184 6224 6455 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07183 11074 10891 6224 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07182 6224 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07181 11074 10888 6224 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07180 6142 6224 5996 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07179 11074 7023 7024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07178 7026 7451 7025 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07177 7022 7025 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07176 10902 10915 10908 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07175 10904 10915 10912 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07174 10905 10909 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07173 10907 10912 10906 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07172 11074 10901 10903 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07171 853 3413 1048 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07170 1048 2473 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07169 2474 1048 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07168 11074 4064 4065 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07167 11074 4463 4065 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07166 4065 5304 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07165 4063 4065 4062 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07164 11074 5600 3323 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07163 3324 8661 3325 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07162 3698 3325 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07161 11074 6809 5995 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07160 5994 6806 6222 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07159 6141 6222 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07158 11074 8650 8521 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07157 8522 8652 8653 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07156 8651 8653 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07155 11074 2741 2742 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07154 2744 2746 2743 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07153 3311 2743 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07152 11074 5719 3544 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07151 3543 5919 3707 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07150 4653 3707 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07149 5787 10029 5786 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07148 5789 5919 5790 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07147 11074 8643 5788 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07146 8316 5790 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07145 5315 5320 5314 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07144 5317 5313 5316 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07143 11074 6182 5318 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07142 5312 5316 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07141 5943 6191 6106 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07140 11074 6387 5944 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07139 5946 6192 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07138 6106 6190 5945 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07137 5947 6192 6191 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07136 6190 6387 5942 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07135 4853 7478 4852 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07134 4854 9560 5007 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07133 11074 10028 4855 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07132 5273 5007 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_07131 11074 8124 511 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07130 512 3092 513 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07129 510 513 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07128 9312 9509 9150 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07127 9150 9347 9312 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07126 11074 9594 9150 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07125 9310 9312 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07124 1807 1802 1630 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07123 1630 1801 1807 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07122 11074 2679 1629 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07121 3419 3423 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07120 3421 3422 3420 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07119 3414 3424 3417 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07118 11074 3413 3414 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07117 11074 5262 3424 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07116 3422 3424 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07115 11074 5034 3423 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07114 3420 3424 3419 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07113 3415 3420 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07112 11074 3416 3418 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07111 3417 3422 3416 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07110 3413 3417 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07109 11074 3417 3413 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07108 8418 8419 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07107 8226 8229 8228 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07106 8224 8420 8410 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07105 11074 8411 8224 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07104 11074 10638 8420 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07103 8229 8420 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07102 11074 9030 8419 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07101 8228 8420 8418 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07100 8223 8228 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07099 11074 8225 8227 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07098 8410 8229 8225 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07097 8411 8410 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07096 11074 8410 8411 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07095 11074 7098 4989 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07094 9987 4989 4806 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07093 11074 4989 9987 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07092 11074 4989 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07091 11024 4989 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07090 11074 7098 5225 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07089 10915 5225 5224 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07088 11074 5225 10915 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07087 11074 5225 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07086 11024 5225 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07085 11074 7098 7073 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07084 10774 7073 7074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07083 11074 7073 10774 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07082 11074 7073 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07081 11024 7073 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07080 11074 7098 7076 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07079 10197 7076 7075 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07078 11074 7076 10197 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07077 11074 7076 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07076 11024 7076 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07075 11074 5611 5612 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07074 7098 5612 5486 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07073 11074 5612 7098 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07072 11074 5612 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07071 11024 5612 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07070 2348 5600 2347 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07069 2349 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07068 2351 5719 2350 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07067 2499 2498 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07066 2498 2346 2351 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07065 2792 2500 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07064 11074 2499 2792 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07063 9100 9430 9097 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07062 9097 9095 9100 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07061 11074 9747 9096 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07060 1747 1881 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07059 11074 3714 1747 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07058 1747 6220 1745 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07057 1746 4014 1747 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07056 4781 5181 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07055 4954 7109 4780 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07054 433 434 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07053 430 435 432 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07052 426 436 428 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07051 11074 729 426 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07050 11074 5262 436 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07049 435 436 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07048 11074 743 434 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07047 432 436 433 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07046 427 432 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07045 11074 429 431 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07044 428 435 429 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07043 729 428 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07042 11074 428 729 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07041 10238 10596 10237 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07040 10237 10595 10238 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07039 11074 10312 10237 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07038 10600 10238 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07037 2186 5898 2185 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07036 2187 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07035 2189 7514 2188 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07034 2590 2184 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_07033 2184 2183 2189 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07032 3924 3945 3923 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07031 3923 3925 3924 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07030 11074 3922 3923 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07029 4948 3924 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07028 6018 6249 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07027 6016 6250 6248 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07026 6015 6252 6245 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07025 11074 6246 6015 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07024 11074 8048 6252 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07023 6250 6252 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_07022 11074 7131 6249 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_07021 6248 6252 6018 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07020 6014 6248 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07019 11074 6247 6017 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07018 6245 6250 6247 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07017 6246 6245 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07016 11074 6245 6246 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07015 7040 10027 7038 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07014 7039 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07013 7036 7037 7040 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07012 8213 8709 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07011 8212 8713 8214 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07010 9026 10687 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07009 9678 9667 9027 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07008 9018 10687 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07007 9392 9382 9017 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_07006 4175 5191 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07005 4178 5191 4337 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_07004 11074 7484 4173 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07003 4339 4336 4176 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07002 4177 4337 4339 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07001 4335 4339 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_07000 11074 4339 4335 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06999 4336 7484 4174 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06998 5874 8051 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06997 5873 6574 5875 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06996 10972 10974 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06995 10966 10973 10971 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06994 10964 10975 10965 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06993 11074 10963 10964 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06992 11074 11051 10975 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06991 10973 10975 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06990 11074 10970 10974 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06989 10971 10975 10972 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06988 10967 10971 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06987 11074 10969 10968 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06986 10965 10973 10969 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06985 10963 10965 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06984 11074 10965 10963 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06983 7287 7685 7286 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06982 7288 7684 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06981 8834 7465 7287 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06980 8234 10689 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06979 8750 9080 8235 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06978 1012 1248 1013 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06977 11074 1006 1008 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06976 11074 1248 1014 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06975 1010 5732 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06974 1011 1009 1010 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06973 1007 1005 1012 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06972 1008 1006 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06971 5734 5736 5733 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06970 11074 5739 5732 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06969 11074 5736 5740 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06968 5737 6788 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06967 5738 5742 5737 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06966 5735 11018 5734 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06965 5732 5739 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06964 6363 10704 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06963 6569 9716 6364 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06962 5278 5293 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06961 5279 5275 5276 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06960 5277 6278 5279 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06959 11074 10606 5277 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06958 5277 5273 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06957 5398 6221 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06956 5542 6220 5397 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06955 11074 5541 5542 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06954 5756 5542 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06953 2633 2982 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06952 2635 3625 2634 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06951 11074 3632 2635 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06950 2632 2635 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06949 11074 6215 5374 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06948 5375 6214 5524 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06947 5523 5524 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06946 4311 2434 2280 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06945 2280 2435 4311 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06944 11074 2688 2279 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06943 4135 5727 4134 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06942 4136 5728 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06941 4323 10995 4135 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06940 3920 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06939 3941 4316 3921 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06938 3919 4307 3941 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06937 11074 5124 3919 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06936 3919 3917 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06935 8835 8893 7862 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06934 7862 8644 8835 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06933 11074 8070 7861 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06932 7633 7445 7259 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06931 7259 7667 7633 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06930 11074 10774 7258 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06929 10384 10700 10386 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06928 10385 10392 10384 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06927 10387 10701 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06926 10382 10384 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06925 11074 10693 10383 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06924 10385 10694 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06923 7968 9710 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06922 8042 8429 7967 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06921 1683 1841 1682 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06920 11074 1842 1839 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06919 11074 1841 1685 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06918 1686 5544 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06917 1687 1845 1686 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06916 1684 1844 1683 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06915 1839 1842 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06914 1440 1841 1439 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06913 11074 1436 1437 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06912 11074 1841 1443 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06911 1444 5707 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06910 1441 1442 1444 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06909 1438 1826 1440 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06908 1437 1436 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06907 4164 9560 4162 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06906 4163 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06905 6251 9308 4164 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06904 4158 8922 4156 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06903 4157 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06902 7465 8921 4158 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06901 2137 9560 2135 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06900 2136 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06899 2572 5898 2137 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06898 9260 10414 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06897 9432 10686 9261 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06896 5472 5600 5471 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06895 5473 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06894 5475 9560 5474 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06893 5906 5599 5476 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06892 6068 6574 6067 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06891 6069 8770 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06890 6064 10704 6070 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06889 6176 7852 6065 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06888 6084 6221 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06887 8636 6220 6085 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06886 11074 10774 10779 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06885 10775 10779 10776 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06884 11074 10838 10775 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06883 10773 10776 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06882 11074 10776 10773 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06881 5242 7478 5241 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06880 5243 6277 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06879 5238 8643 5244 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06878 5240 5851 5239 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06877 11074 2989 2830 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06876 2831 7432 2990 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06875 3635 2990 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06874 11074 3925 3515 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06873 3516 3945 3674 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06872 3675 3674 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06871 9896 10013 9895 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06870 9897 10015 10012 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06869 11074 10014 9898 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06868 10005 10012 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06867 9882 10542 9881 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06866 9883 10566 9990 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06865 11074 10541 9884 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06864 9989 9990 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06863 1673 1841 1675 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06862 11074 1832 2047 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06861 11074 1841 1678 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06860 1676 5732 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06859 1677 1833 1676 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06858 1674 2038 1673 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06857 2047 1832 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06856 972 1841 971 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06855 11074 1263 1260 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06854 11074 1841 979 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06853 975 5531 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06852 976 1264 975 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06851 973 1456 972 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06850 1260 1263 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06849 1464 1841 1463 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06848 11074 1460 1461 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06847 11074 1841 1467 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06846 1465 3277 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06845 1466 1470 1465 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06844 1462 2432 1464 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06843 1461 1460 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06842 936 1284 935 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06841 11074 1241 1431 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06840 11074 1284 939 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06839 932 4910 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06838 933 1243 932 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06837 930 1423 936 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06836 1431 1241 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06835 351 1284 354 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06834 11074 353 347 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06833 11074 1284 355 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06832 349 4905 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06831 350 356 349 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06830 352 348 351 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06829 347 353 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06828 4153 6277 4154 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06827 4155 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06826 7069 8643 4153 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06825 2173 2172 2174 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06824 2174 2177 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06823 2581 2174 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06822 11074 4929 3847 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06821 3845 3844 3848 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06820 3858 5150 3856 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_06819 3848 3846 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06818 3843 4929 3846 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_06817 4272 3854 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_06816 3859 3849 3855 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06815 3851 5150 3850 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06814 3853 3858 3852 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06813 3857 4530 3859 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06812 11074 4929 3462 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06811 3459 3635 3460 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06810 3640 5150 3468 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_06809 3460 3636 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06808 3458 4929 3636 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_06807 4275 3642 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_06806 3469 3637 3461 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06805 3463 5150 3467 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06804 3465 3640 3464 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06803 3466 4535 3469 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_06802 7707 8092 7706 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06801 7708 8709 7710 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06800 11074 8713 7709 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06799 7704 7710 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06798 544 1284 542 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06797 11074 696 925 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06796 11074 1284 546 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06795 547 5510 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06794 543 650 547 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06793 545 916 544 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06792 925 696 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06791 1015 1284 1017 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06790 11074 1283 1280 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06789 11074 1284 1021 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06788 1018 5544 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06787 1019 1285 1018 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06786 1016 1493 1015 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06785 1280 1283 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06784 2127 6275 2126 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06783 2128 6276 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06782 2470 6277 2127 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06781 8469 10710 8468 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06780 8470 11076 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06779 8466 9405 8471 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06778 8477 10700 8467 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06777 6603 9057 6602 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06776 6601 8059 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06775 6599 8746 6598 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06774 6905 9433 6600 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06773 7218 8453 7221 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06772 7222 9080 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06771 7220 8770 7219 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06770 7217 9433 7216 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06769 6090 6232 6089 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06768 6091 6457 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06767 6088 6251 6087 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06766 10578 6227 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06765 6227 6086 6088 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06764 11074 6537 6539 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06763 6541 7532 6540 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06762 6538 6540 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06761 11074 10697 6688 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06760 6689 7798 6865 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06759 6866 6865 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06758 11074 10915 1505 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06757 1506 1519 1507 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06756 1504 1507 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06755 10617 10619 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06754 11074 10891 10617 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06753 10617 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06752 11074 10888 10617 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06751 10618 10617 10457 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06750 4767 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06749 4943 4944 4768 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06748 4769 4942 4943 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06747 11074 5124 4769 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06746 4769 4940 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06745 8509 9287 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06744 8641 8834 8510 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06743 11074 8645 8641 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06742 8862 8641 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06741 11074 6259 6026 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06740 6027 8733 6258 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06739 7129 6258 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06738 11074 489 237 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06737 5919 237 106 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06736 11074 237 5919 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06735 11074 237 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06734 11024 237 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06733 11074 489 490 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06732 2133 490 488 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06731 11074 490 2133 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06730 11074 490 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06729 11024 490 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06728 11074 238 236 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06727 489 236 105 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06726 11074 236 489 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06725 11074 236 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06724 11024 236 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06723 11074 2697 2437 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06722 10888 2437 2281 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06721 11074 2437 10888 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06720 11074 2437 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06719 11024 2437 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06718 11074 2697 2698 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06717 6132 2698 2696 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06716 11074 2698 6132 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06715 11074 2698 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06714 11024 2698 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06713 11074 2450 2438 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06712 2697 2438 2282 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06711 11074 2438 2697 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06710 11074 2438 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06709 11024 2438 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06708 11074 7721 3990 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06707 3991 5719 3992 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06706 4654 3992 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06705 1835 1837 1679 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06704 1679 1834 1835 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06703 11074 2688 1679 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06702 5528 1835 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06701 8483 8617 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06700 8619 8834 8484 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06699 11074 8616 8619 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06698 8824 8619 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06697 5820 5818 5819 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06696 5819 9379 5820 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06695 11074 10684 5819 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06694 6498 5820 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06693 3315 5599 3314 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06692 3316 9308 3315 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06691 3318 3969 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06690 3693 3315 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06689 11074 3974 3317 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06688 3316 3967 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06687 10312 9955 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06686 10231 9633 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06685 11074 11072 9071 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06684 9072 10701 9075 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06683 9095 9075 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06682 3593 6278 3592 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06681 3594 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06680 3596 5911 3595 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06679 4047 3741 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06678 3741 3604 3596 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06677 1725 2741 1724 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06676 1726 6243 1872 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06675 11074 2728 1723 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06674 1871 1872 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06673 468 1545 467 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06672 469 472 470 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06671 11074 5837 465 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06670 466 470 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06669 2611 8821 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06668 2613 10545 2612 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06667 11074 2609 2613 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06666 2610 2613 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06665 3471 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06664 4286 3879 3472 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06663 3470 4290 4286 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06662 11074 5124 3470 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06661 3470 4285 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06660 363 365 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06659 361 366 364 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06658 359 367 358 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06657 11074 706 359 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06656 11074 2673 367 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06655 366 367 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06654 11074 368 365 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06653 364 367 363 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06652 357 364 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06651 11074 360 362 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06650 358 366 360 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06649 706 358 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06648 11074 358 706 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06647 5457 5591 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06646 5456 5592 5589 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06645 5453 5594 5586 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06644 11074 6163 5453 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06643 11074 8048 5594 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06642 5592 5594 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06641 11074 6164 5591 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06640 5589 5594 5457 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06639 5454 5589 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06638 11074 5587 5455 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06637 5586 5592 5587 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06636 6163 5586 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06635 11074 5586 6163 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06634 5962 6203 6117 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06633 11074 6993 5963 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06632 5965 6413 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06631 6117 6204 5964 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06630 5966 6413 6203 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06629 6204 6993 5961 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06628 1180 9020 1179 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06627 1181 5600 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06626 1178 5918 1177 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06625 1574 1305 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06624 1305 1176 1178 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06623 10024 9612 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06622 5464 7514 5463 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06621 5467 7478 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06620 5466 9597 5465 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06619 6574 5596 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06618 5596 5462 5466 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06617 5166 6803 5167 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06616 5167 7437 5166 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06615 11074 8937 5167 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06614 5165 5166 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06613 3614 3612 3434 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06612 3434 4501 3614 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06611 11074 3610 3434 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06610 3611 3614 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06609 529 686 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06608 527 687 684 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06607 526 688 680 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06606 11074 691 526 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06605 11074 2673 688 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06604 687 688 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06603 11074 690 686 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06602 684 688 529 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06601 525 684 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06600 11074 683 528 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06599 680 687 683 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06598 691 680 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06597 11074 680 691 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06596 10478 10659 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06595 10477 10660 10658 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06594 10475 10661 10654 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06593 11074 10652 10475 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06592 11074 11051 10661 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06591 10660 10661 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06590 11074 10680 10659 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06589 10658 10661 10478 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06588 10476 10658 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06587 11074 10655 10479 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06586 10654 10660 10655 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06585 10652 10654 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06584 11074 10654 10652 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06583 2558 5746 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06582 2717 2693 2559 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06581 5895 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06580 5897 6861 5896 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06579 5894 6574 5897 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06578 11074 7840 5894 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06577 5894 9424 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_06576 10484 10670 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06575 10482 10671 10666 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06574 10480 10672 10663 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06573 11074 10662 10480 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06572 11074 11051 10672 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06571 10671 10672 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06570 11074 10668 10670 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06569 10666 10672 10484 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06568 10481 10666 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06567 11074 10665 10483 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06566 10663 10671 10665 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06565 10662 10663 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06564 11074 10663 10662 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06563 3426 8824 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06562 8309 8817 3427 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06561 3525 3693 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06560 3694 8297 3526 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06559 10256 3413 479 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06558 11074 2473 481 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06557 480 481 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06556 1706 2119 1707 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06555 1708 1866 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06554 2688 1864 1706 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06553 4559 5140 4564 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06552 11074 4554 4555 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06551 11074 5140 4566 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06550 4562 4617 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06549 4563 4561 4562 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06548 4560 4553 4559 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06547 4555 4554 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06546 519 668 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06545 516 669 666 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06544 515 670 663 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06543 11074 4254 515 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06542 11074 5083 670 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06541 669 670 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06540 11074 2610 668 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06539 666 670 519 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06538 517 666 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06537 11074 664 518 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06536 663 669 664 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06535 4254 663 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06534 11074 663 4254 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06533 11074 10018 9578 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06532 9580 9594 9581 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06531 9579 9581 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06530 10827 10959 10829 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06529 11074 10826 10824 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06528 11074 10959 10833 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06527 10830 10847 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06526 10831 10835 10830 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06525 10828 10825 10827 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06524 10824 10826 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06523 10856 10959 10855 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06522 11074 10852 10853 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06521 11074 10959 10858 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06520 10859 10877 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06519 10860 10864 10859 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06518 10857 10854 10856 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06517 10853 10852 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06516 10883 10959 10881 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06515 11074 10878 10879 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06514 11074 10959 10885 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06513 10886 10917 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06512 10882 10887 10886 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06511 10884 10880 10883 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06510 10879 10878 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06509 10949 10959 10946 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06508 11074 10943 10944 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06507 11074 10959 10952 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06506 10947 10951 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06505 10948 10953 10947 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06504 10950 10945 10949 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06503 10944 10943 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06502 10926 10959 10925 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06501 11074 10922 10923 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06500 11074 10959 10928 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06499 10929 10977 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06498 10930 10931 10929 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06497 10927 10924 10926 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06496 10923 10922 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06495 10282 10959 10281 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06494 11074 10280 10646 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06493 11074 10959 10287 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06492 10285 11012 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06491 10286 10284 10285 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06490 10283 10641 10282 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06489 10646 10280 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06488 827 5086 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06487 4240 1401 828 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06486 6451 6468 6336 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06485 11074 9987 6338 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06484 6337 6338 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06483 756 2473 643 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06482 11074 3413 757 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06481 644 757 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06480 11074 3391 2781 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06479 2778 2781 2777 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06478 11074 2776 2778 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06477 3069 2777 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06476 11074 2777 3069 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06475 2873 3037 2871 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06474 2872 3036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06473 3959 3035 2873 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06472 11074 4926 2808 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06471 2809 3830 2972 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06470 2971 2972 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06469 5970 7711 5969 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06468 5971 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06467 5967 9597 5972 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06466 6215 8848 5968 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06465 3156 5144 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06464 3158 3155 3157 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06463 9130 9296 9129 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06462 9131 9298 9299 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06461 11074 9297 9132 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06460 9295 9299 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06459 10957 10959 10955 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06458 11074 10954 10970 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06457 11074 10959 10960 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06456 10961 11039 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06455 10956 10962 10961 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06454 10958 10963 10957 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06453 10970 10954 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06452 7794 10689 7799 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06451 7800 11066 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06450 7796 10399 7795 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06449 7798 9716 7797 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06448 1137 1552 1136 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06447 1140 5809 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06446 1139 7041 1138 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06445 1867 1299 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06444 1299 1135 1139 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06443 5429 6275 5432 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06442 5433 10029 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06441 5431 7478 5430 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06440 5816 5563 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06439 5563 5428 5431 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06438 11074 5528 5530 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06437 5382 5530 5529 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06436 11074 6437 5382 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06435 5527 5529 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06434 11074 5529 5527 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06433 8828 8833 8827 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06432 8832 8831 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06431 8830 8824 8829 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06430 10541 8826 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06429 8826 8825 8830 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06428 8267 9566 7873 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06427 7873 8644 8267 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06426 11074 8081 7872 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06425 11074 9605 6999 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06424 7001 6998 7000 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06423 6997 7000 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06422 11074 3092 240 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06421 107 240 239 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06420 11074 8124 107 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06419 238 239 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06418 11074 239 238 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06417 10511 10710 10513 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06416 10514 10709 10711 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06415 11074 10708 10512 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06414 11067 10711 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06413 11074 2432 2277 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06412 2278 7701 2433 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06411 3008 2433 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06410 11074 2038 1672 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06409 1671 7701 1829 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06408 2691 1829 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06407 5695 5701 5698 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06406 11074 5693 5696 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06405 5699 6201 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06404 5698 5694 5697 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06403 5700 6201 5701 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06402 5694 5693 5692 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06401 11074 5665 5666 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06400 5668 5670 5669 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06399 5667 5669 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06398 11074 6493 4697 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06397 4699 5607 4698 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06396 4694 4698 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06395 3994 5918 3546 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06394 3546 5911 3994 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06393 11074 4654 3545 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06392 7433 9552 7255 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06391 7255 7437 7433 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06390 11074 9300 7255 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06389 7432 7433 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06388 2270 2423 6192 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06387 11074 9305 2271 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06386 2273 6105 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06385 6192 2424 2272 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06384 2274 6105 2423 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06383 2424 9305 2269 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06382 9251 10698 9250 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06381 9253 10078 9425 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06380 11074 10708 9252 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06379 9430 9425 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06378 5299 6179 5298 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06377 5300 5302 5305 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06376 11074 5908 5301 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06375 5295 5305 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06374 4725 4727 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06373 4482 4728 4484 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06372 4479 4729 4724 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06371 11074 8124 4479 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06370 11074 5262 4729 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06369 4728 4729 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06368 11074 4726 4727 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06367 4484 4729 4725 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06366 4480 4484 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06365 11074 4481 4483 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06364 4724 4728 4481 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06363 8124 4724 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06362 11074 4724 8124 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06361 11074 10774 7579 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06360 7578 7579 7580 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06359 11074 10567 7578 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06358 10172 7580 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06357 11074 7580 10172 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06356 6526 8762 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06355 6525 6866 6526 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06354 11074 6524 6525 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06353 10030 10608 9817 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06352 9817 10606 10030 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06351 11074 10945 9817 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06350 9932 10030 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06349 2923 3077 2922 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06348 2924 3076 3078 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06347 11074 4349 2925 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06346 4057 3078 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06345 1588 9020 1590 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06344 1589 5600 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06343 1585 9308 1587 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06342 1583 1586 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06341 1586 1584 1585 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06340 6568 9716 6567 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06339 6566 10704 6565 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06338 11074 9747 6563 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06337 6564 6565 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06336 441 452 445 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06335 446 464 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06334 443 745 442 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06333 7701 444 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06332 444 440 443 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06331 3927 4602 3926 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06330 3926 4142 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06329 3925 3926 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06328 7138 7141 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06327 7137 7140 7139 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06326 7133 7143 7132 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06325 11074 7516 7133 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06324 11074 8048 7143 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06323 7140 7143 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06322 11074 7521 7141 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06321 7139 7143 7138 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06320 7134 7139 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06319 11074 7136 7135 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06318 7132 7140 7136 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06317 7516 7132 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06316 11074 7132 7516 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06315 2358 7478 2357 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06314 2359 5599 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06313 2361 8126 2360 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06312 2601 2503 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06311 2503 2356 2361 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06310 43 174 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06309 42 175 173 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06308 40 176 169 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06307 11074 708 40 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06306 11074 2673 176 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06305 175 176 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06304 11074 377 174 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06303 173 176 43 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06302 41 173 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06301 11074 170 44 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06300 169 175 170 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06299 708 169 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06298 11074 169 708 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06297 7326 7495 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06296 7323 7496 7494 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06295 7322 7497 7490 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06294 11074 7749 7322 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06293 11074 10638 7497 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06292 7496 7497 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06291 11074 7752 7495 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06290 7494 7497 7326 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06289 7324 7494 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06288 11074 7492 7325 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06287 7490 7496 7492 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06286 7749 7490 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06285 11074 7490 7749 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06284 5082 5081 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06283 5077 5085 5080 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06282 5074 5084 5075 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06281 11074 5488 5074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06280 11074 5083 5084 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06279 5085 5084 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06278 11074 5487 5081 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06277 5080 5084 5082 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06276 5078 5080 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06275 11074 5076 5079 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06274 5075 5085 5076 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06273 5488 5075 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06272 11074 5075 5488 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06271 6349 6497 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06270 11019 6499 6350 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06269 8573 10687 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06268 8749 8748 8574 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06267 7811 9083 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06266 7813 9080 7812 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06265 4879 5321 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06264 5040 5934 4878 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06263 10433 10558 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06262 10556 10560 10434 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06261 11074 10561 10556 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06260 10808 10556 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06259 5565 6545 5434 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06258 11074 8409 5566 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06257 5435 5566 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06256 2847 4617 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06255 4410 4553 2848 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06254 8924 8922 8923 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06253 8925 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06252 8919 8921 8926 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06251 10013 8918 8920 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06250 1522 7721 1523 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06249 1524 7711 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06248 1865 1862 1522 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06247 9218 9972 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06246 9411 9409 9217 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06245 7969 10687 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06244 8046 8407 7970 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06243 6361 8733 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06242 7142 6867 6362 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06241 565 1248 564 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06240 11074 721 722 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06239 11074 1248 569 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06238 567 5531 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06237 568 653 567 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06236 566 711 565 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06235 722 721 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06234 3552 8922 3550 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06233 3551 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06232 8709 5898 3552 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06231 10168 11075 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06230 10170 11072 10169 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06229 6101 8244 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06228 6182 6574 6100 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06227 11074 2788 2592 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06226 2592 2495 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06225 2321 3079 2592 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06224 7043 7041 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06223 8635 7042 7044 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06222 1641 7426 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06221 2974 1810 1642 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06220 3269 3274 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06219 3268 3273 3270 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06218 3264 3275 3267 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06217 11074 8305 3264 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06216 11074 5083 3275 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06215 3273 3275 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_06214 11074 3272 3274 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_06213 3270 3275 3269 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06212 3265 3270 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06211 11074 3266 3271 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06210 3267 3273 3266 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06209 8305 3267 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06208 11074 3267 8305 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06207 9771 10566 9770 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06206 9772 10218 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06205 9768 10542 9767 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06204 10184 10541 9769 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06203 9995 10583 9778 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06202 9778 10564 9995 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06201 11074 10565 9778 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06200 9991 9995 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06199 5383 5736 5385 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06198 11074 5534 5531 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06197 11074 5736 5388 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06196 5386 6449 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06195 5387 5536 5386 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06194 5384 10680 5383 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06193 5531 5534 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06192 58 1248 59 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06191 11074 198 195 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06190 11074 1248 60 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06189 56 3277 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06188 57 199 56 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06187 55 724 58 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06186 195 198 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06185 6207 6210 6081 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06184 6082 10258 6207 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06183 6083 6451 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06182 6121 6207 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06181 11074 10256 6080 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06180 6082 10269 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06179 4811 5583 4812 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06178 4813 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06177 6230 5599 4811 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06176 10259 10268 10144 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06175 11074 10774 10146 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06174 10145 10146 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06173 4840 7711 4839 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06172 4841 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06171 4843 8921 4842 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06170 4998 5293 4838 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06169 4848 9309 4847 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06168 4849 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06167 4845 9560 4850 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06166 5001 8921 4846 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06165 5306 6177 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06164 5304 5926 5303 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06163 4464 5897 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06162 4463 6171 4462 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06161 11074 7484 3527 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06160 3528 3695 3696 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06159 3958 3696 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06158 11074 5718 3880 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06157 3878 5153 3883 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06156 3879 3883 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06155 11074 4311 4127 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06154 4128 6811 4313 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06153 4312 4313 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06152 11074 4410 3495 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06151 3496 3928 3663 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06150 3905 3663 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06149 8232 9418 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06148 8431 9417 8233 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06147 961 1284 965 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06146 11074 960 963 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06145 11074 1284 968 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06144 966 5707 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06143 967 964 966 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06142 962 959 961 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06141 963 960 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06140 589 1284 587 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06139 11074 742 743 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06138 11074 1284 591 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06137 592 5732 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06136 588 656 592 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06135 590 729 589 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06134 743 742 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06133 378 1284 380 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06132 11074 383 377 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06131 11074 1284 384 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06130 381 5531 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06129 382 385 381 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06128 379 708 378 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06127 377 383 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06126 417 1284 420 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06125 11074 423 419 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06124 11074 1284 424 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06123 421 3277 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06122 422 425 421 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06121 418 726 417 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06120 419 423 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06119 3281 7042 3278 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06118 11074 3276 3277 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06117 11074 7042 3283 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06116 3279 10995 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06115 3280 3284 3279 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06114 3282 8297 3281 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06113 3277 3276 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06112 1539 7042 1538 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06111 1540 6243 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06110 1535 2741 1541 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06109 1537 1881 1536 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06108 7031 10604 7018 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06107 7018 8091 7031 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06106 11074 8930 7017 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06105 2920 4029 2918 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06104 2919 3070 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06103 4036 3370 2920 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06102 2415 2435 2033 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06101 2033 2434 2415 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06100 11074 4325 2031 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06099 8514 10031 8513 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06098 8515 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06097 8511 8643 8516 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06096 9526 8642 8512 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06095 5363 5727 5362 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06094 5364 5728 5520 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06093 11074 10024 5361 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06092 5519 5520 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06091 7273 7455 7276 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06090 7274 7459 7456 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06089 11074 7672 7275 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06088 8095 7456 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06087 6094 6251 6093 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06086 6095 6232 6231 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06085 11074 6230 6092 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06084 8644 6231 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_06083 896 1248 894 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06082 11074 891 892 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06081 11074 1248 898 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06080 899 4910 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06079 895 893 899 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06078 897 902 896 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06077 892 891 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06076 4528 5736 4527 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06075 11074 4913 4910 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06074 11074 5736 4534 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06073 4531 6401 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06072 4529 4914 4531 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06071 4525 10257 4528 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_06070 4910 4913 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06069 9503 9514 9501 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06068 11074 10774 9504 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06067 9502 9504 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06066 5796 7721 5795 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06065 5797 6277 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06064 5793 8643 5792 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06063 6206 5794 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06062 5794 5791 5793 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06061 10695 10693 10495 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06060 10495 10694 10695 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06059 11074 10706 10494 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06058 5337 7484 5336 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06057 5338 8885 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06056 5340 8122 5339 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06055 5500 7655 5341 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06054 11074 6142 5767 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06053 5768 7045 5769 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06052 5766 5769 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06051 4132 4323 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06050 4321 5539 4133 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06049 11074 6213 4321 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06048 4322 4321 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06047 7631 8082 7256 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06046 11074 10915 7435 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06045 7257 7435 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06044 9713 10701 9715 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06043 9714 10694 9713 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06042 9712 10686 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06041 9710 9713 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06040 11074 10702 9711 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06039 9714 9971 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_06038 11074 9305 7227 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06037 7228 7414 7409 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06036 7408 7409 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06035 4340 4348 4179 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06034 4179 4347 4340 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06033 11074 6503 4179 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06032 4450 4340 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06031 5005 5601 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06030 11074 5008 5005 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06029 5005 5002 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06028 11074 5009 5005 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06027 5024 5005 4851 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06026 11074 1456 1457 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06025 1458 7701 1459 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06024 2434 1459 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06023 11074 1403 1404 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06022 1405 7701 1406 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06021 2004 1406 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06020 7741 10027 7747 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06019 7743 10027 7748 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06018 7744 8709 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06017 7746 7748 7745 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06016 11074 8708 7742 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06015 9705 10705 9704 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06014 9706 10378 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06013 9708 11076 9707 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06012 9702 9709 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_06011 9709 9703 9708 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_06010 11074 6243 2902 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06009 2902 3714 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06008 3064 3056 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06007 2902 10018 3056 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06006 3056 4014 2902 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_06005 8996 9005 9002 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06004 11074 8995 8997 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06003 9000 8999 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06002 9002 8998 9001 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_06001 9003 8999 9005 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_06000 8998 8995 8994 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05999 11074 6220 3948 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05998 3949 6221 3950 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05997 5771 3950 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05996 3011 3008 2850 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05995 2850 3009 3011 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05994 11074 6132 2849 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05993 748 2472 601 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05992 601 10256 748 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05991 11074 8713 601 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05990 752 748 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05989 3956 10596 3957 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05988 3957 10595 3956 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05987 11074 10995 3955 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05986 10243 10896 10242 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05985 10244 10258 10243 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05984 10245 10913 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05983 10239 10243 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05982 11074 10256 10246 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05981 10244 10269 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05980 2130 9020 2129 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05979 2131 2133 2134 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05978 11074 5918 2132 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05977 5736 2134 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05976 2252 3193 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05975 2401 3626 2252 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05974 11074 3632 2401 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05973 5753 6803 5754 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05972 5754 7437 5753 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05971 11074 8937 5752 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05970 7608 7606 7607 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05969 7607 7690 7608 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05968 11074 9275 7607 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05967 7605 7608 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05966 2605 7711 2604 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05965 2606 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05964 2608 5599 2607 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05963 2801 2800 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05962 2800 2603 2608 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05961 11018 10366 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05960 10594 9509 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05959 6714 8746 6718 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05958 6715 8059 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05957 6717 8453 6716 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05956 6896 6897 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05955 6897 6713 6717 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05954 7842 9433 7841 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05953 7843 9426 7845 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05952 11074 9716 7844 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05951 7840 7845 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05950 342 1495 346 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05949 346 1494 343 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05948 344 348 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05947 339 338 346 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05946 11074 1489 340 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05945 11074 341 345 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05944 2418 346 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05943 2878 3322 2877 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05942 2879 3311 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05941 2881 3306 2880 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05940 3285 3039 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05939 3039 2876 2881 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05938 5691 5698 5690 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05937 5690 6119 5691 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05936 11074 5703 5690 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05935 6195 5691 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05934 49 183 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05933 47 184 180 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05932 45 185 177 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05931 11074 723 45 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05930 11074 2446 185 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05929 184 185 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05928 11074 397 183 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05927 180 185 49 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05926 46 180 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05925 11074 179 48 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05924 177 184 179 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05923 723 177 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05922 11074 177 723 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05921 6032 6264 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05920 6030 6265 6263 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05919 6029 6266 6260 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05918 11074 6261 6029 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05917 11074 8048 6266 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05916 6265 6266 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05915 11074 6538 6264 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05914 6263 6266 6032 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05913 6028 6263 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05912 11074 6262 6031 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05911 6260 6265 6262 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05910 6261 6260 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05909 11074 6260 6261 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05908 10241 10596 10240 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05907 10240 10595 10241 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05906 11074 10257 10240 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05905 10585 10241 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05904 2073 5557 2072 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05903 2072 2452 2073 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05902 11074 5766 2071 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05901 3512 3941 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05900 3922 3938 3511 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05899 1001 1003 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05898 844 1002 997 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05897 841 1004 992 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05896 11074 1490 841 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05895 11074 2446 1004 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05894 1002 1004 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05893 11074 1265 1003 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05892 997 1004 1001 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05891 842 997 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05890 11074 998 843 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05889 992 1002 998 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05888 1490 992 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05887 11074 992 1490 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05886 10037 10596 9819 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05885 9819 10595 10037 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05884 11074 11018 9819 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05883 10032 10037 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05882 2036 7027 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05881 2081 2035 2037 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05880 4431 6276 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05879 10269 9560 4432 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05878 10081 5556 5415 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05877 5415 5557 10081 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05876 11074 5776 5414 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05875 8939 10908 8940 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05874 8940 9347 8939 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05873 11074 8938 8940 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05872 8937 8939 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05871 3497 3928 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05870 3668 4410 3498 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05869 10464 10628 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05868 10463 10629 10627 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05867 10460 10630 10623 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05866 11074 10909 10460 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05865 11074 10914 10630 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05864 10629 10630 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05863 11074 10995 10628 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05862 10627 10630 10464 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05861 10461 10627 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05860 11074 10624 10462 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05859 10623 10629 10624 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05858 10909 10623 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05857 11074 10623 10909 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05856 11 124 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05855 8 125 123 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05854 7 126 119 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05853 11074 8839 7 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05852 11074 2673 126 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05851 125 126 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05850 11074 4885 124 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05849 123 126 11 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05848 9 123 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05847 11074 121 10 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05846 119 125 121 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05845 8839 119 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05844 11074 119 8839 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05843 4619 10915 4618 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05842 11074 4961 4969 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05841 11074 10915 4625 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05840 4626 5191 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05839 4620 4964 4626 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05838 4616 6465 4619 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05837 4969 4961 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05836 9724 9760 9723 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05835 9723 10694 9724 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05834 11074 10702 9722 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05833 8770 11076 8606 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05832 8606 10710 8770 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05831 11074 10686 8607 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05830 5297 6586 5296 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05829 5296 5292 5297 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05828 11074 5293 5294 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05827 572 1495 728 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05826 728 1494 574 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05825 575 726 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05824 570 723 728 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05823 11074 1489 571 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05822 11074 724 573 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05821 3009 728 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05820 9794 10027 9795 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05819 9796 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05818 10002 10880 9794 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05817 2731 6275 2732 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05816 2733 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05815 3037 4070 2731 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05814 9847 10058 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05813 9844 10060 10056 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05812 9843 10057 10053 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05811 11074 10054 9843 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05810 11074 11051 10057 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05809 10060 10057 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05808 11074 10059 10058 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05807 10056 10057 9847 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05806 9845 10056 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05805 11074 10055 9846 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05804 10053 10060 10055 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05803 10054 10053 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05802 11074 10053 10054 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05801 9113 9271 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05800 9112 9272 9270 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05799 9109 9273 9266 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05798 11074 10213 9109 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05797 11074 10914 9273 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05796 9272 9273 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05795 11074 10177 9271 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05794 9270 9273 9113 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05793 9110 9270 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05792 11074 9267 9111 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05791 9266 9272 9267 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05790 10213 9266 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05789 11074 9266 10213 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05788 2715 10959 2714 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05787 11074 3023 3272 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05786 11074 10959 2721 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05785 2716 3263 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05784 2710 3026 2716 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05783 2708 8305 2715 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05782 3272 3023 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05781 4091 10959 4090 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05780 11074 4269 4496 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05779 11074 10959 4093 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05778 4094 4240 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05777 4095 4242 4094 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05776 4092 7601 4091 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05775 4496 4269 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05774 4521 10959 4520 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05773 11074 4514 4892 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05772 11074 10959 4526 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05771 4522 4524 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05770 4523 4518 4522 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05769 4519 7418 4521 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05768 4892 4514 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05767 1657 10959 1656 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05766 11074 1819 1816 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05765 11074 10959 1658 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05764 1654 2003 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05763 1655 1820 1654 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05762 1653 7425 1657 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05761 1816 1819 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05760 2064 10959 2063 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05759 11074 2066 2062 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05758 11074 10959 2067 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05757 2068 2073 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05756 2069 2070 2068 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05755 2065 7450 2064 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05754 2062 2066 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05753 2021 10959 2020 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05752 11074 2023 2019 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05751 11074 10959 2025 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05750 2026 2024 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05749 2027 2028 2026 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05748 2022 7611 2021 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05747 2019 2023 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05746 6991 8122 6990 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05745 6989 6992 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05744 6998 7655 6991 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05743 1408 3832 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05742 4524 1409 1407 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05741 642 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05740 1042 7514 641 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05739 11074 4553 2660 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05738 2662 4617 2661 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05737 3632 2661 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05736 11074 4915 2626 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05735 2625 3817 2627 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05734 2965 2627 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05733 11074 6246 5173 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05732 5174 5181 5176 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05731 5175 5176 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05730 4752 5522 4751 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05729 4753 5521 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05728 4755 4959 4754 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05727 4916 4954 4750 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05726 3677 3945 3514 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05725 3514 3925 3677 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05724 11074 9987 3513 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05723 2712 10959 2711 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05722 11074 2707 2709 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05721 11074 10959 2722 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05720 2719 2717 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05719 2720 2718 2719 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05718 2713 7466 2712 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05717 2709 2707 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05716 2078 10959 2075 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05715 11074 2080 2074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05714 11074 10959 2082 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05713 2076 2081 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05712 2077 2083 2076 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05711 2079 7474 2078 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05710 2074 2080 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05709 2703 10959 2701 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05708 11074 2699 3019 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05707 11074 10959 2706 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05706 2705 3012 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05705 2702 2700 2705 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05704 2704 7037 2703 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05703 3019 2699 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05702 5423 6275 5422 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05701 5427 10029 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05700 5425 7478 5424 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05699 6483 8409 5426 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05698 5665 10604 4493 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05697 4493 8091 5665 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05696 11074 8642 4492 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05695 2035 2434 2034 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05694 2034 2435 2035 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05693 11074 10888 2032 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05692 4039 6173 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05691 4042 4183 4040 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05690 11074 2728 2302 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05689 2302 4014 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05688 4453 2476 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05687 2302 2572 2476 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05686 2476 3714 2302 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05685 4169 6275 4168 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05684 4170 5583 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05683 4981 7514 4169 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05682 1057 6275 1056 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05681 1058 6276 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05680 1542 1055 1057 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05679 2107 8922 2106 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05678 2108 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05677 2114 3703 2107 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05676 9888 10003 9887 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05675 9889 10002 10001 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05674 11074 10004 9890 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05673 10000 10001 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05672 4195 5718 4194 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05671 4196 5153 4289 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05670 11074 5131 4197 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05669 4288 4289 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05668 4199 6127 4198 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05667 4200 5159 4302 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05666 11074 5131 4201 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05665 4301 4302 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05664 1720 2109 1719 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05663 1721 1870 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05662 1717 1871 1722 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05661 2466 2114 1718 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05660 3333 3331 3332 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05659 3339 3338 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05658 3335 3709 3334 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05657 3337 3994 3336 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05656 9332 9333 9170 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05655 9170 9609 9332 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05654 11074 9603 9169 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05653 11074 2741 2154 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05652 2154 3714 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05651 3063 2153 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05650 2154 2578 2153 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05649 2153 4014 2154 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05648 3582 9309 3581 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05647 3583 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05646 3579 5719 3578 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05645 3739 5918 3580 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05644 7206 8453 7205 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05643 7207 8746 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05642 7202 8770 7208 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05641 7204 9433 7203 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05640 2591 3084 2787 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05639 2787 3082 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05638 2788 2787 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05637 5936 6286 5935 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05636 5935 6905 5936 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05635 11074 5933 5935 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05634 5934 5936 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05633 8878 8864 8868 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05632 8868 8865 8878 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05631 11074 8866 8867 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05630 9427 9980 9257 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05629 9257 9976 9427 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05628 11074 9426 9256 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05627 11074 4014 4006 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05626 11074 4348 4006 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05625 4006 4347 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05624 4005 4006 4004 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05623 8084 8318 7694 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05622 7694 8316 8084 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05621 11074 8970 7692 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05620 5721 5719 5720 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05619 5722 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05618 5716 10028 5723 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05617 5718 8869 5717 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05616 9912 10701 9911 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05615 9913 10078 10077 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05614 11074 10700 9914 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05613 11066 10077 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05612 5092 5093 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05611 11074 10604 5092 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05610 5092 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05609 11074 10888 5092 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05608 5091 5092 5090 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05607 11074 6108 5675 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05606 5676 6762 5677 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05605 5672 5677 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05604 11074 4012 2110 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05603 2111 2121 2112 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05602 2109 2112 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05601 11074 6275 3358 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05600 3360 3379 3359 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05599 3723 3359 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05598 11074 6277 2894 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05597 2895 9309 3048 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05596 3969 3048 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05595 11074 1396 1397 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05594 1398 7701 1399 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05593 2417 1399 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05592 9301 9955 9133 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05591 9133 9347 9301 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05590 11074 9559 9133 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05589 9300 9301 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05588 5550 10608 5407 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05587 5407 10606 5550 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05586 11074 8305 5406 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05585 7413 7411 7229 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05584 7229 7690 7413 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05583 11074 8000 7229 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05582 7410 7413 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05581 7454 7452 7270 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05580 7270 7690 7454 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05579 11074 10239 7270 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05578 7451 7454 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05577 11074 11072 7951 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05576 7952 11076 8159 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05575 8063 8159 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05574 84 1545 83 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05573 85 472 218 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05572 11074 4673 86 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05571 217 218 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05570 5126 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05569 5684 5523 5127 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05568 5125 5128 5684 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05567 11074 5124 5125 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05566 5125 5681 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_05565 8109 8113 7914 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05564 7914 8212 8109 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05563 11074 8112 7914 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05562 8340 8109 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05561 3081 3079 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05560 11074 3355 3081 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05559 6743 6905 6742 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05558 6746 7217 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05557 6745 7212 6744 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05556 6904 6907 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05555 6907 6741 6745 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05554 9998 10614 9783 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05553 9783 10615 9998 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05552 11074 10312 9781 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05551 2954 3100 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05550 2953 3099 3096 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05549 2951 3101 3094 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05548 11074 3092 2951 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05547 11074 5262 3101 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05546 3099 3101 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05545 11074 4370 3100 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05544 3096 3101 2954 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05543 2952 3096 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05542 11074 3095 2955 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05541 3094 3099 3095 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05540 3092 3094 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05539 11074 3094 3092 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05538 7123 7127 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05537 7125 7126 7124 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05536 7118 7128 7119 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05535 11074 7117 7118 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05534 11074 8048 7128 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05533 7126 7128 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05532 11074 7518 7127 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05531 7124 7128 7123 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05530 7120 7124 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05529 11074 7122 7121 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05528 7119 7126 7122 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05527 7117 7119 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05526 11074 7119 7117 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05525 5928 7204 5930 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05524 5930 6286 5928 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05523 11074 5927 5930 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05522 5926 5928 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05521 2586 8124 2585 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05520 2587 3092 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05519 2584 4066 2588 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05518 3379 2786 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05517 2786 2583 2584 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05516 2782 2589 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05515 11074 2590 2782 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05514 1188 6276 1187 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05513 1191 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05512 1190 9020 1189 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05511 2212 1313 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05510 1313 1186 1190 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05509 4861 9309 4860 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05508 4862 5012 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05507 4859 9020 4858 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05506 5292 5013 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05505 5013 4857 4859 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05504 4309 4925 4124 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05503 4124 4318 4309 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05502 11074 4926 4124 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05501 4307 4309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05500 4491 4489 4490 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05499 4490 5496 4491 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05498 11074 6206 4490 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05497 4488 4491 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05496 65 206 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05495 63 207 203 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05494 62 208 200 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05493 11074 726 62 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05492 11074 5262 208 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05491 207 208 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05490 11074 419 206 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05489 203 208 65 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05488 61 203 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05487 11074 202 64 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05486 200 207 202 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05485 726 200 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05484 11074 200 726 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05483 604 1041 602 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05482 603 752 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05481 1287 759 604 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05480 2089 5727 2087 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05479 2088 2456 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05478 2090 2094 2089 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05477 2097 5727 2095 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05476 2096 2093 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05475 2098 2094 2097 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05474 4237 4368 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05473 4370 4369 4238 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05472 5777 5552 5409 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05471 5409 10606 5777 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05470 11074 8918 5408 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05469 1990 6978 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05468 5490 1991 1989 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05467 4214 4327 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05466 4628 8713 4215 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05465 6814 9610 6659 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05464 6659 7437 6814 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05463 11074 9346 6659 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05462 6811 6814 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05461 6674 6838 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05460 6671 6839 6837 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05459 6670 6840 6833 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05458 11074 7085 6670 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05457 11074 8048 6840 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05456 6839 6840 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05455 11074 7089 6838 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05454 6837 6840 6674 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05453 6672 6837 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05452 11074 6835 6673 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05451 6833 6839 6835 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05450 7085 6833 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05449 11074 6833 7085 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05448 2015 2016 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05447 2012 2017 2014 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05446 2010 2018 2009 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05445 11074 7611 2010 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05444 11074 2673 2018 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05443 2017 2018 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05442 11074 2019 2016 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05441 2014 2018 2015 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05440 2008 2014 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05439 11074 2011 2013 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05438 2009 2017 2011 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05437 7611 2009 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05436 11074 2009 7611 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05435 6405 6406 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05434 6321 6324 6323 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05433 6319 6407 6403 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05432 11074 6992 6319 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05431 11074 10914 6407 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05430 6324 6407 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05429 11074 6404 6406 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05428 6323 6407 6405 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05427 6318 6323 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05426 11074 6320 6322 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05425 6403 6324 6320 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05424 6992 6403 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05423 11074 6403 6992 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05422 10566 10583 10439 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05421 10439 10564 10566 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05420 11074 10565 10438 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05419 7445 7444 7264 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05418 7264 7463 7445 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05417 11074 7467 7263 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05416 10509 10707 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05415 11061 10704 10510 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05414 10492 10695 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05413 10692 10691 10493 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05412 9254 9427 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05411 10074 9424 9255 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05410 8563 10687 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05409 9044 9033 8562 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05408 5289 5307 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05407 5288 5897 5287 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05406 3646 5726 2837 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05405 2837 2997 3646 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05404 11074 3236 2836 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05403 4495 4498 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05402 4406 4497 4407 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05401 4402 4499 4494 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05400 11074 7601 4402 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05399 11074 5083 4499 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05398 4497 4499 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05397 11074 4496 4498 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05396 4407 4499 4495 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05395 4403 4407 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05394 11074 4405 4404 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05393 4494 4497 4405 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05392 7601 4494 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05391 11074 4494 7601 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05390 11074 10018 9568 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05389 9569 9603 9570 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05388 10014 9570 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05387 8531 10031 8530 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05386 8532 8661 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05385 8534 9597 8533 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05384 9572 8699 8535 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05383 8560 10687 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05382 9409 9395 8561 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05381 7378 8765 7376 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05380 7377 7531 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05379 7532 8762 7378 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05378 2144 7721 2142 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05377 2143 9560 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05376 2480 10028 2144 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05375 9262 10083 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05374 9747 11072 9263 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05373 8362 9350 8361 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05372 11074 8692 8989 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05371 11074 9350 8364 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05370 8365 8694 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05369 8359 8696 8365 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05368 8360 8691 8362 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05367 8989 8692 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05366 8988 9376 8987 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05365 11074 8984 8999 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05364 11074 9376 8992 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05363 8991 8989 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05362 8990 8993 8991 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05361 8986 8985 8988 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05360 8999 8984 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05359 4871 5033 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05358 5034 5606 4872 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05357 11074 8318 6812 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05356 6658 6812 6810 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05355 11074 10018 6658 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05354 6809 6810 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05353 11074 6810 6809 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05352 6656 7041 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05351 6807 7042 6657 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05350 11074 10772 6807 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05349 6806 6807 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05348 11074 4926 3186 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05347 3187 4274 3189 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05346 3188 3189 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05345 11074 4410 4119 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05344 4120 4555 4294 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05343 4932 4294 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05342 5158 5727 5157 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05341 5160 5728 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05340 5159 10680 5158 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05339 24 1248 26 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05338 11074 148 145 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05337 11074 1248 29 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05336 27 4905 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05335 28 149 27 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05334 25 341 24 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05333 145 148 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05332 9146 9560 9145 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05331 9147 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05330 9149 9308 9148 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05329 9541 10825 9143 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05328 1401 2004 1402 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05327 1402 2006 1401 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05326 11074 10888 1400 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05325 1050 5918 1049 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05324 1051 9020 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05323 2578 7478 1050 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05322 8152 10710 7945 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05321 7945 10083 8152 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05320 11074 11072 7944 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05319 7214 8746 7213 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05318 7215 8059 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05317 7210 8453 7209 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05316 7212 9107 7211 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05315 8958 9350 8957 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05314 11074 8953 8985 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05313 11074 9350 8961 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05312 8959 9335 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05311 8955 8960 8959 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05310 8956 8954 8958 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05309 8985 8953 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05308 5268 5593 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05307 5307 5271 5268 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05306 11074 5878 5307 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05305 2485 4014 2309 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05304 2309 2741 2485 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05303 11074 2487 2309 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05302 3068 2485 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05301 3321 5898 3319 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05300 3320 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05299 3322 4070 3321 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05298 2745 7514 2747 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05297 2748 5898 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05296 2746 8124 2745 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05295 10190 10546 10189 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05294 10191 10551 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05293 10187 10555 10192 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05292 10559 10547 10188 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05291 4513 5736 4512 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05290 11074 4908 4905 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05289 11074 5736 4517 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05288 4515 6106 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05287 4516 4909 4515 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05286 4509 10231 4513 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05285 4905 4908 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05284 8899 9560 8898 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05283 8900 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05282 8896 8921 8895 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05281 9306 10854 8897 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05280 4814 10031 4818 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05279 4819 5012 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05278 4816 9020 4815 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05277 4991 8643 4817 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05276 8887 9309 8886 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05275 8888 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05274 8890 9308 8889 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05273 9532 8885 8891 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05272 4644 7068 4643 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05271 4645 4981 4647 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05270 11074 4658 4646 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05269 4983 4647 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05268 11074 4929 2244 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05267 2242 2393 2243 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05266 2396 3844 2325 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_05265 2243 2394 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05264 2324 4929 2394 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_05263 3606 2398 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_05262 2251 2401 2245 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05261 2247 3844 2246 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05260 2249 2396 2248 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05259 2250 3626 2251 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_05258 5355 5517 5693 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05257 11074 5518 5353 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05256 5356 5684 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05255 5693 5515 5357 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05254 5358 5684 5517 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05253 5515 5518 5354 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05252 331 1248 330 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05251 11074 333 329 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05250 11074 1248 334 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05249 335 5510 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05248 336 337 335 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05247 332 692 331 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05246 329 333 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05245 6466 9987 9362 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05244 6346 9987 6469 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05243 6470 6468 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05242 6472 6469 6471 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05241 11074 6465 6467 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05240 11074 7655 7008 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05239 7009 7007 7010 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05238 7006 7010 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05237 11074 8970 7910 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05236 7911 8388 8104 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05235 8030 8104 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05234 11074 8084 7879 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05233 7880 8638 8083 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05232 8012 8083 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05231 10579 10578 10442 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05230 10442 10577 10579 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05229 11074 10800 10442 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05228 10576 10579 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05227 6980 8893 6979 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05226 6979 7437 6980 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05225 11074 7012 6979 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05224 6978 6980 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05223 301 308 1796 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05222 11074 2385 302 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05221 305 2630 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05220 1796 304 306 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05219 307 2630 308 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05218 304 2385 303 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05217 5503 8918 5344 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05216 11074 10915 5505 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05215 5345 5505 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05214 11074 4255 856 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05213 857 3152 858 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05212 3833 858 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05211 11074 6275 3574 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05210 3573 3735 3733 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05209 4030 3733 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05208 11074 3065 2313 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05207 2314 2782 2488 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05206 2492 2488 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05205 5162 8839 5161 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05204 11074 10915 5163 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05203 5164 5163 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05202 8253 8261 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05201 8251 8613 8250 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05200 11074 8624 8251 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05199 8252 8251 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05198 9293 8862 8863 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05197 8863 9295 9293 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05196 11074 9987 8861 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05195 6077 8122 6076 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05194 6078 7484 6189 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05193 11074 7655 6079 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05192 6105 6189 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05191 11074 10708 9050 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05190 9053 10698 9052 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05189 9051 9052 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05188 7994 10710 7996 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05187 7997 11076 8156 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05186 11074 10700 7995 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05185 8059 8156 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05184 11074 9716 7401 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05183 7402 10399 7541 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05182 9424 7541 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05181 1132 7514 1131 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05180 1133 5911 1298 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05179 11074 8124 1134 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05178 1520 1298 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05177 11074 2104 7673 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05176 7673 2105 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05175 2103 2102 7673 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05174 11074 8684 8542 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05173 8542 10606 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05172 8679 8680 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05171 8542 8690 8680 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05170 8680 8682 8542 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05169 7130 7786 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05168 7131 8053 7130 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05167 11074 7129 7131 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05166 10680 10323 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05165 10995 10908 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05164 5247 5911 5246 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05163 5248 9020 5249 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05162 11074 7721 5245 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05161 10606 5249 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_05160 5321 4047 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05159 11074 4048 5321 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05158 3725 7523 3570 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05157 3569 5901 3725 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05156 3568 6574 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05155 3721 3725 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05154 11074 3723 3567 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05153 3569 3722 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_05152 1548 2099 1547 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05151 1553 1552 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05150 1550 2121 1549 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05149 1545 1551 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_05148 1551 1546 1550 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05147 1106 1219 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05146 1105 1218 1216 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05145 1103 1220 1213 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05144 11074 1403 1103 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05143 11074 2673 1220 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05142 1218 1220 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05141 11074 1235 1219 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05140 1216 1220 1106 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05139 1104 1216 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05138 11074 1214 1107 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05137 1213 1218 1214 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05136 1403 1213 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05135 11074 1213 1403 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05134 10041 10608 9821 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05133 9821 10606 10041 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05132 11074 10963 9821 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05131 10043 10041 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05130 9688 10054 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05129 11074 449 439 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05128 439 451 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05127 1489 438 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05126 439 437 438 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05125 438 466 439 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05124 5705 6201 5706 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05123 5706 5704 5705 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05122 11074 5702 5706 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05121 5703 5705 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05120 4674 4676 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05119 4437 4675 4438 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05118 4433 4677 4672 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05117 11074 4673 4433 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05116 11074 5262 4677 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05115 4675 4677 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05114 11074 6525 4676 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05113 4438 4677 4674 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05112 4434 4438 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05111 11074 4436 4435 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05110 4672 4675 4436 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05109 4673 4672 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05108 11074 4672 4673 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05107 7271 8834 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05106 7455 7652 7272 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05105 4208 4323 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05104 4318 5539 4209 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05103 39 165 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05102 36 166 164 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05101 35 167 160 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05100 11074 951 35 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05099 11074 2673 167 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05098 166 167 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05097 11074 934 165 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05096 164 167 39 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05095 37 164 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05094 11074 162 38 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05093 160 166 162 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05092 951 160 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05091 11074 160 951 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05090 1383 1385 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05089 1381 1384 1382 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05088 1377 1386 1376 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05087 11074 8617 1377 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05086 11074 5083 1386 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05085 1384 1386 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05084 11074 8312 1385 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05083 1382 1386 1383 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05082 1378 1382 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05081 11074 1380 1379 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05080 1376 1384 1380 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05079 8617 1376 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05078 11074 1376 8617 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05077 7729 8708 7728 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05076 11074 7733 7727 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05075 11074 8708 7734 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05074 7731 8297 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05073 7732 7737 7731 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05072 7730 8408 7729 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05071 7727 7733 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05070 2851 6440 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05069 3012 3011 2852 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05068 3557 4335 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05067 3718 5293 3558 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05066 4202 5165 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05065 4306 4305 4203 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05064 9864 10068 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05063 9862 10064 10067 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05062 9861 10065 10063 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05061 11074 10350 9861 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05060 11074 11051 10065 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05059 10064 10065 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05058 11074 10348 10068 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05057 10067 10065 9864 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05056 9860 10067 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05055 11074 10066 9863 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05054 10063 10064 10066 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05053 10350 10063 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05052 11074 10063 10350 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05051 11074 1881 1525 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05050 1526 4981 1527 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05049 1868 1527 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05048 5864 10687 5867 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05047 11074 5870 5866 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05046 11074 10687 5871 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05045 5868 6571 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05044 5869 5872 5868 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05043 5865 5863 5864 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_05042 5866 5870 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05041 7003 7655 7002 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05040 7005 7007 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05039 7004 8930 7003 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05038 6584 10704 6582 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05037 6583 8770 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05036 6585 7852 6584 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05035 11074 9100 8473 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05034 8473 8475 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05033 8472 8474 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05032 8473 9974 8474 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05031 8474 8477 8473 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_05030 5405 8316 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05029 5770 5561 5405 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05028 11074 8318 5770 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05027 4148 7068 4146 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05026 4147 4981 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05025 5181 4658 4148 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05024 11074 7068 7070 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05023 7071 7069 7072 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05022 9347 7072 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05021 9481 9484 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05020 9480 9483 9482 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05019 9476 9485 9475 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05018 11074 9922 9476 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05017 11074 10914 9485 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05016 9483 9485 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_05015 11074 9916 9484 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_05014 9482 9485 9481 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05013 9477 9482 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05012 11074 9479 9478 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05011 9475 9483 9479 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_05010 9922 9475 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05009 11074 9475 9922 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05008 11074 10018 9587 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05007 9588 9613 9589 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05006 10249 9589 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05005 6943 8831 6944 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05004 6944 6942 6943 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05003 11074 10774 6944 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05002 6941 6943 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_05001 6748 9433 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_05000 6908 9716 6747 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04999 4833 10031 4832 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04998 4834 5253 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04997 4836 5918 4835 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04996 4996 8126 4837 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04995 5445 8661 5444 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04994 5446 5579 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04993 5442 6276 5447 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04992 5580 8643 5443 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04991 11074 2473 502 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04990 500 502 501 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04989 11074 3413 500 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04988 499 501 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04987 11074 501 499 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04986 11074 10018 3353 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04985 3353 3714 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04984 3349 3352 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04983 3353 6221 3352 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04982 3352 4014 3353 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04981 8650 8318 8319 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04980 8319 8316 8650 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04979 11074 9335 8317 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04978 11074 10212 10209 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04977 10208 10206 10207 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04976 10570 10207 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04975 5369 6277 5368 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04974 5370 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04973 5372 8643 5371 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04972 5522 9287 5373 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04971 2667 4291 2666 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04970 11074 2993 2996 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04969 11074 4291 2671 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04968 2668 4617 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04967 2669 2994 2668 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04966 2663 4553 2667 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04965 2996 2993 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04964 11074 10018 7870 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04963 7871 8080 8079 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04962 8009 8079 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04961 3985 4665 3984 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04960 3986 6221 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04959 3988 4666 3987 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04958 3983 7069 3989 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04957 6052 10687 6054 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04956 11074 6279 6273 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04955 11074 10687 6055 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04954 6050 9074 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04953 6051 6169 6050 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04952 6053 6493 6052 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04951 6273 6279 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04950 7518 9046 7349 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04949 7349 7525 7518 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04948 11074 7517 7348 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04947 11074 3413 493 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04946 492 493 491 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04945 11074 2473 492 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04944 494 491 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04943 11074 491 494 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04942 11074 5911 4149 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04941 4149 7678 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04940 10614 4329 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04939 4149 4653 4329 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04938 4329 4654 4149 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_04937 1143 1552 1147 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04936 1148 5809 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04935 1145 7041 1144 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04934 1300 2099 1146 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04933 9653 10684 9651 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04932 11074 9655 10073 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04931 11074 10684 9656 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04930 9657 10231 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04929 9652 9658 9657 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04928 9654 10289 9653 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04927 10073 9655 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04926 5772 6455 5773 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04925 5773 5771 5772 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04924 11074 5770 5773 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04923 5774 5772 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04922 3304 3306 3303 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04921 3305 3322 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04920 3301 5771 3300 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04919 7437 3302 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04918 3302 3299 3301 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04917 6623 6766 6622 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04916 6624 6765 6767 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04915 11074 7655 6625 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04914 6764 6767 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04913 5479 7514 5478 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04912 5480 7478 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04911 5482 9597 5481 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04910 6286 5607 5483 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04909 11074 5906 5907 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04908 5909 6176 5910 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04907 5908 5910 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04906 11074 6820 5992 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04905 5993 7430 6219 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04904 6140 6219 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04903 905 1495 911 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04902 911 1494 906 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04901 907 1423 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04900 904 901 911 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04899 11074 1489 900 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04898 11074 902 903 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04897 2006 911 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04896 2988 2986 2827 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04895 2827 3860 2988 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04894 11074 4553 2827 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04893 2985 2988 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04892 3007 2691 2687 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04891 2687 2692 3007 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04890 11074 2688 2686 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04889 4575 4577 4950 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04888 11074 4940 4576 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04887 4583 4943 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04886 4950 4578 4579 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04885 4420 4943 4577 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04884 4578 4940 4419 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04883 8627 8848 8491 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04882 11074 10197 8628 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04881 8490 8628 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04880 11074 7655 7234 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04879 7233 7415 7416 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04878 7421 7416 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04877 1753 9560 1752 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04876 1754 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04875 1751 6275 1750 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04874 1886 1887 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04873 1887 1786 1751 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04872 4444 7711 4443 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04871 4445 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04870 4447 8921 4446 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04869 4679 4678 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04868 4678 4442 4447 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04867 4649 9020 4648 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04866 4651 5600 4650 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04865 11074 5898 4652 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04864 5552 4650 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04863 4076 4080 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04862 4075 4079 4078 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04861 4071 4081 4074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04860 11074 4070 4071 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04859 11074 5262 4081 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04858 4079 4081 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04857 11074 4374 4080 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04856 4078 4081 4076 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04855 4072 4078 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04854 11074 4073 4077 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04853 4074 4079 4073 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04852 4070 4074 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04851 11074 4074 4070 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04850 11074 10915 661 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04849 514 661 660 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04848 11074 4254 514 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04847 2609 660 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04846 11074 660 2609 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04845 9328 10596 9168 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04844 9168 10595 9328 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04843 11074 10024 9168 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04842 9329 9328 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04841 4050 6171 4055 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04840 4056 4054 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04839 4052 4057 4051 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04838 4363 4053 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04837 4053 4049 4052 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04836 11074 3712 4000 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04835 4000 3982 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04834 3553 3710 4000 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04833 11074 4005 4344 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04832 4344 4000 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04831 4001 4451 4344 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04830 11074 5017 4366 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04829 4187 4366 4365 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04828 11074 4364 4187 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04827 4368 4365 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04826 11074 4365 4368 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04825 3385 3739 3389 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04824 3390 3738 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04823 3387 3396 3386 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04822 3382 3388 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04821 3388 3384 3387 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04820 9675 9677 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04819 9670 9676 9674 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04818 9668 9679 9669 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04817 11074 9667 9668 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04816 11074 11051 9679 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04815 9676 9679 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04814 11074 9682 9677 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04813 9674 9679 9675 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04812 9671 9674 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04811 11074 9673 9672 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04810 9669 9676 9673 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04809 9667 9669 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04808 11074 9669 9667 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04807 6805 6803 6655 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04806 6655 8644 6805 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04805 11074 7036 6655 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04804 7459 6805 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04803 2576 3046 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04802 11074 2752 2576 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04801 2576 2575 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04800 11074 3337 2576 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04799 3330 10028 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04798 3338 4654 3329 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04797 3328 5911 3338 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04796 11074 3698 3328 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04795 3326 3969 3338 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04794 11074 5918 3327 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04793 9348 10323 9176 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04792 9176 9347 9348 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04791 11074 9613 9176 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04790 9346 9348 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04789 2219 2223 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04788 2218 2222 2221 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04787 2214 2224 2217 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04786 11074 2473 2214 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04785 11074 5262 2224 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04784 2222 2224 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04783 11074 4063 2223 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04782 2221 2224 2219 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04781 2215 2221 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04780 11074 2216 2220 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04779 2217 2222 2216 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04778 2473 2217 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04777 11074 2217 2473 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04776 2287 2444 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04775 2285 2448 2442 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04774 2284 2447 2440 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04773 11074 7466 2284 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04772 11074 2446 2447 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04771 2448 2447 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04770 11074 2709 2444 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04769 2442 2447 2287 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04768 2283 2442 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04767 11074 2441 2286 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04766 2440 2448 2441 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04765 7466 2440 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04764 11074 2440 7466 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04763 3165 3167 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04762 3161 3168 3166 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04761 3159 3169 3160 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04760 11074 8642 3159 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04759 11074 5083 3169 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04758 3168 3169 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04757 11074 6370 3167 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04756 3166 3169 3165 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04755 3162 3166 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04754 11074 3164 3163 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04753 3160 3168 3164 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04752 8642 3160 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04751 11074 3160 8642 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04750 1054 2099 1053 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04749 1052 1061 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04748 1292 1556 1054 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04747 4659 7721 4660 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04746 4661 7711 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04745 4658 9597 4659 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04744 6284 6286 6075 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04743 6075 6902 6284 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04742 11074 6285 6075 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04741 6180 6284 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04740 5731 5727 5729 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04739 5730 5728 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04738 6214 10594 5731 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04737 1118 1504 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04736 1268 1489 1119 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04735 9627 9938 9629 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04734 9628 10258 9627 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04733 9626 9939 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04732 9624 9627 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04731 11074 10256 9625 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04730 9628 10269 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_04729 611 7721 609 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04728 610 5898 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04727 1556 7514 611 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04726 4440 4679 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04725 4439 9002 4441 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04724 11074 4956 4958 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04723 4782 4958 4957 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04722 11074 5177 4782 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04721 4955 4957 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04720 11074 4957 4955 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04719 7253 9922 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04718 7430 8635 7254 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04717 7252 8636 7430 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04716 11074 8869 7252 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04715 7250 9313 7430 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04714 11074 8633 7251 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04713 4737 4893 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04712 4736 4894 4890 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04711 4734 4895 4887 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04710 11074 7418 4734 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04709 11074 5083 4895 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04708 4894 4895 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04707 11074 4892 4893 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04706 4890 4895 4737 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04705 4735 4890 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04704 11074 4888 4738 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04703 4887 4894 4888 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04702 7418 4887 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04701 11074 4887 7418 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04700 9154 10031 9153 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04699 9155 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04698 9151 10028 9156 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04697 10008 9313 9152 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04696 11074 7670 7671 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04695 7674 7673 7675 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04694 7672 7675 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04693 7823 9412 7821 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04692 7822 11076 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04691 7824 10700 7823 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04690 3374 3379 3373 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04689 3372 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04688 3370 5911 3374 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04687 3392 4048 3393 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04686 3393 4047 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04685 3391 3393 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04684 2086 7042 2084 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04683 2085 3033 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04682 3032 2728 2086 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04681 9992 10772 9776 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04680 9776 10564 9992 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04679 11074 9994 9776 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04678 10182 9992 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04677 11074 4929 2811 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04676 2812 2974 2813 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04675 2977 3844 2820 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_04674 2813 2975 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04673 2810 4929 2975 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_04672 2973 2979 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_04671 2821 3179 2814 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04670 2816 3844 2815 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04669 2818 2977 2817 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04668 2819 3183 2821 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04667 11074 8709 6507 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04666 6502 10366 6508 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04665 6854 6861 6681 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_04664 6508 6852 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04663 6680 8709 6852 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_04662 6851 6857 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_04661 6519 7117 6512 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04660 6514 6861 6513 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04659 6516 6854 6515 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04658 6510 9605 6519 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_04657 5349 5736 5347 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04656 11074 5511 5510 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04655 11074 5736 5351 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04654 5352 7422 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04653 5348 5514 5352 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04652 5350 10312 5349 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04651 5510 5511 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04650 9562 9560 9561 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04649 9563 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04648 9557 9597 9564 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04647 9559 10880 9558 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04646 5678 6465 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04645 6210 9987 5679 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04644 5887 10029 5886 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04643 5888 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04642 5884 5918 5889 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04641 5890 7721 5885 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04640 6709 9433 6708 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04639 6710 9057 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04638 6712 8052 6711 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04637 6895 9716 6707 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04636 6575 6574 6580 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04635 6581 8770 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04634 6577 10704 6576 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04633 6579 9747 6578 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04632 5682 5689 6200 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04631 11074 5681 5683 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04630 5686 5684 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04629 6200 5685 5687 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04628 5688 5684 5689 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04627 5685 5681 5680 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04626 3887 5153 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04625 3886 5718 3885 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04624 11074 6213 3886 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04623 3884 3886 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04622 595 1248 593 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04621 11074 744 1025 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04620 11074 1248 597 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04619 598 5544 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04618 594 659 598 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04617 596 1496 595 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04616 1025 744 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04615 5399 7042 5401 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04614 11074 5547 5544 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04613 11074 7042 5404 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04612 5402 10024 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04611 5403 5548 5402 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04610 5400 8918 5399 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04609 5544 5547 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04608 948 1248 947 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04607 11074 1246 1244 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04606 11074 1248 954 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04605 949 5707 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04604 950 1250 949 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04603 945 1245 948 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04602 1244 1246 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04601 5710 5736 5708 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04600 11074 5712 5707 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04599 11074 5736 5713 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04598 5714 6117 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04597 5709 5715 5714 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04596 5711 10594 5710 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04595 5707 5712 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04594 11074 6131 5747 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04593 5745 8021 5750 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04592 5746 5750 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04591 7443 7444 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04590 11074 10604 7443 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04589 7443 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04588 11074 10888 7443 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04587 7439 7443 7262 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04586 9506 10774 9509 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04585 9510 10774 9513 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04584 9511 9514 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04583 9507 9513 9512 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04582 11074 9505 9508 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04581 2198 5600 2197 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04580 2199 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04579 2201 9560 2200 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04578 2203 9308 2202 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04577 5022 5286 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04576 11074 5288 5022 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04575 5022 5018 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04574 11074 5024 5022 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04573 5017 5022 4869 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04572 11074 3377 3378 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04571 11074 3721 3378 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04570 3378 3375 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04569 4064 3378 3376 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04568 10212 10614 10211 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04567 10211 10615 10212 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04566 11074 10257 10210 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04565 1097 1211 1210 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04564 11074 2967 1098 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04563 1100 2630 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04562 1210 1208 1101 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04561 1102 2630 1211 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04560 1208 2967 1099 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04559 11074 1310 1311 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04558 9314 1311 1184 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04557 11074 1311 9314 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04556 11074 1311 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04555 11024 1311 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04554 11074 1310 1070 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04553 8661 1070 1071 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04552 11074 1070 8661 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04551 11074 1070 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04550 11024 1070 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04549 11074 767 766 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04548 1310 766 623 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04547 11074 766 1310 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04546 11074 766 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04545 11024 766 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04544 11074 9987 8625 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04543 8489 8625 8626 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04542 11074 8623 8489 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04541 8624 8626 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04540 11074 8626 8624 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04539 11074 2473 1063 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04538 1062 3413 1064 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04537 3734 1064 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04536 6561 7825 6562 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04535 6562 6564 6561 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04534 11074 10027 6562 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04533 6560 6561 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04532 11074 6579 5280 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04531 5282 5279 5281 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04530 5283 5281 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04529 11074 10702 9870 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04528 9871 10694 10071 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04527 9974 10071 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04526 11074 5295 4876 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04525 4877 5309 5039 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04524 5038 5039 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04523 11074 8022 7649 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04522 7647 8277 7651 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04521 7648 7651 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04520 11074 10418 9434 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04519 9433 9434 9264 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04518 11074 9434 9433 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04517 11074 9434 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04516 11024 9434 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04515 11074 10418 9108 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04514 9107 9108 9106 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04513 11074 9108 9107 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04512 11074 9108 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04511 11024 9108 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04510 11074 10419 10420 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04509 10418 10420 10417 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04508 11074 10420 10418 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04507 11074 10420 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04506 11024 10420 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04505 9755 10698 9754 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04504 9756 10078 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04503 9758 10701 9757 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04502 10080 9753 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04501 9753 9752 9758 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04500 9738 10705 9737 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04499 9739 10414 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04498 9735 11076 9734 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04497 9732 9736 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04496 9736 9733 9735 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04495 3293 3694 3296 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04494 3297 5550 3298 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04493 11074 3292 3294 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04492 3295 3298 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04491 11074 8092 3977 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04490 3978 3976 3979 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04489 3993 3979 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04488 6491 6819 6492 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04487 6492 6489 6491 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04486 11074 6490 6492 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04485 7766 6491 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04484 631 5809 633 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04483 634 1035 751 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04482 11074 2578 632 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04481 750 751 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04480 7427 9305 7249 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04479 7249 7437 7427 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04478 11074 8882 7249 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04477 7426 7427 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04476 3367 3379 3366 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04475 3368 6278 3371 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04474 11074 5911 3369 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04473 3726 3371 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04472 9701 10350 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04471 11013 11028 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04470 10332 10999 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04469 7802 9046 7804 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04468 7804 7813 7802 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04467 11074 8046 7801 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04466 10675 10990 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04465 6889 6879 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04464 6358 6261 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04463 4680 5863 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04462 5837 4673 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04461 6864 7516 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04460 2493 2796 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04459 11074 2582 2493 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04458 2984 2986 2826 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04457 2826 3860 2984 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04456 11074 4553 2825 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04455 2845 5535 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04454 3242 3007 2846 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04453 4586 4925 4585 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04452 4585 4584 4586 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04451 11074 4926 4585 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04450 4942 4586 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04449 5144 5142 5145 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04448 5145 5143 5144 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04447 11074 10915 5141 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04446 5949 9379 6404 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04445 5951 9379 6194 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04444 5952 6195 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04443 5954 6194 5953 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04442 11074 6765 5950 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04441 1371 1369 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04440 1368 1372 1370 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04439 1364 1373 1363 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04438 11074 1396 1364 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04437 11074 5083 1373 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04436 1372 1373 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04435 11074 1388 1369 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04434 1370 1373 1371 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04433 1366 1370 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04432 11074 1365 1367 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04431 1363 1372 1365 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04430 1396 1363 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04429 11074 1363 1396 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04428 5260 5264 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04427 5257 5263 5261 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04426 5254 5265 5255 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04425 11074 5863 5254 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04424 11074 5262 5265 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04423 5263 5265 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04422 11074 5866 5264 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04421 5261 5265 5260 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04420 5258 5261 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04419 11074 5256 5259 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04418 5255 5263 5256 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04417 5863 5255 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04416 11074 5255 5863 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04415 9808 10027 9807 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04414 9809 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04413 10015 10945 9808 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04412 7391 10080 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04411 7538 10399 7390 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04410 1862 3413 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04409 10781 10786 10782 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04408 10782 10780 10781 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04407 11074 10777 10778 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04406 1996 2657 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04405 1998 2984 1997 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04404 11074 3632 1998 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04403 2406 1998 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04402 3891 4943 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04401 4295 3890 3892 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04400 1711 1865 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04399 2105 2114 1712 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04398 1141 1302 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04397 2104 6243 1142 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04396 2100 7069 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04395 2102 2099 2101 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04394 7676 10700 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04393 7685 10027 7677 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04392 1290 1288 1127 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04391 1127 1287 1290 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04390 11074 1500 1127 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04389 1501 1290 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04388 8329 8675 8332 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04387 11074 8677 8949 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04386 11074 8675 8333 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04385 8334 8679 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04384 8335 8678 8334 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04383 8330 8954 8329 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04382 8949 8677 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04381 6702 10687 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04380 6890 6889 6703 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04379 6705 7167 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04378 6894 8056 6706 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04377 1374 6387 1375 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04376 1375 7408 1374 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04375 11074 5500 1375 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04374 6394 1374 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04373 10592 10608 10448 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04372 10448 10606 10592 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04371 11074 10825 10448 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04370 10591 10592 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04369 3240 3893 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04368 3246 4410 3241 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04367 8246 8247 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04366 8193 8197 8196 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04365 8191 8248 8245 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04364 11074 8623 8191 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04363 11074 10914 8248 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04362 8197 8248 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04361 11074 8252 8247 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04360 8196 8248 8246 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04359 8194 8196 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04358 11074 8192 8195 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04357 8245 8197 8192 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04356 8623 8245 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04355 11074 8245 8623 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04354 11074 9927 9554 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04353 9555 9571 9556 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04352 10215 9556 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04351 8354 8709 8351 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04350 11074 8687 8684 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04349 11074 8709 8356 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04348 8352 10680 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04347 8353 8689 8352 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04346 8355 8685 8354 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04345 8684 8687 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04344 4429 4981 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04343 10608 7068 4430 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04342 1709 1874 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04341 3961 2109 1710 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04340 2909 3062 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04339 3728 3063 2910 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04338 11074 10018 9545 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04337 9544 9559 9546 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04336 10004 9546 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04335 11074 10774 10563 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04334 10437 10563 10562 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04333 11074 10800 10437 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04332 10561 10562 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04331 11074 10562 10561 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04330 9787 10027 9785 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04329 9786 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04328 9925 10825 9787 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04327 11037 11038 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04326 11033 11040 11035 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04325 11031 11041 11030 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04324 11074 11028 11031 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04323 11074 11051 11041 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04322 11040 11041 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04321 11074 11036 11038 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04320 11035 11041 11037 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04319 11029 11035 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04318 11074 11032 11034 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04317 11030 11040 11032 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04316 11028 11030 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04315 11074 11030 11028 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04314 5661 5662 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04313 5658 5663 5660 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04312 5656 5664 5655 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04311 11074 10567 5656 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04310 11074 10914 5664 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04309 5663 5664 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04308 11074 10186 5662 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04307 5660 5664 5661 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04306 5654 5660 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04305 11074 5657 5659 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04304 5655 5663 5657 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04303 10567 5655 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04302 11074 5655 10567 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04301 11074 10018 7235 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04300 7236 7419 7417 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04299 7585 7417 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04298 1293 2472 1033 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04297 1033 10256 1293 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04296 11074 8713 1032 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04295 6555 10687 6554 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04294 11074 6552 7154 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04293 11074 10687 6559 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04292 6557 10080 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04291 6558 6556 6557 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04290 6553 7147 6555 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04289 7154 6552 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04288 6549 10687 6548 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04287 11074 6542 6543 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04286 11074 10687 6551 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04285 6550 7165 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04284 6546 6544 6550 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04283 6547 6545 6549 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04282 6543 6542 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04281 6518 6861 6517 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04280 6517 7747 6518 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04279 11074 6862 6511 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04278 10388 10705 10393 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04277 10394 10414 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04276 10390 11076 10389 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04275 10392 10700 10391 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04274 8401 8403 8400 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04273 8396 8395 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04272 8398 8437 8397 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04271 8394 10704 8399 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04270 7230 8122 7231 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04269 7232 7484 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04268 7414 7655 7230 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04267 4255 10604 4084 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04266 4084 8091 4255 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04265 11074 8885 4083 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04264 9631 10684 9630 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04263 11074 9636 10078 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04262 11074 10684 9637 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04261 9634 9633 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04260 9635 9638 9634 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04259 9632 9945 9631 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04258 10078 9636 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04257 10311 10684 10310 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04256 11074 10303 10698 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04255 11074 10684 10315 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04254 10316 10312 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04253 10305 10304 10316 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04252 10306 10662 10311 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04251 10698 10303 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04250 7400 9432 7398 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04249 7399 8770 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04248 7540 7852 7400 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04247 4104 5119 4103 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04246 4105 5123 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04245 4107 4959 4106 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04244 4274 4954 4102 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04243 7591 7596 8103 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04242 11074 8893 7588 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04241 7592 7594 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04240 8103 7590 7593 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04239 7595 7594 7596 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04238 7590 8893 7589 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04237 7925 8643 7924 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04236 7926 8126 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04235 7922 8124 7921 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04234 8121 9987 7923 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04233 2740 9308 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04232 5207 3040 2737 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04231 2738 2736 5207 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04230 11074 5599 2738 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04229 2734 5898 5207 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04228 11074 3379 2735 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04227 9836 10684 9835 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04226 11074 10051 10709 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04225 11074 10684 9840 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04224 9838 9955 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04223 9839 9957 9838 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04222 9837 10302 9836 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_04221 10709 10051 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04220 5903 8922 5902 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04219 5904 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04218 5899 5898 5905 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04217 5927 7711 5900 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04216 9535 9532 9534 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04215 9536 9547 9538 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04214 11074 9533 9537 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04213 9996 9538 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04212 8612 8613 8481 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04211 8481 8615 8612 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04210 11074 8610 8480 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04209 11074 7176 7168 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04208 7166 7177 7169 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04207 7167 7169 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04206 11074 9083 9086 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04205 9084 11066 9085 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04204 9081 9085 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04203 11074 9395 7080 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04202 7081 7476 7083 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04201 7082 7083 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04200 10603 10772 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04199 11074 10604 10603 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04198 10603 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04197 11074 10888 10603 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04196 10861 10603 10451 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04195 3398 7478 3397 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04194 3399 5599 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04193 3394 8126 3400 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04192 3396 5607 3395 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04191 2928 7711 2927 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04190 2929 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04189 2931 5599 2930 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04188 3151 7478 2926 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04187 6435 9333 6436 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04186 6436 7437 6435 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04185 11074 9321 6434 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04184 9104 11076 8609 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04183 8609 10083 9104 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04182 11074 10708 8608 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04181 6638 6792 6788 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04180 11074 7004 6639 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04179 6640 6789 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04178 6788 6787 6641 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04177 6642 6789 6792 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04176 6787 7004 6637 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04175 11074 9560 2295 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04174 2296 6276 2461 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04173 2736 2461 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04172 1810 2417 1646 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04171 1646 2418 1810 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04170 11074 2688 1645 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04169 10613 10614 10456 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04168 10456 10615 10613 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04167 11074 10680 10455 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04166 7240 7424 7422 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04165 11074 9552 7241 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04164 7243 7421 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04163 7422 7420 7244 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04162 7245 7421 7424 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04161 7420 9552 7242 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04160 11074 6574 4024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04159 4025 7527 4026 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04158 4023 4026 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04157 11074 5293 3562 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04156 3563 4010 3720 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04155 3719 3720 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04154 1701 7042 1700 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04153 1702 3033 1859 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04152 11074 2728 1699 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04151 1864 1859 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04150 7760 8643 7764 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04149 7765 8126 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04148 7762 8124 7761 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04147 8403 7763 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04146 7763 7759 7762 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04145 8240 10701 8239 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04144 8243 10073 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04143 8242 9405 8241 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04142 8458 8457 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04141 8457 8238 8242 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04140 7308 8126 7307 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04139 7309 7478 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04138 7306 9308 7305 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04137 7476 7479 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04136 7479 7304 7306 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04135 5459 5600 5458 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04134 5460 8661 5595 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04133 11074 8643 5461 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04132 5593 5595 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04131 1773 3734 1772 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04130 1774 3735 1896 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04129 11074 5293 1775 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04128 2208 1896 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04127 7982 9412 7981 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04126 7983 11076 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04125 7980 10083 7984 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04124 8051 8149 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04123 8149 7979 7980 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04122 3174 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04121 3607 3175 3172 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04120 3173 3188 3607 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04119 11074 5124 3173 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04118 3173 3606 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_04117 6678 6848 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04116 6677 6849 6845 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04115 6675 6850 6842 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04114 11074 10684 6675 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04113 11074 8048 6850 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04112 6849 6850 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04111 11074 6847 6848 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04110 6845 6850 6678 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04109 6676 6845 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04108 11074 6843 6679 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04107 6842 6849 6843 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04106 10684 6842 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04105 11074 6842 10684 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04104 1577 8661 1581 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04103 1582 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04102 1579 6276 1578 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04101 1575 1580 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04100 1580 1576 1579 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04099 7361 9412 7364 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04098 7365 11076 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04097 7363 9405 7362 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04096 7527 7528 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_04095 7528 7360 7363 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04094 7300 8126 7302 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04093 7303 7478 7477 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04092 11074 10028 7301 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04091 8100 7477 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_04090 3357 6221 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04089 11074 3714 3357 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04088 3357 7041 3356 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04087 3354 4014 3357 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04086 10784 10783 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04085 10786 10915 10785 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04084 3230 3004 2842 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04083 2842 5743 3230 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04082 11074 3219 2841 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04081 4292 4925 4118 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04080 4118 4291 4292 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04079 11074 4926 4118 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04078 4290 4292 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04077 3601 3749 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04076 3600 3750 3748 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04075 3598 3751 3744 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04074 11074 4066 3598 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04073 11074 5262 3751 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04072 3750 3751 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04071 11074 4476 3749 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04070 3748 3751 3601 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04069 3599 3748 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04068 11074 3745 3602 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04067 3744 3750 3745 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04066 4066 3744 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04065 11074 3744 4066 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04064 9203 9389 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04063 9200 9391 9388 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04062 9199 9390 9384 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04061 11074 9382 9199 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04060 11074 11051 9390 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04059 9391 9390 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04058 11074 9394 9389 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04057 9388 9390 9203 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04056 9201 9388 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04055 11074 9385 9202 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04054 9384 9391 9385 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04053 9382 9384 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04052 11074 9384 9382 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04051 2464 2576 2298 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04050 2298 2469 2464 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04049 11074 4327 2297 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04048 8291 9313 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04047 11074 8699 8291 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04046 8291 8930 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04045 11074 8297 8291 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04044 8290 8885 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04043 11074 8642 8290 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04042 8290 9304 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04041 11074 8918 8290 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04040 555 1495 710 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04039 710 1494 556 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04038 558 708 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04037 553 706 710 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04036 11074 1489 554 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04035 11074 711 557 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04034 2435 710 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04033 4805 5240 4988 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04032 4988 8409 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04031 4986 4988 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04030 6485 6483 6484 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04029 6488 6487 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04028 6486 8691 6485 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04027 6505 10027 6509 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04026 6504 7498 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04025 6506 6503 6505 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04024 8599 11066 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04023 8765 9977 8599 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04022 11074 8768 8765 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04021 5674 5671 5673 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04020 5673 7690 5674 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04019 11074 6121 5673 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04018 5670 5674 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04017 8633 6867 5810 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04016 5810 5809 8633 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04015 11074 8092 5808 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_04014 11074 6376 4485 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04013 4487 4488 4486 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04012 5143 4486 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_04011 1693 1852 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04010 1692 1853 1851 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04009 1690 1854 1847 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04008 11074 7474 1690 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04007 11074 2446 1854 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04006 1853 1854 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_04005 11074 2074 1852 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_04004 1851 1854 1693 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04003 1691 1851 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04002 11074 1848 1694 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04001 1847 1853 1848 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_04000 7474 1847 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03999 11074 1847 7474 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03998 862 864 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03997 825 863 860 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03996 823 865 859 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03995 11074 8885 823 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03994 11074 5083 865 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03993 863 865 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03992 11074 867 864 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03991 860 865 862 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03990 824 860 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03989 11074 861 826 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03988 859 863 861 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03987 8885 859 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03986 11074 859 8885 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03985 6570 6585 6572 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03984 6573 8767 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03983 6571 6569 6570 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03982 1468 1504 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03981 1841 7701 1469 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03980 1543 1542 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03979 3710 4981 1544 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03978 3980 4665 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03977 3982 4658 3981 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03976 1419 1420 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03975 1417 1421 1418 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03974 1412 1422 1415 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03973 11074 7425 1412 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03972 11074 2673 1422 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03971 1421 1422 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03970 11074 1816 1420 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03969 1418 1422 1419 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03968 1413 1418 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03967 11074 1416 1414 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03966 1415 1421 1416 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03965 7425 1415 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03964 11074 1415 7425 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03963 11074 10018 9797 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03962 9798 10017 10016 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03961 10009 10016 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03960 11074 8915 8910 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03959 8911 8913 8914 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03958 8912 8914 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03957 2890 8709 2888 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03956 2889 3047 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03955 3046 4012 2890 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03954 2891 6277 2892 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03953 2893 5911 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03952 3047 3706 2891 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03951 2113 6243 2115 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03950 2116 2114 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03949 2575 2121 2113 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03948 1161 5911 1159 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03947 1160 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03946 1870 3092 1161 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03945 11074 8340 8345 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03944 8338 9335 8339 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03943 8346 10027 8211 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03942 8339 8337 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03941 8210 8340 8337 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_03940 9341 8336 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_03939 8349 8341 8342 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03938 8344 10027 8343 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03937 8348 8346 8347 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03936 8350 10231 8349 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03935 10497 10697 10496 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03934 10498 11066 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03933 11058 10699 10497 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03932 10507 11076 10506 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03931 10508 10705 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03930 10706 11072 10507 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03929 3561 3967 3559 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03928 3560 3719 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03927 3738 5918 3561 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03926 3531 6277 3529 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03925 3530 6276 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03924 4327 8643 3531 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03923 6175 6286 6066 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03922 6066 6902 6175 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03921 11074 6285 6063 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03920 11074 6127 4770 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03919 4771 5159 4946 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03918 4944 4946 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03917 8932 9309 8931 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03916 8933 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03915 8935 10028 8934 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03914 10247 8930 8936 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03913 11074 1520 1521 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03912 11074 1537 1521 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03911 1521 7082 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03910 1519 1521 1518 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03909 9599 10029 9598 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03908 9604 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03907 9601 9597 9600 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03906 9603 10945 9602 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03905 6727 9057 6726 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03904 6728 9080 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03903 6730 8770 6729 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03902 6902 9433 6725 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03901 5913 6278 5912 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03900 5914 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03899 5916 9020 5915 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03898 6282 5911 5917 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03897 6721 8746 6720 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03896 6722 9057 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03895 6724 8770 6723 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03894 6901 9433 6719 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03893 5156 5727 5154 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03892 5155 5728 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03891 5153 11018 5156 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03890 10133 10566 10132 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03889 10136 10218 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03888 10135 10542 10134 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03887 10547 10193 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03886 10193 10131 10135 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03885 11074 8746 6695 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03884 6696 10399 6878 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03883 6877 6878 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03882 9590 10029 9595 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03881 9596 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03880 9592 10028 9591 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03879 9594 10924 9593 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03878 2164 6220 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03877 11074 3714 2164 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03876 2164 7042 2162 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03875 2163 4014 2164 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03874 11074 2581 2779 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03873 11074 3716 2779 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03872 2779 2582 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03871 4037 2779 2780 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03870 3888 5153 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03869 3889 5718 3888 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03868 11074 6213 3889 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03867 5100 5098 5101 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03866 5101 6195 5100 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03865 11074 10915 5099 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03864 8270 8848 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03863 8269 8834 8268 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03862 11074 8267 8269 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03861 9298 8269 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03860 4632 6259 4633 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03859 4633 4983 4632 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03858 11074 5194 4633 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03857 4631 4632 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03856 11074 1075 1072 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03855 5600 1072 1073 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03854 11074 1072 5600 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03853 11074 1072 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03852 11024 1072 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03851 11074 1075 1076 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03850 6276 1076 1074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03849 11074 1076 6276 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03848 11074 1076 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03847 11024 1076 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03846 11074 770 771 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03845 1075 771 627 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03844 11074 771 1075 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03843 11074 771 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03842 11024 771 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03841 11074 4356 3409 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03840 8922 3409 3408 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03839 11074 3409 8922 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03838 11074 3409 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03837 11024 3409 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03836 11074 4356 3742 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03835 9309 3742 3597 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03834 11074 3742 9309 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03833 11074 3742 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03832 11024 3742 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03831 11074 4356 3736 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03830 10031 3736 3584 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03829 11074 3736 10031 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03828 11074 3736 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03827 11024 3736 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03826 11074 4356 4357 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03825 5583 4357 4184 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03824 11074 4357 5583 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03823 11074 4357 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03822 11024 4357 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03821 11074 3410 3412 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03820 4356 3412 3411 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03819 11074 3412 4356 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03818 11074 3412 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03817 11024 3412 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03816 11074 1545 599 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03815 600 4995 746 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03814 745 746 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03813 11074 1826 1667 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03812 1668 7701 1827 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03811 2680 1827 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03810 8593 9433 8592 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03809 8595 9087 8761 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03808 11074 9716 8594 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03807 8760 8761 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03806 11074 9597 3571 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03805 3572 3735 3732 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03804 4031 3732 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03803 8883 9633 8884 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03802 8884 9347 8883 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03801 11074 9306 8884 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03800 8882 8883 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03799 7341 7514 7344 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03798 7345 7721 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03797 7343 10028 7342 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03796 10697 7515 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03795 7515 7340 7343 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03794 11074 5926 4721 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03793 4719 4717 4718 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03792 4720 4718 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03791 3347 8922 3346 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03790 3351 9314 3350 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03789 11074 3703 3348 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03788 3712 3350 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03787 5779 5782 5778 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03786 5780 5777 5781 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03785 11074 5774 5775 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03784 5776 5781 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03783 8391 8392 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03782 8217 8222 8221 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03781 8216 8393 8385 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03780 11074 8388 8216 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03779 11074 10638 8393 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03778 8222 8393 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03777 11074 8390 8392 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03776 8221 8393 8391 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03775 8218 8221 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03774 11074 8220 8219 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03773 8385 8222 8220 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03772 8388 8385 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03771 11074 8385 8388 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03770 1568 7678 1567 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03769 1569 2133 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03768 1565 7514 1570 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03767 1890 1566 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03766 1566 1564 1565 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03765 3703 2473 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03764 3706 8124 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03763 1055 4066 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03762 10302 10662 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03761 9945 10289 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03760 9639 9947 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03759 10374 11075 10373 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03758 10375 10378 10377 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03757 11074 10686 10376 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03756 10704 10377 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03755 4424 7041 4427 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03754 4428 5809 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03753 4426 10018 4425 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03752 5202 4613 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03751 4613 4423 4426 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03750 5418 9560 5417 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03749 5419 6276 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03748 5421 6275 5420 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03747 8318 5559 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03746 5559 5416 5421 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03745 5359 5684 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03744 5702 5518 5360 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03743 1112 1227 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03742 1110 1228 1225 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03741 1109 1229 1222 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03740 11074 1813 1109 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03739 11074 2673 1229 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03738 1228 1229 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03737 11074 1230 1227 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03736 1225 1229 1112 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03735 1108 1225 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03734 11074 1224 1111 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03733 1222 1228 1224 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03732 1813 1222 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03731 11074 1222 1813 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03730 10045 10596 9822 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03729 9822 10595 10045 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03728 11074 10680 9822 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03727 10042 10045 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03726 7719 9395 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03725 5671 7601 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03724 3804 7418 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03723 7411 7425 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03722 487 2473 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03721 11074 3413 487 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03720 773 4070 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03719 11074 4066 773 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03718 2594 3382 2598 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03717 2599 2597 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03716 2596 2592 2595 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03715 5015 2789 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03714 2789 2593 2596 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03713 4411 4555 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03712 4919 4410 4412 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03711 11050 11053 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03710 11045 11052 11049 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03709 11043 11056 11044 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03708 11074 11042 11043 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03707 11074 11051 11056 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03706 11052 11056 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03705 11074 11059 11053 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03704 11049 11056 11050 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03703 11046 11049 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03702 11074 11048 11047 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03701 11044 11052 11048 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03700 11042 11044 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03699 11074 11044 11042 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03698 9585 9582 9583 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03697 9584 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03696 9586 10924 9585 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03695 7053 9605 7054 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03694 7054 8644 7053 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03693 11074 7061 7054 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03692 7447 7053 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03691 2579 3983 2751 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03690 2751 2761 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03689 2752 2751 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03688 2577 3983 2749 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03687 2749 2753 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03686 2750 2749 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03685 1688 7701 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03684 1855 1844 1689 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03683 10546 10772 9777 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03682 9777 10564 10546 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03681 11074 9994 9775 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03680 4421 5159 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03679 4584 6127 4422 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03678 9124 9285 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03677 9121 9286 9284 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03676 9120 9288 9280 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03675 11074 9287 9120 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03674 11074 10914 9288 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03673 9286 9288 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03672 11074 9292 9285 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03671 9284 9288 9124 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03670 9122 9284 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03669 11074 9281 9123 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03668 9280 9286 9281 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03667 9287 9280 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03666 11074 9280 9287 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03665 8325 8327 8324 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03664 11074 8320 8670 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03663 11074 8327 8331 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03662 8326 8328 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03661 8322 8321 8326 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03660 8323 8694 8325 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03659 8670 8320 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03658 7905 8026 7902 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03657 11074 8102 8328 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03656 11074 8026 7907 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03655 7903 10257 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03654 7904 8028 7903 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03653 7906 8642 7905 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03652 8328 8102 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03651 7023 10604 7016 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03650 7016 8091 7023 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03649 11074 8297 7015 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03648 2145 3379 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03647 4012 9597 2146 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03646 1651 8012 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03645 1815 1822 1652 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03644 3041 3967 2884 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03643 2883 9597 3041 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03642 2885 5599 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03641 3695 3041 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03640 11074 3040 2882 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03639 2883 3698 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03638 3259 6811 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03637 3664 4311 3260 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03636 11008 11010 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03635 11002 11009 11007 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03634 11000 11011 11001 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03633 11074 10999 11000 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03632 11074 11051 11011 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03631 11009 11011 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03630 11074 11006 11010 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03629 11007 11011 11008 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03628 11003 11007 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03627 11074 11005 11004 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03626 11001 11009 11005 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03625 10999 11001 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03624 11074 11001 10999 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03623 11074 9297 8272 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03622 8271 9296 8273 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03621 8865 8273 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03620 11074 7667 7260 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03619 7261 7445 7438 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03618 9297 7438 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03617 11074 10027 8927 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03616 8928 10700 8929 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03615 10577 8929 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03614 8381 8712 8380 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03613 11074 8706 8977 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03612 11074 8712 8389 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03611 8386 8970 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03610 8387 8707 8386 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03609 8382 8703 8381 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03608 8977 8706 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03607 8372 8709 8371 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03606 11074 8366 8703 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03605 11074 8709 8376 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03604 8377 10594 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03603 8378 8373 8377 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03602 8367 8697 8372 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_03601 8703 8366 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03600 1748 3379 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03599 2741 5918 1749 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03598 10405 10705 10406 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03597 10407 10414 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03596 10694 10708 10405 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03595 9550 10027 9548 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03594 9549 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03593 9547 10854 9550 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03592 3818 4954 3823 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03591 3824 4959 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03590 3820 3817 3819 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03589 3822 4915 3821 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03588 4131 4323 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03587 4320 5539 4131 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03586 11074 6213 4320 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03585 2621 2624 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03584 2551 2623 2555 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03583 2550 2622 2614 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03582 11074 8090 2550 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03581 11074 5083 2622 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03580 2623 2622 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03579 11074 4881 2624 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03578 2555 2622 2621 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03577 2552 2555 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03576 11074 2554 2553 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03575 2614 2623 2554 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03574 8090 2614 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03573 11074 2614 8090 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03572 9988 10218 9766 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03571 9766 9989 9988 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03570 11074 9987 9766 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03569 10179 9988 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03568 6386 9304 6384 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03567 6385 7415 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03566 6387 7655 6386 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03565 7583 8072 7581 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03564 11074 10197 7584 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03563 7582 7584 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03562 4686 7514 4685 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03561 4687 7721 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03560 4689 8643 4688 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03559 4684 6163 4683 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03558 3454 5727 3453 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03557 3455 5728 3631 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03556 11074 10312 3452 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03555 3630 3631 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03554 11074 5554 5555 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03553 8424 5555 5413 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03552 11074 5555 8424 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03551 11074 5555 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03550 11024 5555 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03549 11074 5199 5201 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03548 8145 5201 5200 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03547 11074 5201 8145 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03546 11074 5201 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03545 11024 5201 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03544 11074 8424 8425 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03543 11051 8425 8423 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03542 11074 8425 11051 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03541 11074 8425 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03540 11024 8425 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03539 11074 8424 8422 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03538 10638 8422 8421 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03537 11074 8422 10638 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03536 11074 8422 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03535 11024 8422 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03534 11074 8424 8147 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03533 8048 8147 7938 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03532 11074 8147 8048 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03531 11074 8147 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03530 11024 8147 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03529 11074 8145 8146 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03528 8047 8146 7937 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03527 11074 8146 8047 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03526 11074 8146 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03525 11024 8146 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03524 11074 8424 8289 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03523 10914 8289 8288 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03522 11074 8289 10914 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03521 11074 8289 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03520 11024 8289 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03519 11074 8424 8287 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03518 8286 8287 8285 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03517 11074 8287 8286 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03516 11074 8287 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03515 11024 8287 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03514 1955 1960 7594 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03513 11074 7484 1952 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03512 1956 1958 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03511 7594 1954 1957 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03510 1959 1958 1960 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03509 1954 7484 1953 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03508 11074 11061 11062 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03507 11064 11071 11065 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03506 11063 11065 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03505 11074 6819 5813 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03504 5812 5813 5814 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03503 11074 5811 5812 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03502 6233 5814 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03501 11074 5814 6233 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03500 11074 4070 1082 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03499 1081 1082 1080 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03498 11074 4066 1081 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03497 1079 1080 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03496 11074 1080 1079 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03495 4061 4057 4059 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03494 4060 5295 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03493 4250 4058 4061 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03492 4827 7514 4826 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03491 4828 7721 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03490 4830 8643 4829 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03489 4995 6879 4831 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03488 3450 4939 3449 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03487 3451 4508 3629 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03486 11074 5131 3448 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03485 3628 3629 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03484 5114 5719 5113 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03483 5115 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03482 5117 9308 5116 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03481 5119 8623 5118 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03480 8093 7652 7650 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03479 11074 9987 7654 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03478 7653 7654 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03477 7807 9051 7806 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03476 7808 10399 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03475 7810 8052 7809 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03474 7805 9716 7803 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03473 9030 9046 9032 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03472 9032 9029 9030 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03471 11074 9028 9031 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03470 11074 6379 6380 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03469 6383 7410 6382 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03468 6381 6382 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03467 6802 7460 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03466 11074 10604 6802 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03465 6802 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03464 11074 10888 6802 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03463 6798 6802 6654 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03462 4820 4994 5012 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03461 11074 7484 4821 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03460 4823 5191 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03459 5012 4992 4824 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03458 4825 5191 4994 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03457 4992 7484 4822 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03456 6631 6786 6789 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03455 11074 9605 6632 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03454 6634 6784 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03453 6789 6783 6635 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03452 6636 6784 6786 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03451 6783 9605 6633 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03450 10263 10621 10262 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03449 10264 10258 10263 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03448 10260 10259 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03447 10255 10263 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03446 11074 10256 10261 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03445 10264 10269 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_03444 11074 7439 7028 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03443 7029 7033 7030 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03442 7027 7030 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03441 11074 7068 4801 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03440 4802 4981 4982 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03439 5214 4982 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03438 11074 7041 2291 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03437 2290 5809 2455 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03436 2454 2455 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03435 11074 4070 625 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03434 626 4066 769 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03433 767 769 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03432 11074 3734 3364 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03431 3363 3735 3365 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03430 3722 3365 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03429 8284 10838 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03428 8652 8635 8282 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03427 8283 8636 8652 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03426 11074 8617 8283 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03425 8280 8885 8652 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03424 11074 8633 8281 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03423 4533 5519 4532 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03422 4532 5525 4533 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03421 11074 4553 4532 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03420 4530 4533 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03419 5537 9605 5389 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03418 5389 7437 5537 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03417 11074 9323 5389 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03416 5535 5537 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03415 3286 3295 3289 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03414 3290 3956 3291 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03413 11074 3285 3287 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03412 3288 3291 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03411 9181 9358 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03410 9178 9360 9357 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03409 9177 9359 9352 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03408 11074 9350 9177 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03407 11074 10638 9359 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03406 9360 9359 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03405 11074 9355 9358 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03404 9357 9359 9181 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03403 9179 9357 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03402 11074 9354 9180 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03401 9352 9360 9354 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03400 9350 9352 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03399 11074 9352 9350 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03398 9210 9402 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03397 9207 9404 9401 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03396 9206 9403 9397 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03395 11074 9395 9206 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03394 11074 11051 9403 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03393 9404 9403 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03392 11074 9411 9402 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03391 9401 9403 9210 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03390 9208 9401 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03389 11074 9398 9209 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03388 9397 9404 9398 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03387 9395 9397 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03386 11074 9397 9395 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03385 6478 6477 6480 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03384 6480 10027 6478 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03383 11074 6499 6479 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03382 7353 9412 7352 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03381 7354 11076 7524 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03380 11074 10700 7355 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03379 7523 7524 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03378 10082 10698 9878 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03377 9878 10083 10082 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03376 11074 10708 9878 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03375 9980 10082 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03374 4125 4955 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03373 4310 4631 4126 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03372 11074 4952 4310 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03371 4925 4310 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03370 3002 5753 2839 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03369 2839 3000 3002 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03368 11074 3236 2839 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03367 2998 3002 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03366 887 889 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03365 831 888 885 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03364 829 890 884 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03363 11074 902 829 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03362 11074 2673 890 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03361 888 890 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03360 11074 892 889 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03359 885 890 887 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03358 830 885 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03357 11074 886 832 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03356 884 888 886 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03355 902 884 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03354 11074 884 902 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03353 11074 10591 10836 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03352 10836 10584 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03351 10444 10585 10836 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03350 1409 2417 1411 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03349 1411 2418 1409 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03348 11074 10888 1410 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03347 2191 5901 2196 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03346 2192 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03345 2194 5898 2193 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03344 2589 2195 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_03343 2195 2190 2194 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03342 6368 7848 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03341 6591 7852 6367 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03340 10422 10555 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03339 10545 10547 10423 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03338 3155 7484 1614 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03337 11074 9987 1791 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03336 1613 1791 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03335 8568 8743 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03334 8566 8745 8740 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03333 8564 8744 8738 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03332 11074 8748 8564 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03331 11074 11051 8744 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03330 8745 8744 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03329 11074 8751 8743 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03328 8740 8744 8568 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03327 8565 8740 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03326 11074 8741 8567 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03325 8738 8745 8741 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03324 8748 8738 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03323 11074 8738 8748 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03322 9098 10701 9099 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03321 9099 10083 9098 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03320 11074 10708 9099 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03319 9426 9098 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03318 3003 3009 2685 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03317 2685 3008 3003 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03316 11074 4325 2684 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03315 3258 5181 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03314 4929 5842 3257 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03313 3870 5522 3868 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03312 3869 5521 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03311 3871 4617 3870 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03310 2857 3020 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03309 2856 3021 3018 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03308 2853 3022 3014 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03307 11074 7037 2853 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03306 11074 5083 3022 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03305 3021 3022 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03304 11074 3019 3020 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03303 3018 3022 2857 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03302 2854 3018 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03301 11074 3015 2855 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03300 3014 3021 3015 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03299 7037 3014 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03298 11074 3014 7037 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03297 845 1504 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03296 1248 1495 846 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03295 4454 4997 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03294 5002 4453 4455 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03293 10436 10571 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03292 10560 10559 10435 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03291 5366 5727 5365 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03290 5367 5728 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03289 5521 10024 5366 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03288 4089 4265 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03287 4087 4260 4262 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03286 4086 4268 4258 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03285 11074 9304 4086 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03284 11074 5083 4268 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03283 4260 4268 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03282 11074 5494 4265 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03281 4262 4268 4089 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03280 4085 4262 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03279 11074 4261 4088 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03278 4258 4260 4261 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03277 9304 4258 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03276 11074 4258 9304 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03275 11074 10018 8519 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03274 8520 8648 8649 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03273 8647 8649 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03272 7381 9421 7379 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03271 7380 8155 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03270 7533 10399 7381 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03269 847 1504 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03268 1284 1494 848 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03267 3549 5600 3547 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03266 3548 8661 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03265 3709 8643 3549 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03264 7162 9080 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03263 7161 8453 7159 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03262 11074 4929 2255 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03261 2253 3688 2254 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03260 2407 5490 2327 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03259 2254 2404 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03258 2326 4929 2404 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_03257 2403 2409 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_03256 2262 2406 2256 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03255 2258 5490 2257 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03254 2260 2407 2259 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03253 2261 2985 2262 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03252 11074 4929 2649 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03251 2643 4142 2644 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03250 2650 5490 2557 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03249 2644 2645 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03248 2556 4929 2645 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_03247 2962 2642 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_03246 2654 2646 2647 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03245 2648 5490 2651 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03244 2653 2650 2652 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03243 2655 2984 2654 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03242 11074 5522 4110 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03241 4111 5521 4282 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03240 4281 4282 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03239 2058 2059 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03238 2055 2060 2057 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03237 2051 2061 2053 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03236 11074 7450 2051 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03235 11074 2446 2061 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03234 2060 2061 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_03233 11074 2062 2059 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_03232 2057 2061 2058 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03231 2052 2057 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03230 11074 2054 2056 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03229 2053 2060 2054 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03228 7450 2053 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03227 11074 2053 7450 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03226 6945 8833 6949 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03225 6950 8831 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03224 6947 8824 6946 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03223 9993 8817 6948 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03222 4253 8824 4082 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03221 4082 8817 4253 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03220 11074 10915 4082 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03219 8313 4253 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03218 7832 9433 7830 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03217 7831 8458 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03216 7828 9716 7832 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03215 9939 10652 9901 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03214 11074 10774 9940 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03213 9902 9940 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03212 4712 6278 4711 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03211 4713 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03210 4715 9020 4714 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03209 6285 5918 4716 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03208 9080 10073 9082 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03207 9082 10701 9080 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03206 11074 10708 9079 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03205 2426 2692 1670 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03204 1670 2691 2426 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03203 11074 4325 1669 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03202 2767 5727 2766 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03201 2765 5728 2768 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03200 11074 10257 2764 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03199 2986 2768 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03198 11074 4929 2233 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03197 2232 5490 2234 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03196 2388 2974 2323 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03195 2234 2386 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03194 2322 4929 2386 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_03193 2385 2390 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_03192 2241 2632 2235 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03191 2237 2974 2236 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03190 2238 2388 2239 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03189 2240 3621 2241 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03188 11074 4929 1978 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03187 1974 1993 1976 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03186 1988 2974 1987 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_03185 1976 1977 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03184 1975 4929 1977 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_03183 2967 1985 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_03182 1986 2640 1979 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03181 1981 2974 1980 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03180 1983 1988 1982 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03179 1984 3625 1986 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_03178 9811 10029 9810 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03177 9815 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03176 9813 10028 9812 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03175 10017 10641 9814 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03174 4015 4014 4016 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03173 4016 4012 4015 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03172 11074 4013 4016 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03171 4701 4015 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03170 9528 9526 9527 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03169 9529 9925 9531 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03168 11074 9540 9530 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03167 10206 9531 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03166 2344 2578 2343 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03165 2345 2470 2471 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03164 11074 8713 2342 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03163 5818 2471 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03162 11074 2480 2306 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03161 2306 4014 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03160 3062 2479 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03159 2306 4012 2479 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03158 2479 3714 2306 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03157 11074 4451 4681 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03156 11074 4450 4681 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03155 4681 4452 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03154 4708 4681 4682 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03153 8022 8318 7899 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03152 7899 8316 8022 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03151 11074 8694 7898 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03150 4097 4270 5098 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03149 11074 4272 4098 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03148 4099 4277 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03147 5098 4271 4100 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03146 4101 4277 4270 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03145 4271 4272 4096 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03144 11074 5608 5291 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03143 9560 5291 5290 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03142 11074 5291 9560 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03141 11074 5291 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03140 11024 5291 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03139 11074 5608 5609 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03138 9020 5609 5477 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03137 11074 5609 9020 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03136 11074 5609 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03135 11024 5609 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03134 11074 5608 5597 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03133 10029 5597 5468 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03132 11074 5597 10029 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03131 11074 5597 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03130 11024 5597 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03129 11074 5035 5036 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03128 5608 5036 4873 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03127 11074 5036 5608 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03126 11074 5036 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03125 11024 5036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03124 11074 762 761 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03123 5898 761 619 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03122 11074 761 5898 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03121 11074 761 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03120 11024 761 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03119 11074 762 763 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03118 5911 763 620 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03117 11074 763 5911 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03116 11074 763 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03115 11024 763 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03114 11074 762 760 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03113 6275 760 618 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03112 11074 760 6275 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03111 11074 760 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03110 11024 760 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03109 11074 494 496 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03108 762 496 495 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03107 11074 496 762 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03106 11074 496 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03105 11024 496 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03104 8106 7719 7705 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03103 7705 7701 8106 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03102 11074 7702 7703 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03101 11074 7835 7818 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03100 7819 8054 7820 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03099 8151 7820 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03098 9241 10701 9240 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03097 9242 10073 9422 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03096 11074 10700 9243 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03095 9421 9422 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03094 10233 10568 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03093 11074 10604 10233 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03092 10233 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03091 11074 10888 10233 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03090 10279 10233 10236 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03089 6218 8654 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03088 11074 10604 6218 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03087 6218 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03086 11074 10888 6218 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_03085 6137 6218 5991 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03084 10553 10551 10430 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03083 10430 10780 10553 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03082 11074 10774 10430 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03081 10550 10553 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03080 11074 1067 765 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03079 5918 765 622 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03078 11074 765 5918 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03077 11074 765 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03076 11024 765 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03075 11074 1067 764 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03074 5599 764 621 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03073 11074 764 5599 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03072 11074 764 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03071 11024 764 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03070 11074 1067 1069 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03069 7678 1069 1068 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03068 11074 1069 7678 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03067 11074 1069 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03066 11024 1069 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03065 11074 499 498 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03064 1067 498 497 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03063 11074 498 1067 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03062 11074 498 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03061 11024 498 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03060 11074 1610 1612 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03059 6277 1612 1611 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03058 11074 1612 6277 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03057 11074 1612 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03056 11024 1612 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03055 11074 1610 1316 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03054 7711 1316 1193 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03053 11074 1316 7711 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03052 11074 1316 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03051 11024 1316 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03050 11074 1610 1312 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03049 5719 1312 1185 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03048 11074 1312 5719 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03047 11074 1312 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03046 11024 1312 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03045 11074 1079 1078 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03044 1610 1078 1077 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03043 11074 1078 1610 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03042 11074 1078 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03041 11024 1078 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03040 8831 8654 8524 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03039 8524 10564 8831 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03038 11074 8912 8523 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03037 9055 10083 9054 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03036 9058 10709 9060 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03035 11074 10700 9056 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03034 9083 9060 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_03033 11074 3063 2907 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03032 2908 3062 3061 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03031 3070 3061 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03030 11074 5918 3380 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03029 3381 3379 3383 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03028 4038 3383 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03027 11074 3739 3590 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03026 3591 3738 3740 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03025 4717 3740 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03024 11074 5581 5250 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03023 5901 5250 5251 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03022 11074 5250 5901 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03021 11074 5250 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03020 11024 5250 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03019 11074 5581 5582 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03018 6278 5582 5448 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03017 11074 5582 6278 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03016 11074 5582 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03015 11024 5582 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03014 11074 5577 5578 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03013 5581 5578 5441 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03012 11074 5578 5581 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03011 11074 5578 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03010 11024 5578 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03009 10044 9610 9611 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03008 9611 9609 10044 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03007 11074 9613 9608 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_03006 11074 3057 2770 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03005 2770 3714 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03004 3065 2769 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03003 2770 3033 2769 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03002 2769 4014 2770 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_03001 11074 11072 7949 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_03000 7950 10710 8158 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02999 8062 8158 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02998 11074 6277 3340 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02997 3341 5600 3342 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02996 3704 3342 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02995 1768 5599 1771 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02994 1769 3735 1895 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02993 11074 5293 1770 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02992 1898 1895 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02991 454 1545 453 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02990 455 472 456 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02989 11074 6261 450 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02988 451 456 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02987 10777 10771 8820 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02986 11074 10915 8818 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02985 8819 8818 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02984 1452 1454 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02983 1450 1453 1451 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02982 1446 1455 1445 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02981 11074 2432 1446 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02980 11074 2446 1455 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02979 1453 1455 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02978 11074 1461 1454 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02977 1451 1455 1452 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02976 1447 1451 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02975 11074 1449 1448 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02974 1445 1453 1449 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02973 2432 1445 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02972 11074 1445 2432 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02971 11074 9033 7770 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02970 7770 8748 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02969 7769 8407 7770 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02968 11074 8388 7740 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02967 7740 7739 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02966 7738 8409 7740 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02965 6244 6851 6013 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02964 6013 6518 6244 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02963 11074 6243 6013 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02962 6152 6244 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02961 9229 10378 9232 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02960 9233 9419 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02959 9231 11075 9230 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02958 9418 9420 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02957 9420 9228 9231 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02956 7691 7689 7693 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02955 7693 7690 7691 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02954 11074 10255 7693 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02953 8096 7691 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02952 7019 7450 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02951 7606 7611 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02950 7689 7466 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02949 3625 3837 3446 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02948 3446 4567 3625 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02947 11074 4553 3444 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02946 3873 3875 3874 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02945 3874 4539 3873 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02944 11074 3872 3874 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02943 6201 3873 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02942 7936 8141 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02941 7934 8142 8139 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02940 7933 8144 8136 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02939 11074 8409 7933 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02938 11074 10638 8144 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02937 8142 8144 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02936 11074 8734 8141 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02935 8139 8144 7936 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02934 7932 8139 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02933 11074 8138 7935 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02932 8136 8142 8138 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02931 8409 8136 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02930 11074 8136 8409 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02929 11074 3337 2469 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02928 2469 2466 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02927 2299 2750 2469 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02926 1128 4981 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02925 1291 1881 1129 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02924 7475 7474 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02923 7452 7037 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02922 10575 10800 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02921 10839 10838 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02920 10772 10771 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02919 10619 4254 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02918 1776 5898 1780 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02917 1777 5600 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02916 1779 6277 1778 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02915 2211 1902 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02914 1902 1789 1779 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02913 2933 9309 2936 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02912 2937 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02911 2935 5918 2934 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02910 3084 3085 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02909 3085 2932 2935 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02908 5138 6214 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02907 5140 6215 5139 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02906 1478 1479 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02905 1475 1480 1477 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02904 1473 1481 1472 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02903 11074 1844 1473 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02902 11074 2446 1481 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02901 1480 1481 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02900 11074 1839 1479 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02899 1477 1481 1478 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02898 1471 1477 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02897 11074 1474 1476 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02896 1472 1480 1474 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02895 1844 1472 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02894 11074 1472 1844 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02893 6037 6269 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02892 6036 6270 6268 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02891 6033 6272 6267 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02890 11074 6493 6033 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02889 11074 8048 6272 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02888 6270 6272 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02887 11074 6273 6269 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02886 6268 6272 6037 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02885 6034 6268 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02884 11074 6271 6035 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02883 6267 6270 6271 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02882 6493 6267 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02881 11074 6267 6493 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02880 4657 5911 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02879 11074 7678 4657 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02878 4657 4653 4656 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02877 4655 4654 4657 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02876 6096 6240 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02875 6827 6486 6097 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02874 6359 8733 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02873 6537 6358 6360 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02872 6489 5811 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02871 5757 5552 5172 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02870 5172 10606 5757 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02869 11074 9304 5171 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02868 2616 9379 2618 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02867 11074 2958 2956 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02866 11074 9379 2619 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02865 2620 2964 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02864 2615 2961 2620 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02863 2617 2957 2616 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02862 2956 2958 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02861 3214 6431 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02860 4936 3213 3215 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02859 9806 10027 9804 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02858 9805 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02857 10011 10641 9806 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02856 8369 8708 8368 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02855 11074 8701 8697 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02854 11074 8708 8379 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02853 8374 8699 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02852 8375 8702 8374 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02851 8370 8983 8369 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02850 8697 8701 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02849 4027 7527 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02848 4029 6574 4028 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02847 2330 6140 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02846 2427 2426 2331 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02845 3480 3651 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02844 3652 4314 3479 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02843 1798 1964 1623 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02842 1622 2637 1798 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02841 1624 2962 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02840 1805 1798 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02839 11074 1796 1621 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02838 1622 3611 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02837 8857 8858 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02836 8853 8859 8855 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02835 8851 8860 8850 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02834 11074 8848 8851 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02833 11074 10914 8860 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02832 8859 8860 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02831 11074 8856 8858 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02830 8855 8860 8857 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02829 8849 8855 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02828 11074 8852 8854 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02827 8850 8859 8852 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02826 8848 8850 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02825 11074 8850 8848 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02824 6240 5816 5817 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02823 5817 6150 6240 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02822 11074 7480 5815 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02821 8414 8733 8412 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02820 11074 8727 8724 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02819 11074 8733 8416 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02818 8417 8728 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02817 8413 8729 8417 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02816 8415 8725 8414 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02815 8724 8727 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02814 6605 10704 6604 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02813 6606 8770 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02812 6906 9747 6605 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02811 6643 7648 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02810 6793 6791 6644 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02809 2560 5809 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02808 3029 7041 2561 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02807 5196 10029 5195 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02806 5197 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02805 5192 10028 5198 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02804 5194 5191 5193 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02803 10982 10986 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02802 10981 10985 10984 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02801 10976 10987 10979 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02800 11074 10990 10976 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02799 11074 11051 10987 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02798 10985 10987 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02797 11074 10989 10986 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02796 10984 10987 10982 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02795 10978 10984 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02794 11074 10980 10983 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02793 10979 10985 10980 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02792 10990 10979 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02791 11074 10979 10990 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02790 11074 10613 10453 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02789 10454 10611 10612 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02788 10610 10612 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02787 7634 7633 7635 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02786 7635 9297 7634 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02785 11074 7631 7632 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02784 7723 7721 7722 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02783 7724 8038 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02782 7726 8126 7725 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02781 8112 9308 7720 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02780 7335 10687 7334 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02779 11074 7512 7509 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02778 11074 10687 7339 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02777 7337 7817 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02776 7338 7513 7337 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02775 7336 7739 7335 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02774 7509 7512 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02773 5844 10687 5843 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02772 11074 5846 5841 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02771 11074 10687 5847 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02770 5848 6877 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02769 5849 5850 5848 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02768 5845 5842 5844 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02767 5841 5846 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02766 6533 10687 6532 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02765 11074 6528 6530 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02764 11074 10687 6536 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02763 6534 7526 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02762 6535 6531 6534 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02761 6529 6527 6533 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02760 6530 6528 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02759 11074 9729 7829 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02758 7826 7829 7827 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02757 11074 8152 7826 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02756 7825 7827 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02755 11074 7827 7825 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02754 4593 4954 4592 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02753 4595 4631 4594 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02752 11074 4955 4591 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02751 5131 4594 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02750 7112 10687 7111 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02749 11074 7107 7108 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02748 11074 10687 7113 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02747 7114 8429 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02746 7115 7116 7114 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02745 7110 7109 7112 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02744 7108 7107 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02743 10599 9552 9553 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02742 9553 9609 10599 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02741 11074 9559 9551 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02740 1762 1890 1891 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02739 1891 1893 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02738 3079 1891 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02737 1571 1574 1572 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02736 1572 1575 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02735 2167 1572 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02734 4348 2140 2141 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02733 2141 2138 4348 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02732 11074 10258 2139 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02731 9725 10705 9730 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02730 9731 10701 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02729 9727 10395 9726 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02728 9729 11072 9728 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02727 6073 6574 6072 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02726 6074 7848 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02725 6179 7852 6073 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02724 1030 9020 1029 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02723 1031 6276 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02722 5809 5911 1030 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02721 2763 3050 2762 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02720 2762 2761 2763 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02719 11074 11042 2760 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02718 8629 9298 8266 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02717 8266 8865 8629 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02716 11074 10197 8265 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02715 8543 8713 8712 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02714 8545 8713 8714 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02713 8546 9016 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02712 8548 8714 8547 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02711 11074 8709 8544 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02710 8202 8862 8201 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02709 8203 8262 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02708 8199 9298 8200 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02707 8817 8254 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02706 8254 8198 8199 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02705 3939 3947 3945 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02704 11074 3938 3940 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02703 3943 3941 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02702 3945 3942 3944 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02701 3946 3941 3947 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02700 3942 3938 3935 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02699 10409 11076 10411 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02698 10413 10709 10412 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02697 11074 10708 10410 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02696 10408 10412 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02695 11074 10031 3972 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02694 3973 9314 3975 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02693 3974 3975 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02692 11074 2168 2169 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02691 2170 4453 2171 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02690 2490 2171 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02689 1533 9597 1532 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02688 1530 1529 1533 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02687 1534 3967 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02686 1528 1533 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02685 11074 1862 1531 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02684 1530 5599 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_02683 7020 7019 7021 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02682 7021 7690 7020 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02681 11074 8903 7021 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02680 7046 7020 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02679 10403 10705 10402 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02678 10400 10414 10404 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02677 11074 10708 10401 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02676 10399 10404 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02675 4230 5297 4229 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02674 4231 4465 4362 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02673 11074 4361 4232 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02672 4369 4362 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02671 5561 6241 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02670 11074 5811 5561 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02669 4535 5519 4537 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02668 4537 5525 4535 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02667 11074 4553 4536 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02666 9325 10366 9166 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02665 9166 9347 9325 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02664 11074 10017 9166 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02663 9323 9325 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02662 585 739 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02661 584 740 736 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02660 582 741 734 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02659 11074 1005 582 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02658 11074 5262 741 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02657 740 741 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02656 11074 1008 739 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02655 736 741 585 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02654 583 736 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02653 11074 735 586 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02652 734 740 735 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02651 1005 734 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02650 11074 734 1005 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02649 8590 9424 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02648 8758 8756 8591 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02647 8589 9724 8758 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02646 11074 9421 8589 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02645 8587 8760 8758 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02644 11074 9073 8588 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02643 9718 10710 9717 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02642 9719 10395 9721 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02641 11074 11072 9720 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02640 9716 9721 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02639 11074 4005 5009 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02638 5009 4003 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02637 4002 4451 5009 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02636 2205 2203 2204 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02635 2206 2213 2210 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02634 11074 3349 2207 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02633 5302 2210 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02632 9191 9372 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02631 9190 9373 9370 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02630 9188 9374 9367 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02629 11074 9376 9188 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02628 11074 10638 9374 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02627 9373 9374 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02626 11074 9375 9372 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02625 9370 9374 9191 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02624 9189 9370 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02623 11074 9368 9192 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02622 9367 9373 9368 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02621 9376 9367 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02620 11074 9367 9376 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02619 6453 6454 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02618 6342 6345 6344 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02617 6340 6456 6452 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02616 11074 6468 6340 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02615 11074 10914 6456 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02614 6345 6456 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02613 11074 10257 6454 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02612 6344 6456 6453 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02611 6339 6344 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02610 11074 6341 6343 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02609 6452 6345 6341 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02608 6468 6452 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02607 11074 6452 6468 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02606 11074 10228 10589 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02605 10589 10139 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02604 10140 10232 10589 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02603 23 142 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02602 20 143 141 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02601 19 144 137 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02600 11074 341 19 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02599 11074 2673 144 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02598 143 144 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02597 11074 145 142 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02596 141 144 23 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02595 21 141 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02594 11074 139 22 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02593 137 143 139 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02592 341 137 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02591 11074 137 341 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02590 7778 7779 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02589 7775 7780 7777 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02588 7771 7781 7773 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02587 11074 8407 7771 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02586 11074 8048 7781 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02585 7780 7781 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02584 11074 7802 7779 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02583 7777 7781 7778 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02582 7772 7777 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02581 11074 7774 7776 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02580 7773 7780 7774 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02579 8407 7773 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02578 11074 7773 8407 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02577 8007 9552 7610 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02576 7610 8644 8007 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02575 11074 8009 7609 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02574 7293 8092 7291 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02573 7292 8709 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02572 8107 8713 7293 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02571 8215 8411 8357 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02570 8357 9033 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02569 8358 8357 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02568 10837 10836 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02567 10847 10832 10834 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02566 8453 10698 8452 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02565 8452 10083 8453 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02564 11074 10708 8451 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02563 4792 4972 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02562 4789 4974 4971 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02561 4788 4973 4966 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02560 11074 5191 4788 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02559 11074 5262 4973 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02558 4974 4973 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02557 11074 4969 4972 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02556 4971 4973 4792 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02555 4790 4971 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02554 11074 4968 4791 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02553 4966 4974 4968 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02552 5191 4966 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02551 11074 4966 5191 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02550 4743 4902 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02549 4741 4904 4900 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02548 4739 4903 4896 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02547 11074 8918 4739 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02546 11074 5083 4903 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02545 4904 4903 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02544 11074 5097 4902 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02543 4900 4903 4743 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02542 4740 4900 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02541 11074 4899 4742 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02540 4896 4904 4899 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02539 8918 4896 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02538 11074 4896 8918 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02537 10544 10542 10421 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02536 10421 10541 10544 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02535 11074 10774 10421 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02534 10540 10544 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02533 8341 8358 7909 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02532 7909 8103 8341 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02531 11074 8206 7908 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02530 11059 11057 11060 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02529 11060 11058 11059 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02528 11074 11054 11055 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02527 3540 5918 3541 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02526 3542 6277 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02525 3976 3706 3540 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02524 88 1545 87 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02523 89 472 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02522 220 4673 88 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02521 3692 4976 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02520 11074 3958 3692 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02519 3692 3959 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02518 11074 4979 3692 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02517 3688 3692 3524 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02516 11074 7068 2886 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02515 2887 3047 3045 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02514 3044 3045 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02513 11074 4410 3482 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02512 3481 3893 3653 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02511 3658 3653 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02510 9574 9572 9573 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02509 9575 9586 9577 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02508 11074 9579 9576 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02507 9571 9577 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02506 8299 8922 8304 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02505 8300 8661 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02504 8302 10028 8301 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02503 8657 8297 8303 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02502 8363 8708 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02501 8690 8709 8363 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02500 11074 10606 8690 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02499 11074 7084 7077 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02498 7078 7476 7079 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02497 7702 7079 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02496 8406 8437 8404 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02495 8405 8403 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02494 8402 10704 8406 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02493 1510 5898 1508 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02492 1509 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02491 2728 7711 1510 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02490 6365 10399 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02489 6592 9716 6366 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02488 79 747 78 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02487 80 482 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02486 452 219 79 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02485 463 1545 461 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02484 462 472 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02483 464 5837 463 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02482 11074 5842 3238 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02481 3237 5181 3239 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02480 3236 3239 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02479 3437 5119 3440 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02478 3438 5123 3619 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02477 11074 5131 3439 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02476 3617 3619 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02475 9022 9020 9021 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02474 9023 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02473 9025 10028 9024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02472 9613 10963 9019 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02471 1158 7478 1156 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02470 1157 5599 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02469 1881 8126 1158 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02468 1515 5809 1514 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02467 1516 4981 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02466 1513 7041 1517 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02465 2462 1512 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02464 1512 1511 1513 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02463 11074 2472 1043 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02462 1043 2474 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02461 1041 1044 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02460 1043 1042 1044 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02459 1044 10256 1043 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02458 10006 10614 9789 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02457 9789 10615 10006 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02456 11074 10024 9788 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02455 11074 7050 7049 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02454 7047 7046 7048 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02453 7045 7048 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02452 11074 6798 6441 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02451 6443 7022 6442 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02450 6440 6442 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02449 3963 3962 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02448 11074 10596 3963 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02447 3963 3961 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02446 11074 10595 3963 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02445 5168 3963 3960 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02444 11074 2602 2797 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02443 11074 2601 2797 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02442 2797 2801 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02441 2799 2797 2798 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02440 8603 9057 8602 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02439 8605 9421 8769 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02438 11074 9433 8604 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02437 8768 8769 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02436 1059 4070 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02435 11074 8124 1059 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02434 1059 3092 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02433 11074 4066 1059 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02432 1061 1059 1060 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02431 11074 2791 2793 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02430 2795 2792 2794 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02429 3403 2794 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02428 3429 3609 3814 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02427 11074 3606 3430 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02426 3432 3607 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02425 3814 3605 3431 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02424 3433 3607 3609 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02423 3605 3606 3428 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02422 4731 6941 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02421 4883 9993 4730 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02420 11074 4880 4883 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02419 4881 4883 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02418 8439 10698 8438 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02417 8441 10073 8440 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02416 11074 11072 8436 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02415 8437 8440 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02414 11074 9716 9258 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02413 9259 9433 9431 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02412 9750 9431 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02411 11074 1881 1741 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02410 1741 3714 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02409 2147 1879 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02408 1741 6220 1879 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02407 1879 4014 1741 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02406 7868 8623 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02405 8078 8834 7869 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02404 11074 8007 8078 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02403 8262 8078 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02402 2363 7711 2366 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02401 2367 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02400 2365 7478 2364 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02399 2602 2504 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02398 2504 2362 2365 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02397 5450 6275 5449 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02396 5451 5583 5584 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02395 11074 7514 5452 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02394 6861 5584 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02393 1432 1433 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02392 1429 1435 1430 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02391 1425 1434 1424 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02390 11074 1423 1425 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02389 11074 2673 1434 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02388 1435 1434 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02387 11074 1431 1433 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02386 1430 1434 1432 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02385 1426 1430 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02384 11074 1427 1428 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02383 1424 1435 1427 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02382 1423 1424 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02381 11074 1424 1423 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02380 7918 8116 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02379 7917 8117 8115 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02378 7915 8119 8114 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02377 11074 8122 7915 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02376 11074 10638 8119 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02375 8117 8119 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02374 11074 8120 8116 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02373 8115 8119 7918 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02372 7916 8115 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02371 11074 8118 7919 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02370 8114 8117 8118 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02369 8122 8114 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02368 11074 8114 8122 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02367 10542 10568 10204 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02366 10204 10564 10542 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02365 11074 10610 10202 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02364 6348 6506 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02363 6487 6496 6347 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02362 11074 7484 5579 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02361 5579 11042 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02360 5252 6493 5579 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02359 5562 7749 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02358 6259 6246 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02357 8654 8090 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02356 10568 10567 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02355 10583 9922 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02354 10890 10213 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02353 5785 7041 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02352 5783 7042 5784 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02351 11074 10619 5783 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02350 5782 5783 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02349 1117 1257 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02348 1114 1259 1256 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02347 1113 1258 1252 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02346 11074 1826 1113 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02345 11074 2446 1258 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02344 1259 1258 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02343 11074 1437 1257 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02342 1256 1258 1117 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02341 1115 1256 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02340 11074 1253 1116 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02339 1252 1259 1253 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02338 1826 1252 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02337 11074 1252 1826 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02336 11074 6859 5836 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02335 10687 5836 5835 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02334 11074 5836 10687 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02333 11074 5836 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02332 11024 5836 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02331 11074 6859 6860 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02330 8733 6860 6682 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02329 11074 6860 8733 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02328 11074 6860 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02327 11024 6860 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02326 11074 6255 6256 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02325 6859 6256 6019 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02324 11074 6256 6859 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02323 11074 6256 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02322 11024 6256 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02321 7668 7667 7669 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02320 7669 9379 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02319 8094 7669 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02318 10230 10608 10229 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02317 10229 10606 10230 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02316 11074 10854 10229 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02315 10228 10230 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02314 6379 10604 3807 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02313 3807 8091 6379 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02312 11074 9304 3806 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02311 1555 3413 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02310 2138 2473 1554 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02309 5541 8623 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02308 6116 8617 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02307 5093 8839 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02306 4975 7085 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02305 6651 8090 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02304 6796 8635 6652 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02303 6653 8636 6796 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02302 11074 7652 6653 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02301 6649 8297 6796 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02300 11074 8633 6650 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02299 5748 2412 1661 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02298 1661 2413 5748 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02297 11074 4325 1659 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02296 4189 4277 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02295 4500 4272 4190 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02294 1634 1805 1635 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02293 1636 2998 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02292 1806 1804 1634 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02291 7155 7158 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02290 7150 7157 7156 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02289 7148 7160 7149 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02288 11074 7147 7148 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02287 11074 8048 7160 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02286 7157 7160 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02285 11074 7154 7158 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02284 7156 7160 7155 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02283 7151 7156 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02282 11074 7153 7152 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02281 7149 7157 7153 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02280 7147 7149 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02279 11074 7149 7147 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02278 8601 9429 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02277 8767 9732 8600 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02276 10488 10687 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02275 11054 11042 10489 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02274 8751 9046 8576 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02273 8576 8750 8751 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02272 11074 8749 8575 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02271 2338 3379 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02270 10258 6275 2339 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02269 2328 8014 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02268 2416 2415 2329 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02267 11074 3007 2843 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02266 2844 5535 3006 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02265 3654 3006 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02264 2834 2996 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02263 3219 4410 2835 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02262 8877 8880 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02261 8875 8879 8876 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02260 8871 8881 8870 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02259 11074 8869 8871 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02258 11074 10914 8881 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02257 8879 8881 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02256 11074 8878 8880 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02255 8876 8881 8877 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02254 8874 8876 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02253 11074 8873 8872 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02252 8870 8879 8873 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02251 8869 8870 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02250 11074 8870 8869 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02249 9622 10027 9621 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02248 9623 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02247 10248 10963 9622 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02246 11074 7615 7616 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02245 7617 7618 7619 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02244 8081 7619 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02243 4014 9987 1756 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02242 11074 2481 1888 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02241 1755 1888 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02240 579 1495 731 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02239 731 1494 580 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02238 581 729 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02237 577 984 731 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02236 11074 1489 576 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02235 11074 1005 578 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02234 2692 731 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02233 7957 8651 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02232 8017 8089 7958 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02231 3881 5153 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02230 4291 5718 3882 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02229 11074 7685 7687 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02228 7686 7684 7688 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02227 10564 7688 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02226 7294 7721 7298 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02225 7299 7711 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02224 7296 9308 7295 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02223 7695 8725 7297 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02222 9235 10697 9234 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02221 9239 9421 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02220 9237 9433 9236 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02219 9680 9716 9238 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02218 9063 10073 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02217 9073 10708 9064 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02216 8101 8318 7901 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02215 7901 8316 8101 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02214 11074 8954 7900 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02213 5751 5755 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02212 8816 5748 5749 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02211 2384 2962 2231 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02210 2231 5124 2384 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02209 11074 3615 2230 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02208 3826 4939 3825 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02207 3831 4508 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02206 3828 4959 3827 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02205 3830 4954 3829 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02204 11074 4929 3910 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02203 3904 4312 3903 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02202 3915 4306 3918 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02201 3903 3906 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02200 3902 4929 3906 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_02199 3917 3914 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_02198 3916 3905 3907 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02197 3909 4306 3908 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02196 3912 3915 3911 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02195 3913 4322 3916 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02194 11074 4929 3502 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02193 3499 3664 3501 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02192 3666 4306 3510 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_02191 3501 3667 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02190 3500 4929 3667 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_02189 3938 3670 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_02188 3509 3668 3503 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02187 3505 4306 3504 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02186 3507 3666 3506 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02185 3508 4320 3509 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_02184 8527 8657 8526 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02183 8528 8659 8660 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02182 11074 8658 8529 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02181 8913 8660 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02180 11074 10018 6474 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02179 6474 6476 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02178 7468 6475 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02177 6474 6473 6475 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02176 6475 8713 6474 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02175 9661 10684 9659 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02174 11074 9663 10701 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02173 11074 10684 9664 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02172 9665 10257 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02171 9660 9666 9665 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02170 9662 9947 9661 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_02169 10701 9663 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02168 7280 7670 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02167 7667 7673 7281 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02166 7279 7459 7667 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02165 11074 7460 7279 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02164 7279 7463 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_02163 2093 7678 2092 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02162 2092 5898 2093 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02161 11074 2736 2091 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02160 11074 11066 7946 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02159 7947 8155 8154 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02158 8460 8154 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02157 11074 5837 5838 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02156 5839 10687 5840 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02155 6524 5840 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02154 7186 10399 7185 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02153 7187 9421 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02152 7189 8453 7188 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02151 7534 9716 7184 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02150 10574 10575 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02149 11074 10604 10574 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02148 10574 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02147 11074 10888 10574 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02146 10832 10574 10441 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02145 3556 7465 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02144 11074 3714 3556 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02143 3556 6251 3554 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02142 3555 3718 3556 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02141 7856 9987 9633 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02140 7860 9987 8065 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02139 7857 8072 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02138 7859 8065 7858 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02137 11074 8064 7855 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02136 4608 6221 4612 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02135 4614 5809 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02134 4610 10018 4609 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02133 4956 6220 4611 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02132 4417 7711 4416 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02131 4418 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02130 4415 8921 4414 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02129 4567 4565 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02128 4565 4413 4415 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02127 6119 6778 5974 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02126 5974 6205 6119 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02125 11074 6206 5973 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02124 11074 8453 8456 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02123 8455 9421 8454 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02122 8756 8454 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02121 11074 6959 6620 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02120 6621 7605 6763 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02119 6762 6763 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02118 11074 449 66 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02117 66 451 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02116 1495 210 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02115 66 213 210 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02114 210 217 66 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02113 5801 6241 5799 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02112 11074 6476 5800 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02111 5798 5800 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02110 11074 10027 7389 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02109 7388 7824 7537 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02108 7536 7537 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02107 11074 4439 4171 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02106 4172 4333 4334 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02105 4342 4334 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02104 11074 2098 1502 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02103 1502 1500 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02102 2459 1503 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02101 1502 2090 1503 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02100 1503 1501 1502 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_02099 8838 8839 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02098 8837 8834 8836 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02097 11074 8835 8837 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02096 8833 8837 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02095 8482 8617 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02094 8615 8834 8482 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02093 11074 8616 8615 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02092 9090 10701 9089 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02091 9091 10709 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02090 9093 9405 9092 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02089 9087 9094 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02088 9094 9088 9093 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02087 6951 6958 7415 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02086 11074 8122 6952 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02085 6955 7484 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02084 7415 6954 6956 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02083 6957 7484 6958 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02082 6954 8122 6953 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02081 5577 10915 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02080 11074 8047 5577 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02079 3585 9309 3589 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02078 3586 9314 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02077 3588 5911 3587 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02076 4048 3737 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_02075 3737 3603 3588 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02074 4123 5159 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02073 4304 6127 4123 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02072 11074 6213 4304 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02071 563 718 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02070 560 719 717 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02069 559 720 712 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02068 11074 711 559 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02067 11074 2446 720 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02066 719 720 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02065 11074 722 718 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02064 717 720 563 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02063 561 717 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02062 11074 714 562 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02061 712 719 714 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02060 711 712 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02059 11074 712 711 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02058 8552 8721 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02057 8551 8722 8720 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02056 8549 8723 8716 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02055 11074 9007 8549 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02054 11074 10638 8723 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02053 8722 8723 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02052 11074 9006 8721 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02051 8720 8723 8552 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02050 8550 8720 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02049 11074 8717 8553 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02048 8716 8722 8717 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02047 9007 8716 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02046 11074 8716 9007 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02045 7867 8075 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02044 7866 8076 8074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02043 7863 8077 8071 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02042 11074 8072 7863 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02041 11074 10914 8077 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02040 8076 8077 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02039 11074 10231 8075 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02038 8074 8077 7867 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02037 7864 8074 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02036 11074 8073 7865 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02035 8071 8076 8073 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02034 8072 8071 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02033 11074 8071 8072 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02032 11074 10605 10865 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02031 10865 10599 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02030 10450 10600 10865 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02029 5606 5603 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02028 11074 5931 5606 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02027 5606 5601 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02026 11074 6175 5606 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02025 18 133 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02024 16 134 130 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02023 15 135 127 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02022 11074 692 15 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02021 11074 2673 135 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02020 134 135 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_02019 11074 329 133 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_02018 130 135 18 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02017 14 130 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02016 11074 129 17 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02015 127 134 129 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02014 692 127 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02013 11074 127 692 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_02012 11074 9932 10142 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02011 10142 9332 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02010 9167 9329 10142 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02009 2000 2413 1648 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02008 1648 2412 2000 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02007 11074 10888 1647 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02006 5032 5040 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02005 11074 5029 5032 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02004 5032 5286 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02003 11074 5610 5032 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_02002 5216 5214 5215 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02001 5215 5565 5216 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_02000 11074 5220 5213 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01999 6693 6874 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01998 6692 6875 6872 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01997 6690 6876 6869 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01996 11074 6867 6690 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01995 11074 8048 6876 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01994 6875 6876 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01993 11074 7144 6874 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01992 6872 6876 6693 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01991 6691 6872 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01990 11074 6870 6694 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01989 6869 6875 6870 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01988 6867 6869 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01987 11074 6869 6867 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01986 2229 2380 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01985 2228 2381 2378 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01984 2225 2382 2375 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01983 11074 7484 2225 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01982 11074 5083 2382 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01981 2381 2382 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01980 11074 3158 2380 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01979 2378 2382 2229 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01978 2226 2378 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01977 11074 2376 2227 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01976 2375 2381 2376 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01975 7484 2375 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01974 11074 2375 7484 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01973 9880 9984 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01972 9985 9987 9879 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01971 10446 10589 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01970 10877 10590 10447 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01969 7846 8059 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01968 8475 9107 7847 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01967 9885 9996 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01966 10137 9997 9886 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01965 4598 4954 4597 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01964 4596 4631 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01963 4926 4955 4598 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01962 1972 3817 1970 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01961 1971 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01960 1973 4915 1972 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01959 2989 2413 2264 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01958 2264 2412 2989 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01957 11074 2688 2263 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01956 7663 7665 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01955 7658 7664 7662 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01954 7656 7666 7657 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01953 11074 7655 7656 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01952 11074 10914 7666 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01951 7664 7666 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01950 11074 8030 7665 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01949 7662 7666 7663 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01948 7659 7662 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01947 11074 7661 7660 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01946 7657 7664 7661 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01945 7655 7657 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01944 11074 7657 7655 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01943 5803 5919 5802 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01942 5804 5801 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01941 5806 9020 5805 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01940 7059 9308 5807 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01939 8442 9080 8444 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01938 8445 9702 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01937 8443 9057 8442 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01936 4152 5911 4150 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01935 4151 9020 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01934 8092 7721 4152 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01933 5284 5283 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01932 5286 5891 5285 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01931 3052 3969 2900 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01930 2899 9308 3052 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01929 2901 5599 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01928 3050 3052 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01927 11074 3967 2898 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01926 2899 3704 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01925 3192 5119 3190 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01924 3191 5123 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01923 3193 4617 3192 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01922 3684 3677 3518 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01921 3518 3675 3684 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01920 11074 3952 3517 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01919 6614 6757 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01918 6613 6756 6755 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01917 6611 6758 6751 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01916 11074 8699 6611 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01915 11074 10914 6758 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01914 6756 6758 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01913 11074 6963 6757 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01912 6755 6758 6614 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01911 6612 6755 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01910 11074 6752 6615 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01909 6751 6756 6752 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01908 8699 6751 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01907 11074 6751 8699 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01906 11074 10225 10221 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01905 10224 10222 10223 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01904 10565 10223 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01903 6683 6864 6684 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01902 6685 6861 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01901 6862 6863 6683 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01900 7816 8054 7814 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01899 7815 8754 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01898 7817 7835 7816 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01897 8582 9095 8580 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01896 8581 9066 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01895 8754 10704 8582 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01894 5000 9002 4844 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01893 4844 4998 5000 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01892 11074 5001 4844 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01891 4997 5000 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01890 5187 5202 5186 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01889 5188 5194 5190 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01888 11074 5771 5189 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01887 5185 5190 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01886 11074 4939 3441 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01885 3442 4508 3620 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01884 3618 3620 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01883 5122 5727 5120 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01882 5121 5728 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01881 5123 10312 5122 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01880 872 9379 870 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01879 11074 866 867 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01878 11074 9379 873 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01877 874 4489 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01876 871 868 874 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01875 869 8885 872 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01874 867 866 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01873 6374 9379 6373 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01872 11074 6369 6370 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01871 11074 9379 6378 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01870 6377 6376 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01869 6375 6371 6377 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01868 6372 8642 6374 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01867 6370 6369 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01866 5325 9379 5324 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01865 11074 5492 5487 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01864 11074 9379 5329 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01863 5327 5490 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01862 5328 5493 5327 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01861 5326 5488 5325 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01860 5487 5492 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01859 4668 4665 4667 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01858 4670 4991 4669 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01857 11074 4666 4671 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01856 7457 4669 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01855 7369 10399 7368 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01854 7370 8155 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01853 7529 8052 7369 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01852 4347 2474 2301 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01851 2301 2472 4347 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01850 11074 4327 2300 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01849 459 1545 457 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01848 458 472 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01847 460 6261 459 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01846 5330 9379 5332 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01845 11074 5498 5494 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01844 11074 9379 5335 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01843 5333 5496 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01842 5334 5499 5333 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01841 5331 9304 5330 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01840 5494 5498 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01839 7892 9560 7891 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01838 7893 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01837 7895 10028 7894 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01836 8938 8305 7896 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01835 10274 10774 10323 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01834 10157 10774 10273 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01833 10275 10652 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01832 10277 10273 10276 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01831 11074 10789 10278 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01830 6609 8064 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01829 7404 10197 6610 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01828 10588 10839 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01827 11074 10604 10588 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01826 10588 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01825 11074 10888 10588 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01824 10590 10588 10445 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01823 6959 10604 6961 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01822 6961 8091 6959 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01821 11074 8699 6960 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01820 11074 6493 5267 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01819 11074 11042 5267 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01818 5267 7484 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01817 5269 5267 5266 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01816 8485 8840 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01815 8620 10197 8486 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01814 11074 6817 5988 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01813 5989 6796 6216 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01812 6130 6216 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01811 9904 10083 9903 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01810 9906 10698 10069 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01809 11074 10700 9905 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01808 10689 10069 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01807 11074 5091 5087 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01806 5088 5667 5089 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01805 5086 5089 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01804 5104 6116 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01803 11074 10604 5104 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01802 5104 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01801 11074 10888 5104 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01800 5103 5104 5102 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01799 9614 10774 10366 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01798 9618 10774 9620 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01797 9619 10268 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01796 9616 9620 9615 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01795 11074 10620 9617 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01794 11074 7042 5178 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01793 5179 7041 5180 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01792 5177 5180 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01791 11074 219 81 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01790 82 482 216 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01789 215 216 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01788 2679 5753 2678 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01787 2678 3000 2679 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01786 11074 3236 2677 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01785 9068 10709 9067 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01784 9069 10073 9070 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01783 11074 10686 9065 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01782 9066 9070 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01781 6617 6766 6616 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01780 6619 6760 6761 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01779 11074 7655 6618 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01778 6759 6761 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01777 2353 9597 2352 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01776 2355 3735 2502 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01775 11074 5293 2354 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01774 2500 2502 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01773 8585 9405 8584 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01772 8586 10698 8755 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01771 11074 10708 8583 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01770 9057 8755 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01769 34 155 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01768 32 157 154 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01767 30 158 150 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01766 11074 348 30 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01765 11074 2673 158 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01764 157 158 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01763 11074 347 155 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01762 154 158 34 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01761 31 154 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01760 11074 153 33 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01759 150 157 153 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01758 348 150 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01757 11074 150 348 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01756 9986 9922 9114 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01755 11074 10774 9274 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01754 9115 9274 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01753 5231 5911 5230 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01752 5233 5600 5234 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01751 11074 6277 5232 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01750 5229 5234 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01749 1165 9314 1169 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01748 1166 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01747 1168 5600 1167 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01746 1573 1303 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01745 1303 1164 1168 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01744 7448 8869 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01743 6109 8848 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01742 6455 9287 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01741 3213 2680 2030 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01740 2030 2681 3213 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01739 11074 2688 2029 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01738 3877 4288 3876 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01737 3876 4290 3877 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01736 11074 4285 3876 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01735 3875 3877 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01734 7333 7506 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01733 7330 7508 7505 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01732 7329 7507 7501 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01731 11074 7739 7329 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01730 11074 8048 7507 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01729 7508 7507 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01728 11074 7509 7506 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01727 7505 7507 7333 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01726 7331 7505 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01725 11074 7503 7332 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01724 7501 7508 7503 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01723 7739 7501 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01722 11074 7501 7739 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01721 7248 10027 7246 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01720 7247 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01719 8080 7425 7248 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01718 6995 7004 6996 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01717 6996 6997 6995 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01716 11074 6994 6996 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01715 6993 6995 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01714 4448 4996 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01713 4452 5580 4449 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01712 6863 7117 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01711 8995 9007 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01710 5851 7147 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01709 5564 6527 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01708 7460 7652 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01707 7444 8082 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01706 2045 2049 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01705 2044 2048 2046 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01704 2040 2050 2039 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01703 11074 2038 2040 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01702 11074 2446 2050 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01701 2048 2050 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01700 11074 2047 2049 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01699 2046 2050 2045 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01698 2041 2046 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01697 11074 2043 2042 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01696 2039 2048 2043 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01695 2038 2039 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01694 11074 2039 2038 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01693 5859 5861 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01692 5854 5860 5858 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01691 5852 5862 5853 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01690 11074 6545 5852 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01689 11074 8048 5862 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01688 5860 5862 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01687 11074 6543 5861 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01686 5858 5862 5859 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01685 5855 5858 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01684 11074 5857 5856 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01683 5853 5860 5857 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01682 6545 5853 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01681 11074 5853 6545 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01680 10871 10875 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01679 10870 10874 10873 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01678 10866 10876 10868 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01677 11074 10880 10866 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01676 11074 10914 10876 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01675 10874 10876 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01674 11074 10879 10875 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01673 10873 10876 10871 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01672 10867 10873 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01671 11074 10869 10872 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01670 10868 10874 10869 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01669 10880 10868 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01668 11074 10868 10880 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01667 7269 10027 7267 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01666 7268 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01665 8648 7450 7269 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01664 2340 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01663 2472 8126 2341 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01662 8893 8642 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01661 2791 1898 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01660 11074 1899 2791 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01659 2791 2208 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01658 11074 2209 2791 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01657 2840 6130 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01656 3425 3003 2838 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01655 9984 9993 9774 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01654 9774 10200 9984 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01653 11074 9991 9773 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01652 1149 4981 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01651 1301 1302 1150 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01650 1297 1292 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01649 11074 1293 1297 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01648 1297 1528 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01647 11074 1291 1297 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01646 1500 1297 1130 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01645 7163 7533 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01644 7165 7828 7164 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01643 7965 8128 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01642 8390 8402 7966 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01641 7735 8121 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01640 8128 8388 7736 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01639 10499 10698 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01638 10699 10708 10500 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01637 10419 10414 10415 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01636 10415 11075 10419 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01635 11074 10686 10416 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01634 3735 8124 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01633 11074 3092 3735 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01632 3735 4066 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01631 11074 4070 3735 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01630 11074 7109 4778 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01629 4779 5181 4953 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01628 4952 4953 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01627 7625 7629 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01626 7624 7628 7627 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01625 7620 7630 7622 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01624 11074 8082 7620 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01623 11074 10914 7630 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01622 7628 7630 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01621 11074 7634 7629 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01620 7627 7630 7625 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01619 7621 7627 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01618 11074 7623 7626 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01617 7622 7628 7623 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01616 8082 7622 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01615 11074 7622 8082 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01614 8308 10027 8306 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01613 8307 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01612 8659 8305 8308 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01611 11074 7740 7327 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01610 7328 7770 7499 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01609 7498 7499 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01608 9825 11019 9823 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01607 11074 10046 9946 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01606 11074 11019 9827 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01605 9828 10257 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01604 9824 9950 9828 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01603 9826 9947 9825 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01602 9946 10046 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01601 9830 11019 9829 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01600 11074 10050 10292 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01599 11074 11019 9832 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01598 9833 10231 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01597 9834 9953 9833 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01596 9831 10289 9830 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01595 10292 10050 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01594 10300 11019 10299 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01593 11074 10294 10668 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01592 11074 11019 10301 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01591 10297 10312 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01590 10298 10296 10297 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01589 10295 10662 10300 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01588 10668 10294 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01587 9848 11019 9852 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01586 11074 10061 10059 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01585 11074 11019 9853 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01584 9850 10024 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01583 9851 9964 9850 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01582 9849 10054 9848 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01581 10059 10061 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01580 10352 11019 10351 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01579 11074 10347 10348 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01578 11074 11019 10355 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01577 10356 10594 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01576 10357 10354 10356 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01575 10353 10350 10352 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01574 10348 10347 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01573 9183 10684 9182 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01572 11074 9364 9419 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01571 11074 10684 9185 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01570 9186 9362 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01569 9187 9365 9186 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01568 9184 9639 9183 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01567 9419 9364 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01566 4745 6277 4744 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01565 4746 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01564 4748 10028 4747 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01563 4915 8839 4749 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01562 11016 11019 11015 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01561 11074 11014 11036 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01560 11074 11019 11022 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01559 11020 11018 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01558 11021 11023 11020 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01557 11017 11028 11016 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01556 11036 11014 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01555 10338 11019 10344 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01554 11074 10679 11006 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01553 11074 11019 10349 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01552 10345 10680 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01551 10346 10678 10345 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01550 10339 10999 10338 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01549 11006 10679 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01548 7521 9046 7351 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01547 7351 8050 7521 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01546 11074 7520 7350 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01545 5921 6278 5920 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01544 5922 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01543 5924 5918 5923 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01542 5933 7514 5925 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01541 9997 10614 9784 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01540 9784 10615 9997 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01539 11074 10231 9782 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01538 1999 2657 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01537 2646 2984 1999 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01536 11074 3632 2646 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01535 4763 5719 4762 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01534 4764 8922 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01533 4766 8921 4765 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01532 4939 8617 4761 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01531 6459 7465 6462 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01530 6461 7615 6460 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01529 11074 8713 6458 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01528 6457 6460 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01527 2869 3033 2868 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01526 2870 10018 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01525 2867 7042 2866 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01524 5727 3034 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01523 3034 2865 2867 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01522 7750 8733 7753 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01521 11074 7756 7752 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01520 11074 8733 7757 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01519 7754 8042 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01518 7755 7758 7754 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01517 7751 7749 7750 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01516 7752 7756 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01515 10336 10684 10335 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01514 11074 10334 10414 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01513 11074 10684 10341 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01512 10342 10680 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01511 10343 10340 10342 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01510 10337 10999 10336 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01509 10414 10334 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01508 2334 2462 2333 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01507 2335 3044 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01506 2337 2727 2336 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01505 5728 2463 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01504 2463 2332 2337 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01503 8864 9296 8503 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01502 8503 9297 8864 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01501 11074 10197 8502 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01500 10075 9979 9751 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01499 9751 9750 10075 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01498 11074 9747 9748 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01497 8432 8430 8435 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01496 8433 8431 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01495 8427 8426 8434 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01494 8429 8443 8428 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01493 6446 6444 6449 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01492 11074 9610 6447 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01491 6450 7006 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01490 6449 6445 6448 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01489 6335 7006 6444 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01488 6445 9610 6334 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01487 9276 9486 9118 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01486 9117 10258 9276 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01485 9119 9503 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01484 9275 9276 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01483 11074 10256 9116 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01482 9117 10269 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01481 6193 6109 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01480 11074 10604 6193 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01479 6193 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01478 11074 10888 6193 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01477 6108 6193 5948 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01476 1824 2680 1666 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01475 1666 2681 1824 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01474 11074 10888 1665 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01473 2316 2493 2315 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01472 2317 2492 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01471 2319 2491 2318 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01470 3377 2490 2320 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01469 1822 2681 1662 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01468 1662 2680 1822 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01467 11074 4325 1660 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01466 1088 1205 4489 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01465 11074 3611 1089 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01464 1091 1210 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01463 4489 1203 1092 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01462 1093 1210 1205 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01461 1203 3611 1090 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01460 10218 10890 10219 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01459 10219 10564 10218 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01458 11074 10215 10220 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01457 10257 9362 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01456 11074 6574 5470 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01455 5469 6896 5598 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01454 5601 5598 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01453 11074 1844 1680 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01452 1681 7701 1838 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01451 1837 1838 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01450 5743 9605 5744 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01449 5744 7437 5743 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01448 11074 9323 5741 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01447 9292 9293 9128 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01446 9128 9290 9292 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01445 11074 9291 9127 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01444 7988 11076 7987 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01443 7989 10698 8153 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01442 11074 10700 7990 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01441 8155 8153 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01440 11074 7514 1047 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01439 1046 5919 1045 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01438 1529 1045 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01437 2912 3065 2911 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01436 2913 3064 3067 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01435 11074 3066 2914 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01434 3076 3067 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01433 8675 8725 7913 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01432 7913 8106 8675 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01431 11074 8107 7912 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01430 6595 6591 6594 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01429 6597 6592 6596 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01428 11074 6908 6593 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01427 6590 6596 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01426 2430 2691 2276 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01425 2276 2692 2430 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01424 11074 2688 2276 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01423 3004 2430 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01422 4305 3008 2690 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01421 2690 3009 4305 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01420 11074 2688 2689 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01419 54 192 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01418 53 193 190 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01417 50 194 187 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01416 11074 724 50 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01415 11074 2446 194 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01414 193 194 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01413 11074 195 192 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01412 190 194 54 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01411 51 190 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01410 11074 188 52 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01409 187 193 188 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01408 724 187 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01407 11074 187 724 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01406 475 753 474 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01405 476 750 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01404 478 1871 477 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01403 472 473 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01402 473 471 478 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01401 956 1495 958 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01400 958 1494 957 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01399 955 959 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01398 952 951 958 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01397 11074 1489 946 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01396 11074 1245 953 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01395 2681 958 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01394 1498 1493 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01393 1857 1494 1499 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01392 1497 1495 1857 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01391 11074 1496 1497 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01390 1492 1490 1857 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01389 11074 1489 1491 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01388 2638 2968 2639 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01387 2639 3611 2638 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01386 11074 2637 2639 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01385 2636 2638 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01384 112 251 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01383 111 252 250 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01382 109 253 246 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01381 11074 244 109 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01380 11074 5262 253 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01379 252 253 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01378 11074 2373 251 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01377 250 253 112 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01376 110 250 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01375 11074 247 113 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01374 246 252 247 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01373 244 246 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01372 11074 246 244 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01371 9496 9497 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01370 9494 9499 9498 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01369 9492 9500 9491 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01368 11074 9489 9492 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01367 11074 10914 9500 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01366 9499 9500 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01365 11074 10312 9497 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01364 9498 9500 9496 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01363 9490 9498 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01362 11074 9493 9495 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01361 9491 9499 9493 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01360 9489 9491 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01359 11074 9491 9489 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01358 11074 10899 10918 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01357 10918 10900 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01356 10898 10897 10918 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01355 10034 9605 9607 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01354 9607 9609 10034 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01353 11074 10017 9606 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01352 1764 5901 1763 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01351 1765 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01350 1767 5719 1766 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01349 1893 1894 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01348 1894 1788 1767 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01347 4984 5564 4804 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01346 4804 4983 4984 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01345 11074 4986 4803 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01344 1024 1027 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01343 852 1026 1022 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01342 849 1028 1020 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01341 11074 1496 849 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01340 11074 5262 1028 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01339 1026 1028 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01338 11074 1025 1027 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01337 1022 1028 1024 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01336 850 1022 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01335 11074 1023 851 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01334 1020 1026 1023 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01333 1496 1020 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01332 11074 1020 1496 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01331 9040 9043 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01330 9036 9042 9041 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01329 9034 9045 9035 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01328 11074 9033 9034 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01327 11074 11051 9045 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01326 9042 9045 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01325 11074 9047 9043 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01324 9041 9045 9040 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01323 9037 9041 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01322 11074 9039 9038 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01321 9035 9042 9039 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01320 9033 9035 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01319 11074 9035 9033 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01318 5830 5831 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01317 5827 5833 5832 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01316 5825 5834 5824 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01315 11074 6819 5825 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01314 11074 8048 5834 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01313 5833 5834 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01312 11074 5829 5831 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01311 5832 5834 5830 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01310 5823 5832 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01309 11074 5826 5828 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01308 5824 5833 5826 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01307 6819 5824 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01306 11074 5824 6819 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01305 298 5488 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01304 299 5488 300 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01303 11074 2957 294 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01302 297 293 295 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01301 296 300 297 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01300 1958 297 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01299 11074 297 1958 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01298 293 2957 292 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01297 8597 9433 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01296 8762 9746 8598 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01295 8596 9750 8762 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01294 11074 9081 8596 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01293 8596 9087 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01292 10862 10865 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01291 10917 10861 10863 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01290 10265 10608 10266 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01289 10266 10606 10265 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01288 11074 10924 10266 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01287 10899 10265 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01286 3154 3804 3153 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01285 3153 7690 3154 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01284 11074 7403 3153 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01283 3152 3154 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01282 6281 6286 6056 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01281 6056 7176 6281 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01280 11074 6280 6056 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01279 6171 6281 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01278 4787 5202 4785 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01277 4786 5194 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01276 4960 5771 4787 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01275 4599 4952 4600 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01274 4601 4631 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01273 5124 4955 4599 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01272 2803 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01271 2964 2965 2804 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01270 2802 3615 2964 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01269 11074 2962 2802 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01268 2802 5124 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_01267 1087 1200 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01266 1086 1201 1198 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01265 1083 1202 1195 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01264 11074 2957 1083 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01263 11074 5083 1202 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01262 1201 1202 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01261 11074 2956 1200 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01260 1198 1202 1087 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01259 1084 1198 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01258 11074 1196 1085 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01257 1195 1201 1196 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01256 2957 1195 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01255 11074 1195 2957 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01254 9742 10701 9740 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01253 9741 10078 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01252 9743 11072 9742 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01251 10143 10142 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01250 10951 10618 10141 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01249 5484 6177 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01248 5610 6180 5485 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01247 2784 3081 2785 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01246 2783 3349 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01245 3072 2782 2784 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01244 6669 6829 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01243 6667 6831 6826 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01242 6665 6830 6822 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01241 11074 8691 6665 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01240 11074 10638 6830 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01239 6831 6830 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01238 11074 6827 6829 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01237 6826 6830 6669 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01236 6666 6826 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01235 11074 6824 6668 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01234 6822 6831 6824 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01233 8691 6822 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01232 11074 6822 8691 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01231 6630 6774 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01230 6627 6775 6773 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01229 6626 6776 6769 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01228 11074 9313 6626 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01227 11074 10914 6776 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01226 6775 6776 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_01225 11074 6777 6774 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01224 6773 6776 6630 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01223 6628 6773 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01222 11074 6770 6629 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01221 6769 6775 6770 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01220 9313 6769 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01219 11074 6769 9313 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01218 8616 9305 7587 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01217 7587 8644 8616 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01216 11074 7585 7586 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01215 11074 7058 7062 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01214 7060 7059 7064 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01213 7061 7064 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01212 10959 2464 2294 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01211 2294 2459 10959 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01210 11074 9987 2293 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01209 8822 10555 8823 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01208 8823 10547 8822 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01207 11074 10915 8823 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01206 8821 8822 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01205 11074 8691 4793 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01204 4794 4984 4977 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01203 4976 4977 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01202 1991 2004 1644 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01201 1644 2006 1991 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01200 11074 2688 1643 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01199 11074 9541 7011 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01198 7013 7063 7014 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01197 7012 7014 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01196 6415 9379 6423 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01195 11074 6781 6777 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01194 11074 9379 6426 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01193 6424 6778 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01192 6417 6782 6424 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01191 6416 9313 6415 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01190 6777 6781 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01189 6965 9379 6964 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01188 11074 6962 6963 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01187 11074 9379 6968 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01186 6969 6967 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01185 6970 6973 6969 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01184 6966 8699 6965 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01183 6963 6962 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01182 8259 8862 8258 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01181 8260 8262 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01180 8256 9298 8255 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01179 8613 8865 8257 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01178 7942 9433 7941 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01177 7943 9421 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01176 8054 8152 7942 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01175 1037 7514 1036 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01174 1034 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01173 1035 1862 1037 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01172 2288 3032 2449 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01171 2449 3029 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01170 2450 2449 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01169 5975 9379 5977 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01168 11074 6212 6427 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01167 11074 9379 5980 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01166 5978 6205 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01165 5979 6126 5978 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01164 5976 8930 5975 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_01163 6427 6212 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01162 10253 10247 10252 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01161 10250 10248 10254 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01160 11074 10249 10251 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01159 10611 10254 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01158 5649 8824 5651 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01157 5652 8833 5653 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01156 11074 8817 5650 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01155 6942 5653 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01154 8496 9298 8495 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01153 8497 8862 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01152 8499 9296 8498 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01151 9290 8631 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01150 8631 8494 8499 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01149 8685 9033 8208 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01148 11074 8930 8209 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01147 8207 8209 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01146 9868 9975 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01145 10070 10692 9869 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01144 11074 10687 10070 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01143 9972 10070 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01142 11074 10080 9101 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01141 9102 9104 9105 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01140 9103 9105 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01139 7834 8059 7833 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01138 7836 8458 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01137 7835 9433 7834 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01136 1559 2481 1560 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01135 1560 10915 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01134 3714 1560 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01133 4009 11042 4011 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01132 4011 7484 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01131 4010 4011 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01130 11074 8124 3091 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01129 2950 3091 3090 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01128 11074 3092 2950 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01127 3410 3090 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01126 11074 3090 3410 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01125 8901 9316 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01124 8906 10197 8902 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01123 2729 10256 2730 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01122 2730 10269 2729 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01121 11074 2728 2730 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01120 3035 2729 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01119 1967 2965 1968 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01118 1966 3615 1967 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01117 1969 5131 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01116 1964 1967 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01115 11074 2962 1965 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01114 1966 5124 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01113 5107 5719 5111 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01112 5112 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01111 5109 9308 5108 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01110 5105 5110 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01109 5110 5106 5109 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01108 8915 10614 8917 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01107 8917 10615 8915 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01106 11074 10995 8916 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01105 11074 8151 7939 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01104 7940 8758 8150 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01103 8053 8150 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01102 10893 10890 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01101 11074 10891 10893 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01100 10893 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01099 11074 10888 10893 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01098 10919 10893 10889 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01097 6058 9107 6057 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01096 6062 8770 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01095 6060 6574 6059 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01094 6173 7852 6061 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01093 9487 9505 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01092 9486 10774 9488 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01091 2569 8709 2573 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01090 2574 2572 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01089 2571 4012 2570 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01088 3036 2739 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01087 2739 2568 2571 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01086 10139 9305 9144 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01085 9144 9609 10139 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01084 11074 9306 9142 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01083 11074 8097 7890 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01082 7889 8096 8098 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01081 8021 8098 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01080 10458 10620 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01079 10621 10774 10459 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01078 8157 10710 7948 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01077 7948 10083 8157 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01076 11074 11072 7948 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01075 8060 8157 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01074 11074 6590 6587 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01073 6589 6898 6588 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01072 6586 6588 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01071 11074 5934 5319 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01070 5322 5321 5323 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01069 5320 5323 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01068 11074 3057 2874 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01067 2875 10018 3038 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01066 3306 3038 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01065 5987 6214 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01064 6128 6215 5987 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01063 11074 6213 6128 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01062 9245 10701 9248 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01061 9249 10078 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01060 9247 10083 9246 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01059 9429 9423 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01058 9423 9244 9247 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01057 11074 1813 1649 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01056 1650 7701 1814 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01055 2413 1814 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01054 3184 3630 3185 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01053 3185 5105 3184 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01052 11074 4553 3185 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01051 3183 3184 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01050 10180 10179 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01049 10178 10184 10181 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01048 11074 10176 10178 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01047 10177 10178 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01046 4693 6276 4692 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01045 4696 8661 4695 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01044 11074 5898 4691 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01043 5275 4695 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01042 4469 4465 4468 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01041 4474 5032 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01040 4471 5297 4470 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01039 4723 4722 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01038 4722 4466 4471 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01037 4211 5771 4210 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01036 4213 5202 4326 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01035 11074 8092 4212 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01034 4325 4326 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01033 11074 9987 1963 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01032 1962 1963 1961 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01031 11074 8617 1962 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01030 8310 1961 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01029 11074 1961 8310 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01028 11074 9382 9016 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01027 9016 9667 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01026 9013 9033 9016 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01025 4808 5918 4807 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01024 4809 9020 4990 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01023 11074 7478 4810 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01022 5226 4990 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01021 4225 4359 4227 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01020 4228 4720 4358 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01019 11074 4710 4226 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01018 4364 4358 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01017 2946 5898 2945 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01016 2947 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01015 2949 7711 2948 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01014 3088 3089 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01013 3089 2944 2949 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01012 7192 7204 7197 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01011 7193 7536 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01010 7195 7837 7194 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01009 7190 7196 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01008 7196 7191 7195 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01007 6732 8472 6736 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01006 6733 6904 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01005 6735 7190 6734 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01004 6898 6899 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_01003 6899 6731 6735 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01002 923 926 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_01001 835 928 917 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_01000 833 929 915 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00999 11074 916 833 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00998 11074 2673 929 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00997 928 929 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00996 11074 925 926 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00995 917 929 923 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00994 834 917 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00993 11074 920 836 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00992 915 928 920 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00991 916 915 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00990 11074 915 916 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00989 5440 5573 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00988 5439 5574 5571 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00987 5436 5575 5568 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00986 11074 5842 5436 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00985 11074 8048 5575 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00984 5574 5575 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00983 11074 5841 5573 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00982 5571 5575 5440 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00981 5437 5571 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00980 11074 5569 5438 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00979 5568 5574 5569 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00978 5842 5568 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00977 11074 5568 5842 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00976 9305 8885 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00975 6760 7484 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00974 9552 9304 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00973 9333 8918 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00972 9566 8699 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00971 9605 9313 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00970 4361 3082 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00969 11074 3084 4361 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00968 5152 6435 5151 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00967 5151 5528 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00966 5150 5151 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00965 4296 4298 4121 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00964 4121 4948 4296 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00963 11074 4295 4121 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00962 4539 4296 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00961 977 978 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00960 839 980 970 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00959 838 981 969 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00958 11074 1456 838 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00957 11074 2446 981 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00956 980 981 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00955 11074 1260 978 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00954 970 981 977 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00953 837 970 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00952 11074 974 840 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00951 969 980 974 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00950 1456 969 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00949 11074 969 1456 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00948 7614 9582 7612 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00947 7613 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00946 7618 7611 7614 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00945 6473 6241 6005 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00944 6005 6233 6473 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00943 11074 7474 6004 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00942 7959 8092 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00941 8026 8713 7960 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00940 10235 10596 10234 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00939 10234 10595 10235 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00938 11074 10231 10234 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00937 10232 10235 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00936 2906 3065 2904 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00935 2905 3064 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00934 3071 3066 2906 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00933 3077 1583 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00932 11074 1573 3077 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00931 3077 1574 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00930 11074 1575 3077 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00929 3995 3993 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00928 4451 3994 3996 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00927 6765 6992 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00926 6766 8122 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00925 9610 8930 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00924 6803 8297 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00923 3402 2590 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00922 11074 3355 3402 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00921 3402 2589 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00920 11074 3079 3402 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00919 2806 3607 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00918 3610 2973 2807 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00917 10937 10941 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00916 10936 10940 10939 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00915 10932 10942 10935 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00914 11074 10945 10932 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00913 11074 11051 10942 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00912 10940 10942 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00911 11074 10944 10941 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00910 10939 10942 10937 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00909 10933 10939 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00908 11074 10934 10938 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00907 10935 10940 10934 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00906 10945 10935 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00905 11074 10935 10945 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00904 1704 1861 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00903 2094 1862 1705 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00902 1703 3040 2094 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00901 11074 7678 1703 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00900 1703 5898 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00899 7963 8394 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00898 8120 8123 7964 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00897 5412 10029 5410 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00896 5411 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00895 6228 8643 5412 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00894 5237 8661 5235 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00893 5236 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00892 6243 8643 5237 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00891 1734 5600 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00890 2140 6277 1735 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00889 3702 3703 3538 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00888 3537 4653 3702 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00887 3539 3704 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00886 10595 3702 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00885 11074 5599 3536 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00884 3537 5898 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00883 11074 3213 2664 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00882 2665 6431 2670 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00881 3198 2670 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00880 7641 7645 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00879 7640 7644 7643 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00878 7636 7646 7638 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00877 11074 7652 7636 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00876 11074 10914 7646 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00875 7644 7646 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00874 11074 8019 7645 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00873 7643 7646 7641 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00872 7637 7643 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00871 11074 7639 7642 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00870 7638 7644 7639 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00869 7652 7638 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00868 11074 7638 7652 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00867 11074 10018 8296 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00866 8295 8938 8298 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00865 8658 8298 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00864 11074 10018 7598 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00863 7597 7600 7599 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00862 8070 7599 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00861 10993 11019 10991 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00860 11074 10988 10989 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00859 11074 11019 10996 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00858 10997 10995 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00857 10992 10998 10997 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00856 10994 10990 10993 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00855 10989 10988 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00854 7961 8121 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00853 8123 8122 7962 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00852 617 9020 615 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00851 616 2133 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00850 3033 5911 617 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00849 1740 9314 1738 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00848 1739 2133 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00847 3057 5911 1740 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00846 8089 2418 2266 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00845 2266 2417 8089 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00844 11074 4325 2265 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00843 11074 5119 3176 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00842 3177 5123 3178 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00841 3175 3178 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00840 7087 10687 7090 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00839 11074 7086 7089 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00838 11074 10687 7093 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00837 7091 7784 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00836 7092 7094 7091 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00835 7088 7085 7087 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00834 7089 7086 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00833 6021 7514 6020 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00832 6022 7721 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00831 6024 10028 6023 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00830 6255 10197 6025 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00829 9315 10020 9157 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00828 11074 10774 9317 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00827 9158 9317 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00826 11074 2481 1307 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00825 1182 1307 1306 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00824 11074 9987 1182 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00823 1308 1306 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00822 11074 1306 1308 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00821 10308 10684 10307 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00820 11074 10673 10705 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00819 11074 10684 10317 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00818 10313 10908 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00817 10314 10674 10313 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00816 10309 10675 10308 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00815 10705 10673 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00814 10328 10684 10327 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00813 11074 10676 11075 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00812 11074 10684 10333 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00811 10330 10995 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00810 10331 10677 10330 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00809 10329 10990 10328 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00808 11075 10676 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00807 10322 10684 10321 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00806 11074 10318 10378 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00805 11074 10684 10325 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00804 10326 10323 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00803 10319 10324 10326 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00802 10320 10332 10322 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00801 10378 10318 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00800 2580 2753 2759 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00799 2759 3723 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00798 2761 2759 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00797 1714 1867 1713 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00796 1715 5240 1869 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00795 11074 1868 1716 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00794 1866 1869 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00793 3626 3630 3447 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00792 3447 5105 3626 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00791 11074 4553 3445 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00790 4191 5131 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00789 4277 4281 4192 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00788 4193 4279 4277 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00787 11074 5124 4193 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00786 4193 4275 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00785 11074 4929 3486 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00784 3483 3654 3485 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00783 3656 3664 3494 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_00782 3485 3657 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00781 3484 4929 3657 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_00780 4940 3662 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_00779 3493 3658 3487 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00778 3489 3664 3488 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00777 3491 3656 3490 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00776 3492 4587 3493 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00775 8621 9489 8487 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00774 11074 10197 8622 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00773 8488 8622 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00772 10364 10684 10369 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00771 11074 10358 10395 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00770 11074 10684 10372 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00769 10370 10366 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00768 10371 10367 10370 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00767 10365 11013 10364 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00766 10395 10358 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00765 10362 10684 10359 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00764 11074 10682 11076 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00763 11074 10684 10368 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00762 10360 11018 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00761 10361 10683 10360 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00760 10363 11028 10362 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00759 11076 10682 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00758 5378 6277 5377 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00757 5379 10031 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00756 5381 8643 5380 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00755 5525 5526 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00754 5526 5376 5381 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00753 3197 3871 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00752 3637 4535 3197 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00751 11074 3632 3637 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00750 11074 4929 3250 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00749 3244 3242 3245 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00748 3251 3664 3148 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_00747 3245 3243 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00746 3147 4929 3243 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_00745 3890 3255 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_00744 3256 3246 3247 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00743 3249 3664 3248 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00742 3253 3251 3252 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00741 3254 4304 3256 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00740 4885 6749 4733 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00739 4733 6942 4885 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00738 11074 5162 4732 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00737 9908 10074 9907 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00736 9909 11063 10072 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00735 11074 10075 9910 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00734 9975 10072 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00733 11074 3032 2453 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00732 2289 2453 2451 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00731 11074 2454 2289 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00730 2452 2451 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00729 11074 2451 2452 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00728 10581 10583 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00727 11074 10604 10581 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00726 10581 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00725 11074 10888 10581 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00724 10582 10581 10443 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00723 8506 10213 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00722 8638 8635 8507 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00721 8508 8636 8638 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00720 11074 8848 8508 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00719 8504 8699 8638 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00718 11074 8633 8505 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00717 10198 10571 10199 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00716 10199 10559 10198 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00715 11074 10197 10199 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00714 10558 10198 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00713 3232 5842 3231 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00712 3235 3230 3232 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00711 3233 5181 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00710 3647 3232 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00709 11074 3242 3234 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00708 3235 3884 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00707 3811 3816 5496 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00706 11074 4501 3808 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00705 3812 3814 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00704 5496 3810 3813 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00703 3815 3814 3816 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00702 3810 4501 3809 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00701 8866 8869 8500 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00700 11074 10774 8632 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00699 8501 8632 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00698 11074 5103 3834 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00697 3835 3833 3836 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00696 3832 3836 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00695 11074 9560 1697 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00694 1698 8922 1858 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00693 3040 1858 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00692 6503 6493 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00691 7084 7739 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00690 9379 10774 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00689 6499 8047 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00688 8983 9382 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00687 11074 5607 5272 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00686 5270 5269 5274 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00685 5271 5274 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00684 1096 2962 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00683 1801 1964 1094 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00682 1095 2637 1801 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00681 11074 1796 1095 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00680 1095 3611 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00679 8314 8313 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00678 8311 8309 8315 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00677 11074 8310 8311 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00676 8312 8311 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00675 8645 9333 8518 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00674 8518 8644 8645 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00673 11074 8647 8517 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00672 11074 6220 2903 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_00671 2903 3714 11074 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_00670 3066 3058 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00669 2903 7042 3058 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_00668 3058 4014 2903 11074 sg13_lv_nmos L=0.13U W=1.29U AS=0.3096P AD=0.3096P PS=3.07U PD=3.07U 
Mtr_00667 11074 4710 4186 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00666 4185 4359 4360 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00665 4467 4360 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00664 6477 6476 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00663 6490 6241 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00662 8408 8407 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00661 8708 9033 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00660 8731 8409 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00659 67 215 70 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00658 71 220 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00657 69 745 68 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00656 1494 212 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00655 212 114 69 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00654 8278 10800 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00653 8277 8635 8279 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00652 8276 8636 8277 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00651 11074 8839 8276 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00650 8274 8642 8277 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00649 11074 8633 8275 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00648 10555 10619 10432 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00647 10432 10564 10555 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00646 11074 10554 10431 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00645 11074 10915 3805 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00644 3802 3805 3803 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00643 11074 8090 3802 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00642 4880 3803 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00641 11074 3803 4880 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00640 2457 10256 2292 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00639 2292 10269 2457 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00638 11074 2578 2292 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00637 2456 2457 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00636 3699 3698 3535 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00635 3534 5599 3699 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00634 3533 9308 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00633 10596 3699 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00632 11074 3974 3532 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00631 3534 3967 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00630 2180 9314 2179 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00629 2181 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00628 2176 8922 2182 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00627 2177 2178 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00626 2178 2175 2176 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00625 5253 7484 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00624 11074 11042 5253 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00623 5881 8922 5880 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00622 5882 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00621 5877 8126 5883 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00620 5878 5879 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00619 5879 5876 5877 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00618 1637 1806 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00617 5142 1807 1638 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00616 97 228 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00615 96 229 227 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00614 94 230 223 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00613 11074 6241 94 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00612 11074 5262 230 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00611 229 230 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00610 11074 231 228 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00609 227 230 97 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00608 95 227 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00607 11074 224 98 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00606 223 229 224 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00605 6241 223 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00604 11074 223 6241 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00603 9803 10023 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00602 9800 10025 10022 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00601 9799 10026 10019 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00600 11074 10020 9799 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00599 11074 10914 10026 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00598 10025 10026 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00597 11074 10024 10023 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00596 10022 10026 9803 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00595 9801 10022 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00594 11074 10021 9802 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00593 10019 10025 10021 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00592 10020 10019 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00591 11074 10019 10020 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00590 8249 8839 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00589 8610 8834 8249 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00588 11074 8835 8610 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00587 11074 10033 10147 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00586 10147 10034 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00585 9816 10032 10147 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00584 11074 4344 4345 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00583 4180 4345 4343 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00582 11074 4342 4180 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00581 4465 4343 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00580 11074 4343 4465 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00579 10138 10137 10205 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00578 10205 10214 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00577 10551 10205 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00576 552 703 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00575 549 704 701 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00574 548 705 699 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00573 11074 1245 548 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00572 11074 2673 705 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00571 704 705 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00570 11074 1244 703 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00569 701 705 552 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00568 550 701 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00567 11074 700 551 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00566 699 704 700 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00565 1245 699 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00564 11074 699 1245 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00563 10129 10542 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00562 10171 10541 10130 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00561 8019 8094 7888 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00560 7888 8095 8019 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00559 11074 8093 7887 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00558 10428 10550 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00557 10548 10559 10429 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00556 11074 10773 10548 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00555 10796 10548 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00554 9175 9343 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00553 9173 9345 9339 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00552 9172 9344 9336 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00551 11074 9335 9172 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00550 11074 10914 9344 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00549 9345 9344 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00548 11074 9341 9343 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00547 9339 9344 9175 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00546 9171 9339 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00545 11074 9338 9174 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00544 9336 9345 9338 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00543 9335 9336 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00542 11074 9336 9335 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00541 10809 10810 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00540 10805 10811 10807 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00539 10801 10812 10803 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00538 11074 10800 10801 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00537 11074 10914 10812 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00536 10811 10812 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00535 11074 10808 10810 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00534 10807 10812 10809 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00533 10802 10807 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00532 11074 10804 10806 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00531 10803 10811 10804 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00530 10800 10803 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00529 11074 10803 10800 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00528 10920 10918 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00527 10977 10919 10921 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00526 11074 10043 10158 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00525 10158 10044 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00524 9820 10042 10158 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00523 9062 9080 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00522 9061 9057 9059 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00521 2311 6278 2310 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00520 2312 3735 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00519 2487 5911 2311 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00518 7065 7069 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00517 7067 7068 7066 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00516 11074 9362 7067 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00515 7063 7067 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00514 2659 4915 2658 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00513 2656 3817 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00512 2657 4617 2659 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00511 3180 3193 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00510 3182 3626 3181 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00509 11074 3632 3182 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00508 3179 3182 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00507 8946 8951 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00506 8945 8950 8948 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00505 8941 8952 8943 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00504 11074 8954 8941 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00503 11074 10914 8952 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00502 8950 8952 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00501 11074 8949 8951 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00500 8948 8952 8946 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00499 8944 8948 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00498 11074 8942 8947 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00497 8943 8950 8942 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00496 8954 8943 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00495 11074 8943 8954 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00494 11074 6496 6011 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00493 6012 6506 6242 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00492 6150 6242 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00491 11074 8290 8294 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00490 8293 8291 8292 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00489 8682 8292 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00488 9873 10701 9872 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00487 9874 10073 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00486 9976 10700 9873 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00485 9691 10083 9689 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00484 9690 10698 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00483 9692 10700 9691 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00482 8908 8906 8907 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00481 8905 10258 8908 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00480 8909 9315 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00479 8903 8908 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00478 11074 10256 8904 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00477 8905 10269 11074 11074 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00476 3577 6278 3575 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00475 3576 3735 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00474 4700 3734 3577 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00473 3565 6278 3564 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00472 3566 3735 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00471 4013 5918 3565 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00470 11074 10006 9790 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00469 9791 10005 10007 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00468 10554 10007 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00467 2822 4939 2823 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00466 2824 4508 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00465 2982 4617 2822 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00464 5134 6215 5133 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00463 5135 6214 5137 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00462 11074 5131 5136 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00461 5132 5137 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00460 3930 4318 3929 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00459 11074 3934 3928 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00458 11074 4318 3936 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00457 3932 4617 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00456 3933 3937 3932 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00455 3931 4553 3930 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00454 3928 3934 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00453 6428 6429 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00452 6328 6333 6332 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00451 6327 6430 6425 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00450 11074 8930 6327 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00449 11074 10914 6430 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00448 6333 6430 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00447 11074 6427 6429 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00446 6332 6430 6428 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00445 6329 6332 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00444 11074 6331 6330 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00443 6425 6333 6331 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00442 8930 6425 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00441 11074 6425 8930 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00440 10201 10568 10203 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00439 10203 10564 10201 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00438 11074 10610 10203 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00437 10200 10201 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00436 6001 6232 6000 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00435 6002 6457 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00434 5998 6251 5997 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00433 7684 6230 5999 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00432 9749 9976 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00431 11074 9980 9749 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00430 9749 9743 9744 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00429 9745 9760 9749 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00428 9759 11076 9761 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00427 9762 10709 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00426 9760 10708 9759 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00425 9682 9692 9683 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00424 9683 9680 9682 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00423 11074 9678 9681 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00422 10381 11075 10379 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00421 10380 10378 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00420 10702 10686 10381 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00419 7200 9716 7198 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00418 7199 10704 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00417 7201 9747 7200 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00416 5204 5771 5205 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00415 5203 5202 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00414 5556 8092 5204 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00413 4507 5727 4510 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00412 4511 5728 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00411 4508 10231 4507 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00410 5391 7711 5390 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00409 5392 9309 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00408 5394 8921 5393 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00407 5539 7652 5395 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00406 9866 10709 9865 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00405 9867 10073 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00404 9971 10686 9866 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00403 5209 9609 5208 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00402 5210 5207 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00401 5212 5214 5211 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00400 10892 8092 5206 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00399 4018 10031 4017 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00398 4019 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00397 4021 6277 4020 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00396 4183 8643 4022 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00395 10913 10909 10910 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00394 11074 10915 10916 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00393 10911 10916 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00392 5956 6197 6967 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00391 11074 6200 5957 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00390 5958 6201 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00389 6967 6198 5959 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00388 5960 6201 6197 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00387 6198 6200 5955 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00386 6217 7448 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00385 11074 10604 6217 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00384 6217 10892 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00383 11074 6132 6217 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00382 6131 6217 5990 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00381 7171 9433 7170 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00380 7172 8453 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00379 7174 8052 7173 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00378 7176 9716 7175 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00377 6044 6276 6048 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00376 6049 6278 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00375 6046 6275 6045 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00374 6280 6277 6047 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00373 9899 10789 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00372 9938 10774 9900 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00371 6820 8318 6664 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00370 6664 8316 6820 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00369 11074 6819 6663 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00368 6419 8122 6418 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00367 6421 6992 6420 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00366 11074 7655 6422 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00365 6784 6420 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00364 8097 10604 7886 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00363 7886 8091 8097 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00362 11074 9313 7885 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00361 4710 4708 4709 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00360 4709 6560 4710 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00359 11074 5293 4707 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00358 10894 10901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00357 10896 10915 10895 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00356 11074 6243 3997 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00355 3998 4666 3999 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00354 4003 3999 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00353 4541 4538 6778 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00352 11074 4539 4542 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00351 4544 4543 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00350 6778 4540 4545 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00349 4409 4543 4538 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00348 4540 4539 4408 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00347 11074 11026 10685 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00346 10708 10685 10486 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00345 11074 10685 10708 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00344 11074 10685 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00343 11024 10685 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00342 11074 11026 10681 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00341 10700 10681 10485 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00340 11074 10681 10700 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00339 11074 10681 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00338 11024 10681 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00337 11074 11026 11027 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00336 11072 11027 11025 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00335 11074 11027 11072 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00334 11074 11027 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00333 11024 11027 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00332 11074 11026 10688 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00331 10686 10688 10487 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00330 11074 10688 10686 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00329 11074 10688 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00328 11024 10688 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00327 11074 7766 7768 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00326 11026 7768 7767 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00325 11074 7768 11026 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00324 11074 7768 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00323 11024 7768 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00322 4703 5873 4702 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00321 4705 4701 4704 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00320 11074 4700 4706 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00319 5014 4704 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00318 4032 5293 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00317 4354 4038 4033 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00316 4034 6278 4354 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00315 11074 4030 4034 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00314 4034 4031 11074 11074 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00313 11074 1556 607 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00312 608 1881 758 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00311 759 758 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00310 2682 2680 2683 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00309 2683 2681 2682 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00308 11074 2688 2683 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00307 2997 2682 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00306 11074 1314 768 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00305 7514 768 624 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00304 11074 768 7514 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00303 11074 768 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00302 11024 768 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00301 11074 1314 1315 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00300 8126 1315 1192 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00299 11074 1315 8126 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00298 11074 1315 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00297 11024 1315 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00296 11074 773 772 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00295 1314 772 628 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00294 11074 772 1314 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00293 11074 772 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00292 11024 772 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00291 11074 508 504 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00290 7721 504 503 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00289 11074 504 7721 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00288 11074 504 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00287 11024 504 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00286 11074 508 506 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00285 7478 506 505 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00284 11074 506 7478 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00283 11074 506 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00282 11024 506 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00281 11074 510 509 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00280 508 509 507 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00279 11074 509 508 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00278 11074 509 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00277 11024 509 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00276 11074 8662 8663 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00275 10027 8663 8536 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00274 11074 8663 10027 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00273 11074 8663 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00272 11024 8663 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00271 11074 8662 8656 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00270 9582 8656 8525 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00269 11074 8656 9582 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00268 11074 8656 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00267 11024 8656 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00266 11074 8100 8099 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00265 8662 8099 7897 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00264 11074 8099 8662 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00263 11074 8099 11024 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00262 11024 8099 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00261 7472 7475 7290 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00260 7290 7690 7472 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00259 11074 9624 7290 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00258 7471 7472 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00257 4795 5214 4797 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00256 4798 9609 4978 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00255 11074 8092 4796 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00254 7690 4978 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00253 2168 1886 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00252 11074 1884 2168 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00251 6738 6901 6737 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00250 6739 7540 6903 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00249 11074 6902 6740 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00248 6900 6903 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00247 2149 2776 2148 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00246 2150 2158 2152 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00245 11074 2147 2151 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00244 4333 2152 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00243 5759 5756 5758 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00242 5760 5757 5762 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00241 11074 6141 5761 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00240 5755 5762 11074 11074 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00239 3952 8297 3953 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00238 11074 10915 3954 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00237 3951 3954 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00236 6398 6396 6401 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00235 11074 6394 6395 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00234 6399 6402 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00233 6401 6397 6400 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00232 6317 6402 6396 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00231 6397 6394 6316 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00230 1172 5600 1171 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00229 1175 8661 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00228 1174 6275 1173 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00227 1884 1304 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00226 1304 1170 1174 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00225 1124 1277 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00224 1121 1278 1276 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00223 1120 1279 1272 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00222 11074 1493 1120 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00221 11074 5262 1279 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00220 1278 1279 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00219 11074 1280 1277 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00218 1276 1279 1124 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00217 1122 1276 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00216 11074 1274 1123 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00215 1272 1278 1274 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00214 1493 1272 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00213 11074 1272 1493 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00212 11074 8388 8038 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00211 8038 8411 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00210 7920 9033 8038 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00209 10607 10608 10452 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00208 10452 10606 10607 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00207 11074 10880 10452 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00206 10605 10607 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00205 1604 5600 1608 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00204 1609 5901 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00203 1606 7711 1605 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00202 1899 1607 11074 11074 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00201 1607 1603 1606 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00200 2213 2211 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00199 11074 2212 2213 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00198 11074 5023 4478 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00197 4478 5037 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00196 4477 4476 4478 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00195 6521 6522 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00194 6354 6357 6356 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00193 6352 6523 6520 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00192 11074 6527 6352 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00191 11074 8048 6523 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00190 6357 6523 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00189 11074 6530 6522 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00188 6356 6523 6521 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00187 6351 6356 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00186 11074 6353 6355 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00185 6520 6357 6353 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00184 6527 6520 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00183 11074 6520 6527 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00182 6496 6493 6495 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00181 6495 8713 6496 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00180 11074 8709 6494 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00179 5821 6152 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00178 5829 6151 5822 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00177 7972 10399 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00176 8430 8746 7971 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00175 7366 10399 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00174 8426 9080 7367 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00173 10469 10637 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00172 10467 10639 10635 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00171 10465 10640 10631 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00170 11074 10924 10465 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00169 11074 10638 10640 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00168 10639 10640 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00167 11074 10923 10637 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00166 10635 10640 10469 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00165 10466 10635 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00164 11074 10634 10468 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00163 10631 10639 10634 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00162 10924 10631 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00161 11074 10631 10924 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00160 10225 10614 10227 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00159 10227 10615 10225 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00158 11074 11018 10226 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00157 7057 10027 7055 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00156 7056 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00155 7058 7466 7057 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00154 6098 6518 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00153 6151 6819 6099 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00152 8236 11066 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00151 9029 10689 8237 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00150 612 9020 613 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00149 614 2133 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00148 7042 5918 612 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00147 1744 9314 1742 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00146 1743 2133 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00145 6220 5918 1744 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00144 4058 3728 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00143 11074 4037 4058 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00142 4058 4023 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00141 11074 3726 4058 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00140 447 4995 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00139 449 1545 448 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00138 72 482 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00137 213 219 73 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00136 4141 5181 4140 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00135 11074 4324 4553 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00134 11074 5181 4143 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00133 4138 4628 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00132 4139 4247 4138 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00131 4137 4975 4141 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00130 4553 4324 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00129 4639 5181 4638 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00128 11074 4634 6213 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00127 11074 5181 4642 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00126 4641 4640 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00125 4636 4635 4641 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00124 4637 7085 4639 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00123 6213 4634 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00122 4623 5181 4627 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00121 11074 4615 4617 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00120 11074 5181 4630 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00119 4629 4628 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00118 4622 4621 4629 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00117 4624 5562 4623 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00116 4617 4615 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00115 7604 9582 7602 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00114 7603 10036 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00113 7600 7601 7604 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00112 7358 7529 11074 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00111 7526 7805 7359 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00110 1728 9020 1727 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00109 1729 5600 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00108 2099 9308 1728 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00107 11074 1991 1994 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00106 1992 6978 1995 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00105 1993 1995 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00104 11074 3822 3436 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00103 3435 4926 3616 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00102 3615 3616 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00101 11074 4929 4548 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00100 4546 5150 4547 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00099 4920 4936 4757 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_00098 4547 4917 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00097 4756 4929 4917 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_00096 5518 4922 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_00095 4558 4919 4549 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00094 4551 4936 4550 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00093 4552 4920 4556 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00092 4557 6128 4558 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00091 11074 4929 4570 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00090 4568 5527 4569 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00089 4933 4936 4760 11074 sg13_lv_nmos L=0.13U W=0.62U AS=0.1488P AD=0.1488P PS=1.72U PD=1.72U 
Mtr_00088 4569 4930 11074 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00087 4759 4929 4930 11074 sg13_lv_nmos L=0.13U W=0.47U AS=0.1128P AD=0.1128P PS=1.42U PD=1.42U 
Mtr_00086 5681 4934 11074 11074 sg13_lv_nmos L=0.13U W=2.04U AS=0.4896P AD=0.4896P PS=4.57U PD=4.57U 
Mtr_00085 4582 4932 4571 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00084 4573 4936 4572 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00083 4574 4933 4580 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00082 4581 5148 4582 11074 sg13_lv_nmos L=0.13U W=0.92U AS=0.2208P AD=0.2208P PS=2.32U PD=2.32U 
Mtr_00081 10821 10819 11074 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00080 10816 10822 10820 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00079 10814 10823 10813 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00078 11074 10825 10814 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00077 11074 10914 10823 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00076 10822 10823 11074 11074 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00075 11074 10824 10819 11074 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00074 10820 10823 10821 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00073 10817 10820 11074 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00072 11074 10815 10818 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00071 10813 10822 10815 11074 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00070 10825 10813 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00069 11074 10813 10825 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00068 9296 7448 7266 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00067 7266 7463 9296 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00066 11074 7447 7265 11074 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00065 11074 6220 2896 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00064 2897 3057 3049 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00063 3331 3049 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00062 10076 11067 9875 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00061 9875 10408 10076 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00060 11074 10399 9875 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00059 9977 10076 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00058 8965 9379 8963 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00057 11074 8962 9355 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00056 11074 9379 8967 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00055 8968 9095 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00054 8964 8969 8968 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00053 8966 9350 8965 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00052 9355 8962 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00051 9195 9379 9193 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00050 11074 9377 9375 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00049 11074 9379 9197 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00048 9198 9958 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00047 9194 9381 9198 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00046 9196 9376 9195 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00045 9375 9377 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00044 9008 9379 9010 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00043 11074 9004 9006 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00042 11074 9379 9014 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00041 9011 9051 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00040 9012 9015 9011 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00039 9009 9007 9008 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00038 9006 9004 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00037 101 6241 99 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00036 11074 233 231 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00035 11074 6241 103 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00034 104 241 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00033 100 235 104 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00032 102 6243 101 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00031 231 233 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00030 9222 10684 9219 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00029 11074 9413 9412 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00028 11074 10684 9224 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00027 9220 9509 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00026 9221 9416 9220 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00025 9223 9701 9222 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00024 9412 9413 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00023 9858 10684 9857 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00022 11074 10062 10710 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00021 11074 10684 9859 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00020 9855 10594 11074 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00019 9856 9967 9855 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00018 9854 10350 9858 11074 sg13_lv_nmos L=0.13U W=0.69U AS=0.1656P AD=0.1656P PS=1.87U PD=1.87U 
Mtr_00017 10710 10062 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00016 2723 7711 2724 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00015 2725 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00014 6221 9597 2723 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00013 1153 7514 1154 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00012 1155 5919 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00011 7041 9597 1153 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00010 11074 10018 9134 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00009 9135 9306 9303 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00008 9533 9303 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00007 2641 2982 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00006 2640 3625 2641 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00005 11074 3632 2640 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00004 3457 3871 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00003 3633 4535 3456 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00002 11074 3632 3633 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00001 3849 3633 11074 11074 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
.ends arlet6502_cts_r

