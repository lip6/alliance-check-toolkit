* GuardRing_N18000W13312HFF
* GuardRing_N18000W13312HFF
.subckt GuardRing_N18000W13312HFF conn

.ends GuardRing_N18000W13312HFF
