* tie_diff
* tie_diff
.subckt tie_diff vdd vss

.ends tie_diff
