-- no model for nand2_x0
