* diode_ff
.param
+ sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult = 8.4794e-01    
+ sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult = 9.3896e-01    
+ sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult = 7.9633e-01  
+ sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult = 7.7428e-01 
+ sky130_fd_pr__nfet_01v8__ajunction_mult = 8.4039e-1
+ sky130_fd_pr__nfet_01v8__pjunction_mult = 8.6147e-1
+ sky130_fd_pr__pfet_01v8__ajunction_mult = 0.93001
+ sky130_fd_pr__pfet_01v8__pjunction_mult = 0.93439
