* Gallery
* nand3_x0
.subckt nand3_x0 vdd vss nq i0 i1 i2
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net0 i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos _net1 i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nand3_x0
* nand3_x1
.subckt nand3_x1 vdd vss nq i0 i1 i2
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi1_nmos _net0 i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi2_nmos _net1 i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi2_pmos vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends nand3_x1
* nand2_x1
.subckt nand2_x1 vdd vss nq i0 i1
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi1_nmos _net0 i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends nand2_x1
* nand4_x0
.subckt nand4_x0 vdd vss nq i0 i1 i2 i3
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net0 i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos _net1 i2 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi3_nmos _net2 i3 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi3_pmos nq i3 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nand4_x0
* nand2_x0
.subckt nand2_x0 vdd vss nq i0 i1
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net0 i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nand2_x0
* nand4_x1
.subckt nand4_x1 vdd vss nq i0 i1 i2 i3
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi1_nmos _net0 i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi2_nmos _net1 i2 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi2_pmos vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi3_nmos _net2 i3 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi3_pmos nq i3 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends nand4_x1
* buf_x4
.subckt buf_x4 vdd vss i q
Mstage0_nmos _i_n i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.195um
Mstage0_pmos _i_n i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.755um
Mnmos[0] vss _i_n q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.195um
Mpmos[0] vdd _i_n q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.755um
Mnmos[1] q _i_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.195um
Mpmos[1] q _i_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.755um
Mnmos[2] vss _i_n q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.195um
Mpmos[2] vdd _i_n q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.755um
Mnmos[3] q _i_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.195um
Mpmos[3] q _i_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.755um
.ends buf_x4
* and2_x1
.subckt and2_x1 vdd vss q i0 i1
Mi0_nmos nq i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net0 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mn_pd vss nq q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mq_pu vdd nq q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends and2_x1
* buf_x2
.subckt buf_x2 vdd vss i q
Mstage0_nmos _i_n i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mstage0_pmos _i_n i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnmos[0] vss _i_n q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.195um
Mpmos[0] vdd _i_n q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.755um
Mnmos[1] q _i_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.195um
Mpmos[1] q _i_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.755um
.ends buf_x2
* and3_x1
.subckt and3_x1 vdd vss q i0 i1 i2
Mi0_nmos nq i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos nq i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net0 i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos vdd i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos _net1 i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos nq i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mn_pd vss nq q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mq_pu vdd nq q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends and3_x1
* buf_x1
.subckt buf_x1 vdd vss i q
Mstage0_nmos _i_n i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mstage0_pmos _i_n i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnmos vss _i_n q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.195um
Mpmos vdd _i_n q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.755um
.ends buf_x1
* and4_x1
.subckt and4_x1 vdd vss q i0 i1 i2 i3
Mi0_nmos nq i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net0 i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos _net1 i2 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi3_nmos _net2 i3 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi3_pmos nq i3 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mn_pd vss nq q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mq_pu vdd nq q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends and4_x1
* inv_x4
.subckt inv_x4 vdd vss i nq
Mnmos[0] vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mpmos[0] vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mnmos[1] nq i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mpmos[1] nq i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mnmos[2] vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mpmos[2] vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mnmos[3] nq i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mpmos[3] nq i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends inv_x4
* nor2_x0
.subckt nor2_x0 vdd vss nq i0 i1
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos _net0 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nor2_x0
* inv_x2
.subckt inv_x2 vdd vss i nq
Mnmos[0] vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mpmos[0] vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mnmos[1] nq i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mpmos[1] nq i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends inv_x2
* nor2_x1
.subckt nor2_x1 vdd vss nq i0 i1
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi0_pmos vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi1_pmos _net0 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends nor2_x1
* inv_x1
.subckt inv_x1 vdd vss i nq
Mnmos vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mpmos vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends inv_x1
* nor3_x0
.subckt nor3_x0 vdd vss nq i0 i1 i2
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos _net0 i1 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos vss i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos _net1 i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nor3_x0
* inv_x0
.subckt inv_x0 vdd vss i nq
Mnmos vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mpmos vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends inv_x0
* nor3_x1
.subckt nor3_x1 vdd vss nq i0 i1 i2
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi0_pmos vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi1_pmos _net0 i1 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi2_nmos vss i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi2_pmos _net1 i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends nor3_x1
* decap_w0
.subckt decap_w0 vdd vss
Mnpass vss one zero vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.465um
Mppass one zero vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.025um
.ends decap_w0
* nor4_x0
.subckt nor4_x0 vdd vss nq i0 i1 i2 i3
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos _net0 i1 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos vss i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos _net1 i2 _net2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi3_nmos nq i3 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi3_pmos _net2 i3 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nor4_x0
* zeroone_x1
.subckt zeroone_x1 vdd vss one zero
Mnpass vss one zero vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.465um
Mppass one zero vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.025um
.ends zeroone_x1
* nor4_x1
.subckt nor4_x1 vdd vss nq i0 i1 i2 i3
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi0_pmos vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi1_pmos _net0 i1 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi2_nmos vss i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi2_pmos _net1 i2 _net2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi3_nmos nq i3 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi3_pmos _net2 i3 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends nor4_x1
* one_x1
.subckt one_x1 vdd vss one
Mnpass vss one zero vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.465um
Mppass one zero vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.025um
.ends one_x1
* or2_x1
.subckt or2_x1 vdd vss q i0 i1
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos nq i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos _net0 i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mn_pd vss nq q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mq_pu vdd nq q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends or2_x1
* zero_x1
.subckt zero_x1 vdd vss zero
Mnpass vss one zero vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.465um
Mppass one zero vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.025um
.ends zero_x1
* or3_x1
.subckt or3_x1 vdd vss q i0 i1 i2
Mi0_nmos nq i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos nq i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos vss i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos _net0 i1 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos nq i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos _net1 i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mn_pd vss nq q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mq_pu vdd nq q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends or3_x1
* diode_w1
.subckt diode_w1 vdd vss i

.ends diode_w1
* or4_x1
.subckt or4_x1 vdd vss q i0 i1 i2 i3
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos nq i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos _net0 i1 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos vss i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos _net1 i2 _net2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi3_nmos nq i3 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi3_pmos _net2 i3 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mn_pd vss nq q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mq_pu vdd nq q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends or4_x1
* tie_poly_w4
.subckt tie_poly_w4 vdd vss

.ends tie_poly_w4
* mux2_x1
.subckt mux2_x1 vdd vss i0 i1 cmd q
Mcmd_inv_nmos cmd_n cmd vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mcmd_inv_pmos cmd_n cmd vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mcmd_n_npass _net0 cmd_n _q_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mcmd_ppass _net1 cmd _q_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mcmd_npass _q_n cmd _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mcmd_n_ppass _q_n cmd_n _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net2 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos _net3 i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mq_n_inv_nmos vss _q_n q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.195um
Mq_n_inv_pmos vdd _q_n q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.755um
.ends mux2_x1
* tie_diff_w4
.subckt tie_diff_w4 vdd vss

.ends tie_diff_w4
* and21nor_x0
.subckt and21nor_x0 vdd vss nq i0 i1 i2
Mi0_nmos vss i0 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos _net0 i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net1 i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos vdd i1 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos nq i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos _net0 i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends and21nor_x0
* tie_w4
.subckt tie_w4 vdd vss

.ends tie_w4
* and21nor_x1
.subckt and21nor_x1 vdd vss nq i0 i1 i2
Mi0_nmos vss i0 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi0_pmos _net0 i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi1_nmos _net1 i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi1_pmos vdd i1 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi2_nmos nq i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi2_pmos _net0 i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends and21nor_x1
* fill_w4
.subckt fill_w4 vdd vss

.ends fill_w4
* or21nand_x0
.subckt or21nand_x0 vdd vss nq i0 i1 i2
Mi0_nmos _net0 i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos vss i1 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos _net1 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi2_nmos _net0 i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi2_pmos nq i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends or21nand_x0
* tie_poly_w2
.subckt tie_poly_w2 vdd vss

.ends tie_poly_w2
* or21nand_x1
.subckt or21nand_x1 vdd vss nq i0 i1 i2
Mi0_nmos _net0 i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi0_pmos vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi1_nmos vss i1 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi1_pmos _net1 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mi2_nmos _net0 i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mi2_pmos nq i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends or21nand_x1
* tie_diff_w2
.subckt tie_diff_w2 vdd vss

.ends tie_diff_w2
* xor2_x0
.subckt xor2_x0 vdd vss i0 i1 q
Mi0_nmos0 i0_n i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos0 i0_n i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi0_nmos1 vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos1 vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos0 _net0 i1 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_n_pmos _net1 i1_n q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi0_n_nmos q i0_n _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_n_pmos q i0_n _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_n_nmos _net2 i1_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos0 _net1 i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos1 vss i1 i1_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos1 vdd i1 i1_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends xor2_x0
* tie_w2
.subckt tie_w2 vdd vss

.ends tie_w2
* nexor2_x0
.subckt nexor2_x0 vdd vss i0 i1 nq
Mi0_nmos0 i0_n i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos0 i0_n i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi0_nmos1 vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos1 vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_n_nmos _net0 i1_n nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos0 _net1 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi0_n_nmos nq i0_n _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_n_pmos nq i0_n _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos0 _net2 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_n_pmos _net1 i1_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos1 vss i1 i1_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos1 vdd i1 i1_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nexor2_x0
* fill_w2
.subckt fill_w2 vdd vss

.ends fill_w2
* nsnrlatch_x0
.subckt nsnrlatch_x0 vdd vss nset nrst q nq
Mnset_nmos q nset _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnset_pmos vdd nset q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnq_nmos _net0 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnq_pmos q q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mq_nmos vss q _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mq_pmos vdd q nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnrst_nmos _net1 nset nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnrst_pmos nq nset vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends nsnrlatch_x0
* tie_poly
.subckt tie_poly vdd vss

.ends tie_poly
* nsnrlatch_x1
.subckt nsnrlatch_x1 vdd vss nset nrst q nq
Mnset_nmos q nset _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.465um
Mnset_pmos vdd nset q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.025um
Mnq_nmos _net0 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.465um
Mnq_pmos q q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.025um
Mq_nmos vss q _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.465um
Mq_pmos vdd q nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.025um
Mnrst_nmos _net1 nset nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.465um
Mnrst_pmos nq nset vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.025um
.ends nsnrlatch_x1
* tie_diff
.subckt tie_diff vdd vss

.ends tie_diff
* dff_x1
.subckt dff_x1 vdd vss i clk q
Mclk_nmos _clk_n clk vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_pmos _clk_n clk vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_n_nmos0 vss _clk_n _clk_buf vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_pmos0 vdd _clk_n _clk_buf vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi_nmos _u i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi_pmos _u i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mu_nmos vss _u _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mu_pmos vdd _u _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_n_nmos1 _net0 _clk_n _dff_m vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_buf_pmos0 _net1 _clk_buf _dff_m vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_buf_nmos0 _dff_m _clk_buf _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_pmos1 _dff_m _clk_n _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
My_nmos _net2 _y vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
My_pmos _net3 _y vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mdff_m_nmos vss _dff_m _y vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mdff_m_pmos vdd _dff_m _y vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_buf_nmos1 _y _clk_buf _dff_s vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_pmos2 _y _clk_n _dff_s vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_n_nmos2 _dff_s _clk_n _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_buf_pmos1 _dff_s _clk_buf _net5 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mq_nmos _net4 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mq_pmos _net5 q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mdff_s_nmos vss _dff_s q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.925um
Mdff_s_pmos vdd _dff_s q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.485um
.ends dff_x1
* tie
.subckt tie vdd vss

.ends tie
* dffnr_x1
.subckt dffnr_x1 vdd vss i clk q nrst
Mclk_nmos _clk_n clk vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_pmos _clk_n clk vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_n_nmos0 vss _clk_n _clk_buf vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_pmos0 vdd _clk_n _clk_buf vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi_nmos _u i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi_pmos _u i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mu_nmos vss _u _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mu_pmos vdd _u _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_n_nmos1 _net0 _clk_n _dff_m vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_buf_pmos0 _net1 _clk_buf _dff_m vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_buf_nmos0 _dff_m _clk_buf _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_pmos1 _dff_m _clk_n _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
My_nmos _net2 _y vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
My_pmos _net3 _y vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mdff_m_nmos vss _dff_m _net6 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mdff_m_pmos vdd _dff_m _y vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnrst_nmos0 _net6 nrst _y vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnrst_pmos0 _y nrst vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnrst_pmos1 vdd nrst _net5 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_buf_nmos1 _y _clk_buf _dff_s vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_nmos2 _dff_s _clk_n _net7 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_pmos2 _y _clk_n _dff_s vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnrst_nmos1 _net7 nrst _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_buf_pmos1 _dff_s _clk_buf _net5 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mq_nmos _net4 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mq_pmos _net5 q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mdff_s_nmos vss _dff_s q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.925um
Mdff_s_pmos vdd _dff_s q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.485um
.ends dffnr_x1
* fill
.subckt fill vdd vss

.ends fill
* Gallery
.subckt Gallery vss vdd
Xfill[0] vdd vss fill
Xdffnr_x1[1] vdd vss dffnr_x1[1].[_InstanceNet[i], 'Gallery'] dffnr_x1[1].[_InstanceNet[clk], 'Gallery'] dffnr_x1[1].[_InstanceNet[q], 'Gallery'] dffnr_x1[1].[_InstanceNet[nrst], 'Gallery'] dffnr_x1
Xdffnr_x1[2] vdd vss dffnr_x1[2].[_InstanceNet[i], 'Gallery'] dffnr_x1[2].[_InstanceNet[clk], 'Gallery'] dffnr_x1[2].[_InstanceNet[q], 'Gallery'] dffnr_x1[2].[_InstanceNet[nrst], 'Gallery'] dffnr_x1
Xtie[0] vdd vss tie
Xdff_x1[1] vdd vss dff_x1[1].[_InstanceNet[i], 'Gallery'] dff_x1[1].[_InstanceNet[clk], 'Gallery'] dff_x1[1].[_InstanceNet[q], 'Gallery'] dff_x1
Xfill[2] vdd vss fill
Xtie_diff[0] vdd vss tie_diff
Xnsnrlatch_x1[1] vdd vss nsnrlatch_x1[1].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x1[1].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x1[1].[_InstanceNet[q], 'Gallery'] nsnrlatch_x1[1].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x1
Xdff_x1[2] vdd vss dff_x1[2].[_InstanceNet[i], 'Gallery'] dff_x1[2].[_InstanceNet[clk], 'Gallery'] dff_x1[2].[_InstanceNet[q], 'Gallery'] dff_x1
Xtie_poly[0] vdd vss tie_poly
Xnsnrlatch_x0[1] vdd vss nsnrlatch_x0[1].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x0[1].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x0[1].[_InstanceNet[q], 'Gallery'] nsnrlatch_x0[1].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x0
Xtie[2] vdd vss tie
Xfill_w2[0] vdd vss fill_w2
Xnexor2_x0[1] vdd vss nexor2_x0[1].[_InstanceNet[i0], 'Gallery'] nexor2_x0[1].[_InstanceNet[i1], 'Gallery'] nexor2_x0[1].[_InstanceNet[nq], 'Gallery'] nexor2_x0
Xnsnrlatch_x1[2] vdd vss nsnrlatch_x1[2].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x1[2].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x1[2].[_InstanceNet[q], 'Gallery'] nsnrlatch_x1[2].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x1
Xtie_w2[0] vdd vss tie_w2
Xxor2_x0[1] vdd vss xor2_x0[1].[_InstanceNet[i0], 'Gallery'] xor2_x0[1].[_InstanceNet[i1], 'Gallery'] xor2_x0[1].[_InstanceNet[q], 'Gallery'] xor2_x0
Xtie_diff[2] vdd vss tie_diff
Xtie_diff_w2[0] vdd vss tie_diff_w2
Xor21nand_x1[1] vdd vss or21nand_x1[1].[_InstanceNet[nq], 'Gallery'] or21nand_x1[1].[_InstanceNet[i0], 'Gallery'] or21nand_x1[1].[_InstanceNet[i1], 'Gallery'] or21nand_x1[1].[_InstanceNet[i2], 'Gallery'] or21nand_x1
Xnsnrlatch_x0[2] vdd vss nsnrlatch_x0[2].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x0[2].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x0[2].[_InstanceNet[q], 'Gallery'] nsnrlatch_x0[2].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x0
Xtie_poly_w2[0] vdd vss tie_poly_w2
Xor21nand_x0[1] vdd vss or21nand_x0[1].[_InstanceNet[nq], 'Gallery'] or21nand_x0[1].[_InstanceNet[i0], 'Gallery'] or21nand_x0[1].[_InstanceNet[i1], 'Gallery'] or21nand_x0[1].[_InstanceNet[i2], 'Gallery'] or21nand_x0
Xtie_poly[2] vdd vss tie_poly
Xfill_w4[0] vdd vss fill_w4
Xand21nor_x1[1] vdd vss and21nor_x1[1].[_InstanceNet[nq], 'Gallery'] and21nor_x1[1].[_InstanceNet[i0], 'Gallery'] and21nor_x1[1].[_InstanceNet[i1], 'Gallery'] and21nor_x1[1].[_InstanceNet[i2], 'Gallery'] and21nor_x1
Xnexor2_x0[2] vdd vss nexor2_x0[2].[_InstanceNet[i0], 'Gallery'] nexor2_x0[2].[_InstanceNet[i1], 'Gallery'] nexor2_x0[2].[_InstanceNet[nq], 'Gallery'] nexor2_x0
Xtie_w4[0] vdd vss tie_w4
Xand21nor_x0[1] vdd vss and21nor_x0[1].[_InstanceNet[nq], 'Gallery'] and21nor_x0[1].[_InstanceNet[i0], 'Gallery'] and21nor_x0[1].[_InstanceNet[i1], 'Gallery'] and21nor_x0[1].[_InstanceNet[i2], 'Gallery'] and21nor_x0
Xfill_w2[2] vdd vss fill_w2
Xtie_diff_w4[0] vdd vss tie_diff_w4
Xmux2_x1[1] vdd vss mux2_x1[1].[_InstanceNet[i0], 'Gallery'] mux2_x1[1].[_InstanceNet[i1], 'Gallery'] mux2_x1[1].[_InstanceNet[cmd], 'Gallery'] mux2_x1[1].[_InstanceNet[q], 'Gallery'] mux2_x1
Xxor2_x0[2] vdd vss xor2_x0[2].[_InstanceNet[i0], 'Gallery'] xor2_x0[2].[_InstanceNet[i1], 'Gallery'] xor2_x0[2].[_InstanceNet[q], 'Gallery'] xor2_x0
Xtie_poly_w4[0] vdd vss tie_poly_w4
Xor4_x1[1] vdd vss or4_x1[1].[_InstanceNet[q], 'Gallery'] or4_x1[1].[_InstanceNet[i0], 'Gallery'] or4_x1[1].[_InstanceNet[i1], 'Gallery'] or4_x1[1].[_InstanceNet[i2], 'Gallery'] or4_x1[1].[_InstanceNet[i3], 'Gallery'] or4_x1
Xtie_w2[2] vdd vss tie_w2
Xdiode_w1[0] vdd vss diode_w1[0].[_InstanceNet[i], 'Gallery'] diode_w1
Xor3_x1[1] vdd vss or3_x1[1].[_InstanceNet[q], 'Gallery'] or3_x1[1].[_InstanceNet[i0], 'Gallery'] or3_x1[1].[_InstanceNet[i1], 'Gallery'] or3_x1[1].[_InstanceNet[i2], 'Gallery'] or3_x1
Xor21nand_x1[2] vdd vss or21nand_x1[2].[_InstanceNet[nq], 'Gallery'] or21nand_x1[2].[_InstanceNet[i0], 'Gallery'] or21nand_x1[2].[_InstanceNet[i1], 'Gallery'] or21nand_x1[2].[_InstanceNet[i2], 'Gallery'] or21nand_x1
Xzero_x1[0] vdd vss zero_x1[0].[_InstanceNet[zero], 'Gallery'] zero_x1
Xor2_x1[1] vdd vss or2_x1[1].[_InstanceNet[q], 'Gallery'] or2_x1[1].[_InstanceNet[i0], 'Gallery'] or2_x1[1].[_InstanceNet[i1], 'Gallery'] or2_x1
Xtie_diff_w2[2] vdd vss tie_diff_w2
Xone_x1[0] vdd vss one_x1[0].[_InstanceNet[one], 'Gallery'] one_x1
Xnor4_x1[1] vdd vss nor4_x1[1].[_InstanceNet[nq], 'Gallery'] nor4_x1[1].[_InstanceNet[i0], 'Gallery'] nor4_x1[1].[_InstanceNet[i1], 'Gallery'] nor4_x1[1].[_InstanceNet[i2], 'Gallery'] nor4_x1[1].[_InstanceNet[i3], 'Gallery'] nor4_x1
Xor21nand_x0[2] vdd vss or21nand_x0[2].[_InstanceNet[nq], 'Gallery'] or21nand_x0[2].[_InstanceNet[i0], 'Gallery'] or21nand_x0[2].[_InstanceNet[i1], 'Gallery'] or21nand_x0[2].[_InstanceNet[i2], 'Gallery'] or21nand_x0
Xzeroone_x1[0] vdd vss zeroone_x1[0].[_InstanceNet[one], 'Gallery'] zeroone_x1[0].[_InstanceNet[zero], 'Gallery'] zeroone_x1
Xnor4_x0[1] vdd vss nor4_x0[1].[_InstanceNet[nq], 'Gallery'] nor4_x0[1].[_InstanceNet[i0], 'Gallery'] nor4_x0[1].[_InstanceNet[i1], 'Gallery'] nor4_x0[1].[_InstanceNet[i2], 'Gallery'] nor4_x0[1].[_InstanceNet[i3], 'Gallery'] nor4_x0
Xtie_poly_w2[2] vdd vss tie_poly_w2
Xdecap_w0[0] vdd vss decap_w0
Xnor3_x1[1] vdd vss nor3_x1[1].[_InstanceNet[nq], 'Gallery'] nor3_x1[1].[_InstanceNet[i0], 'Gallery'] nor3_x1[1].[_InstanceNet[i1], 'Gallery'] nor3_x1[1].[_InstanceNet[i2], 'Gallery'] nor3_x1
Xand21nor_x1[2] vdd vss and21nor_x1[2].[_InstanceNet[nq], 'Gallery'] and21nor_x1[2].[_InstanceNet[i0], 'Gallery'] and21nor_x1[2].[_InstanceNet[i1], 'Gallery'] and21nor_x1[2].[_InstanceNet[i2], 'Gallery'] and21nor_x1
Xinv_x0[0] vdd vss inv_x0[0].[_InstanceNet[i], 'Gallery'] inv_x0[0].[_InstanceNet[nq], 'Gallery'] inv_x0
Xnor3_x0[1] vdd vss nor3_x0[1].[_InstanceNet[nq], 'Gallery'] nor3_x0[1].[_InstanceNet[i0], 'Gallery'] nor3_x0[1].[_InstanceNet[i1], 'Gallery'] nor3_x0[1].[_InstanceNet[i2], 'Gallery'] nor3_x0
Xfill_w4[2] vdd vss fill_w4
Xinv_x1[0] vdd vss inv_x1[0].[_InstanceNet[i], 'Gallery'] inv_x1[0].[_InstanceNet[nq], 'Gallery'] inv_x1
Xnor2_x1[1] vdd vss nor2_x1[1].[_InstanceNet[nq], 'Gallery'] nor2_x1[1].[_InstanceNet[i0], 'Gallery'] nor2_x1[1].[_InstanceNet[i1], 'Gallery'] nor2_x1
Xand21nor_x0[2] vdd vss and21nor_x0[2].[_InstanceNet[nq], 'Gallery'] and21nor_x0[2].[_InstanceNet[i0], 'Gallery'] and21nor_x0[2].[_InstanceNet[i1], 'Gallery'] and21nor_x0[2].[_InstanceNet[i2], 'Gallery'] and21nor_x0
Xinv_x2[0] vdd vss inv_x2[0].[_InstanceNet[i], 'Gallery'] inv_x2[0].[_InstanceNet[nq], 'Gallery'] inv_x2
Xnor2_x0[1] vdd vss nor2_x0[1].[_InstanceNet[nq], 'Gallery'] nor2_x0[1].[_InstanceNet[i0], 'Gallery'] nor2_x0[1].[_InstanceNet[i1], 'Gallery'] nor2_x0
Xtie_w4[2] vdd vss tie_w4
Xinv_x4[0] vdd vss inv_x4[0].[_InstanceNet[i], 'Gallery'] inv_x4[0].[_InstanceNet[nq], 'Gallery'] inv_x4
Xand4_x1[1] vdd vss and4_x1[1].[_InstanceNet[q], 'Gallery'] and4_x1[1].[_InstanceNet[i0], 'Gallery'] and4_x1[1].[_InstanceNet[i1], 'Gallery'] and4_x1[1].[_InstanceNet[i2], 'Gallery'] and4_x1[1].[_InstanceNet[i3], 'Gallery'] and4_x1
Xmux2_x1[2] vdd vss mux2_x1[2].[_InstanceNet[i0], 'Gallery'] mux2_x1[2].[_InstanceNet[i1], 'Gallery'] mux2_x1[2].[_InstanceNet[cmd], 'Gallery'] mux2_x1[2].[_InstanceNet[q], 'Gallery'] mux2_x1
Xbuf_x1[0] vdd vss buf_x1[0].[_InstanceNet[i], 'Gallery'] buf_x1[0].[_InstanceNet[q], 'Gallery'] buf_x1
Xand3_x1[1] vdd vss and3_x1[1].[_InstanceNet[q], 'Gallery'] and3_x1[1].[_InstanceNet[i0], 'Gallery'] and3_x1[1].[_InstanceNet[i1], 'Gallery'] and3_x1[1].[_InstanceNet[i2], 'Gallery'] and3_x1
Xtie_diff_w4[2] vdd vss tie_diff_w4
Xbuf_x2[0] vdd vss buf_x2[0].[_InstanceNet[i], 'Gallery'] buf_x2[0].[_InstanceNet[q], 'Gallery'] buf_x2
Xand2_x1[1] vdd vss and2_x1[1].[_InstanceNet[q], 'Gallery'] and2_x1[1].[_InstanceNet[i0], 'Gallery'] and2_x1[1].[_InstanceNet[i1], 'Gallery'] and2_x1
Xor4_x1[2] vdd vss or4_x1[2].[_InstanceNet[q], 'Gallery'] or4_x1[2].[_InstanceNet[i0], 'Gallery'] or4_x1[2].[_InstanceNet[i1], 'Gallery'] or4_x1[2].[_InstanceNet[i2], 'Gallery'] or4_x1[2].[_InstanceNet[i3], 'Gallery'] or4_x1
Xbuf_x4[0] vdd vss buf_x4[0].[_InstanceNet[i], 'Gallery'] buf_x4[0].[_InstanceNet[q], 'Gallery'] buf_x4
Xnand4_x1[1] vdd vss nand4_x1[1].[_InstanceNet[nq], 'Gallery'] nand4_x1[1].[_InstanceNet[i0], 'Gallery'] nand4_x1[1].[_InstanceNet[i1], 'Gallery'] nand4_x1[1].[_InstanceNet[i2], 'Gallery'] nand4_x1[1].[_InstanceNet[i3], 'Gallery'] nand4_x1
Xtie_poly_w4[2] vdd vss tie_poly_w4
Xnand2_x0[0] vdd vss nand2_x0[0].[_InstanceNet[nq], 'Gallery'] nand2_x0[0].[_InstanceNet[i0], 'Gallery'] nand2_x0[0].[_InstanceNet[i1], 'Gallery'] nand2_x0
Xnand4_x0[1] vdd vss nand4_x0[1].[_InstanceNet[nq], 'Gallery'] nand4_x0[1].[_InstanceNet[i0], 'Gallery'] nand4_x0[1].[_InstanceNet[i1], 'Gallery'] nand4_x0[1].[_InstanceNet[i2], 'Gallery'] nand4_x0[1].[_InstanceNet[i3], 'Gallery'] nand4_x0
Xor3_x1[2] vdd vss or3_x1[2].[_InstanceNet[q], 'Gallery'] or3_x1[2].[_InstanceNet[i0], 'Gallery'] or3_x1[2].[_InstanceNet[i1], 'Gallery'] or3_x1[2].[_InstanceNet[i2], 'Gallery'] or3_x1
Xnand2_x1[0] vdd vss nand2_x1[0].[_InstanceNet[nq], 'Gallery'] nand2_x1[0].[_InstanceNet[i0], 'Gallery'] nand2_x1[0].[_InstanceNet[i1], 'Gallery'] nand2_x1
Xnand3_x1[1] vdd vss nand3_x1[1].[_InstanceNet[nq], 'Gallery'] nand3_x1[1].[_InstanceNet[i0], 'Gallery'] nand3_x1[1].[_InstanceNet[i1], 'Gallery'] nand3_x1[1].[_InstanceNet[i2], 'Gallery'] nand3_x1
Xdiode_w1[2] vdd vss diode_w1[2].[_InstanceNet[i], 'Gallery'] diode_w1
Xnand3_x0[0] vdd vss nand3_x0[0].[_InstanceNet[nq], 'Gallery'] nand3_x0[0].[_InstanceNet[i0], 'Gallery'] nand3_x0[0].[_InstanceNet[i1], 'Gallery'] nand3_x0[0].[_InstanceNet[i2], 'Gallery'] nand3_x0
Xnand3_x0[1] vdd vss nand3_x0[1].[_InstanceNet[nq], 'Gallery'] nand3_x0[1].[_InstanceNet[i0], 'Gallery'] nand3_x0[1].[_InstanceNet[i1], 'Gallery'] nand3_x0[1].[_InstanceNet[i2], 'Gallery'] nand3_x0
Xor2_x1[2] vdd vss or2_x1[2].[_InstanceNet[q], 'Gallery'] or2_x1[2].[_InstanceNet[i0], 'Gallery'] or2_x1[2].[_InstanceNet[i1], 'Gallery'] or2_x1
Xnand3_x1[0] vdd vss nand3_x1[0].[_InstanceNet[nq], 'Gallery'] nand3_x1[0].[_InstanceNet[i0], 'Gallery'] nand3_x1[0].[_InstanceNet[i1], 'Gallery'] nand3_x1[0].[_InstanceNet[i2], 'Gallery'] nand3_x1
Xnand2_x1[1] vdd vss nand2_x1[1].[_InstanceNet[nq], 'Gallery'] nand2_x1[1].[_InstanceNet[i0], 'Gallery'] nand2_x1[1].[_InstanceNet[i1], 'Gallery'] nand2_x1
Xzero_x1[2] vdd vss zero_x1[2].[_InstanceNet[zero], 'Gallery'] zero_x1
Xnand4_x0[0] vdd vss nand4_x0[0].[_InstanceNet[nq], 'Gallery'] nand4_x0[0].[_InstanceNet[i0], 'Gallery'] nand4_x0[0].[_InstanceNet[i1], 'Gallery'] nand4_x0[0].[_InstanceNet[i2], 'Gallery'] nand4_x0[0].[_InstanceNet[i3], 'Gallery'] nand4_x0
Xnand2_x0[1] vdd vss nand2_x0[1].[_InstanceNet[nq], 'Gallery'] nand2_x0[1].[_InstanceNet[i0], 'Gallery'] nand2_x0[1].[_InstanceNet[i1], 'Gallery'] nand2_x0
Xnor4_x1[2] vdd vss nor4_x1[2].[_InstanceNet[nq], 'Gallery'] nor4_x1[2].[_InstanceNet[i0], 'Gallery'] nor4_x1[2].[_InstanceNet[i1], 'Gallery'] nor4_x1[2].[_InstanceNet[i2], 'Gallery'] nor4_x1[2].[_InstanceNet[i3], 'Gallery'] nor4_x1
Xnand4_x1[0] vdd vss nand4_x1[0].[_InstanceNet[nq], 'Gallery'] nand4_x1[0].[_InstanceNet[i0], 'Gallery'] nand4_x1[0].[_InstanceNet[i1], 'Gallery'] nand4_x1[0].[_InstanceNet[i2], 'Gallery'] nand4_x1[0].[_InstanceNet[i3], 'Gallery'] nand4_x1
Xbuf_x4[1] vdd vss buf_x4[1].[_InstanceNet[i], 'Gallery'] buf_x4[1].[_InstanceNet[q], 'Gallery'] buf_x4
Xone_x1[2] vdd vss one_x1[2].[_InstanceNet[one], 'Gallery'] one_x1
Xand2_x1[0] vdd vss and2_x1[0].[_InstanceNet[q], 'Gallery'] and2_x1[0].[_InstanceNet[i0], 'Gallery'] and2_x1[0].[_InstanceNet[i1], 'Gallery'] and2_x1
Xbuf_x2[1] vdd vss buf_x2[1].[_InstanceNet[i], 'Gallery'] buf_x2[1].[_InstanceNet[q], 'Gallery'] buf_x2
Xnor4_x0[2] vdd vss nor4_x0[2].[_InstanceNet[nq], 'Gallery'] nor4_x0[2].[_InstanceNet[i0], 'Gallery'] nor4_x0[2].[_InstanceNet[i1], 'Gallery'] nor4_x0[2].[_InstanceNet[i2], 'Gallery'] nor4_x0[2].[_InstanceNet[i3], 'Gallery'] nor4_x0
Xand3_x1[0] vdd vss and3_x1[0].[_InstanceNet[q], 'Gallery'] and3_x1[0].[_InstanceNet[i0], 'Gallery'] and3_x1[0].[_InstanceNet[i1], 'Gallery'] and3_x1[0].[_InstanceNet[i2], 'Gallery'] and3_x1
Xbuf_x1[1] vdd vss buf_x1[1].[_InstanceNet[i], 'Gallery'] buf_x1[1].[_InstanceNet[q], 'Gallery'] buf_x1
Xzeroone_x1[2] vdd vss zeroone_x1[2].[_InstanceNet[one], 'Gallery'] zeroone_x1[2].[_InstanceNet[zero], 'Gallery'] zeroone_x1
Xand4_x1[0] vdd vss and4_x1[0].[_InstanceNet[q], 'Gallery'] and4_x1[0].[_InstanceNet[i0], 'Gallery'] and4_x1[0].[_InstanceNet[i1], 'Gallery'] and4_x1[0].[_InstanceNet[i2], 'Gallery'] and4_x1[0].[_InstanceNet[i3], 'Gallery'] and4_x1
Xinv_x4[1] vdd vss inv_x4[1].[_InstanceNet[i], 'Gallery'] inv_x4[1].[_InstanceNet[nq], 'Gallery'] inv_x4
Xnor3_x1[2] vdd vss nor3_x1[2].[_InstanceNet[nq], 'Gallery'] nor3_x1[2].[_InstanceNet[i0], 'Gallery'] nor3_x1[2].[_InstanceNet[i1], 'Gallery'] nor3_x1[2].[_InstanceNet[i2], 'Gallery'] nor3_x1
Xnor2_x0[0] vdd vss nor2_x0[0].[_InstanceNet[nq], 'Gallery'] nor2_x0[0].[_InstanceNet[i0], 'Gallery'] nor2_x0[0].[_InstanceNet[i1], 'Gallery'] nor2_x0
Xinv_x2[1] vdd vss inv_x2[1].[_InstanceNet[i], 'Gallery'] inv_x2[1].[_InstanceNet[nq], 'Gallery'] inv_x2
Xdecap_w0[2] vdd vss decap_w0
Xnor2_x1[0] vdd vss nor2_x1[0].[_InstanceNet[nq], 'Gallery'] nor2_x1[0].[_InstanceNet[i0], 'Gallery'] nor2_x1[0].[_InstanceNet[i1], 'Gallery'] nor2_x1
Xinv_x1[1] vdd vss inv_x1[1].[_InstanceNet[i], 'Gallery'] inv_x1[1].[_InstanceNet[nq], 'Gallery'] inv_x1
Xnor3_x0[2] vdd vss nor3_x0[2].[_InstanceNet[nq], 'Gallery'] nor3_x0[2].[_InstanceNet[i0], 'Gallery'] nor3_x0[2].[_InstanceNet[i1], 'Gallery'] nor3_x0[2].[_InstanceNet[i2], 'Gallery'] nor3_x0
Xnor3_x0[0] vdd vss nor3_x0[0].[_InstanceNet[nq], 'Gallery'] nor3_x0[0].[_InstanceNet[i0], 'Gallery'] nor3_x0[0].[_InstanceNet[i1], 'Gallery'] nor3_x0[0].[_InstanceNet[i2], 'Gallery'] nor3_x0
Xinv_x0[1] vdd vss inv_x0[1].[_InstanceNet[i], 'Gallery'] inv_x0[1].[_InstanceNet[nq], 'Gallery'] inv_x0
Xinv_x0[2] vdd vss inv_x0[2].[_InstanceNet[i], 'Gallery'] inv_x0[2].[_InstanceNet[nq], 'Gallery'] inv_x0
Xnor3_x1[0] vdd vss nor3_x1[0].[_InstanceNet[nq], 'Gallery'] nor3_x1[0].[_InstanceNet[i0], 'Gallery'] nor3_x1[0].[_InstanceNet[i1], 'Gallery'] nor3_x1[0].[_InstanceNet[i2], 'Gallery'] nor3_x1
Xdecap_w0[1] vdd vss decap_w0
Xnor2_x1[2] vdd vss nor2_x1[2].[_InstanceNet[nq], 'Gallery'] nor2_x1[2].[_InstanceNet[i0], 'Gallery'] nor2_x1[2].[_InstanceNet[i1], 'Gallery'] nor2_x1
Xnor4_x0[0] vdd vss nor4_x0[0].[_InstanceNet[nq], 'Gallery'] nor4_x0[0].[_InstanceNet[i0], 'Gallery'] nor4_x0[0].[_InstanceNet[i1], 'Gallery'] nor4_x0[0].[_InstanceNet[i2], 'Gallery'] nor4_x0[0].[_InstanceNet[i3], 'Gallery'] nor4_x0
Xzeroone_x1[1] vdd vss zeroone_x1[1].[_InstanceNet[one], 'Gallery'] zeroone_x1[1].[_InstanceNet[zero], 'Gallery'] zeroone_x1
Xinv_x1[2] vdd vss inv_x1[2].[_InstanceNet[i], 'Gallery'] inv_x1[2].[_InstanceNet[nq], 'Gallery'] inv_x1
Xnor4_x1[0] vdd vss nor4_x1[0].[_InstanceNet[nq], 'Gallery'] nor4_x1[0].[_InstanceNet[i0], 'Gallery'] nor4_x1[0].[_InstanceNet[i1], 'Gallery'] nor4_x1[0].[_InstanceNet[i2], 'Gallery'] nor4_x1[0].[_InstanceNet[i3], 'Gallery'] nor4_x1
Xone_x1[1] vdd vss one_x1[1].[_InstanceNet[one], 'Gallery'] one_x1
Xnor2_x0[2] vdd vss nor2_x0[2].[_InstanceNet[nq], 'Gallery'] nor2_x0[2].[_InstanceNet[i0], 'Gallery'] nor2_x0[2].[_InstanceNet[i1], 'Gallery'] nor2_x0
Xor2_x1[0] vdd vss or2_x1[0].[_InstanceNet[q], 'Gallery'] or2_x1[0].[_InstanceNet[i0], 'Gallery'] or2_x1[0].[_InstanceNet[i1], 'Gallery'] or2_x1
Xzero_x1[1] vdd vss zero_x1[1].[_InstanceNet[zero], 'Gallery'] zero_x1
Xinv_x2[2] vdd vss inv_x2[2].[_InstanceNet[i], 'Gallery'] inv_x2[2].[_InstanceNet[nq], 'Gallery'] inv_x2
Xor3_x1[0] vdd vss or3_x1[0].[_InstanceNet[q], 'Gallery'] or3_x1[0].[_InstanceNet[i0], 'Gallery'] or3_x1[0].[_InstanceNet[i1], 'Gallery'] or3_x1[0].[_InstanceNet[i2], 'Gallery'] or3_x1
Xdiode_w1[1] vdd vss diode_w1[1].[_InstanceNet[i], 'Gallery'] diode_w1
Xand4_x1[2] vdd vss and4_x1[2].[_InstanceNet[q], 'Gallery'] and4_x1[2].[_InstanceNet[i0], 'Gallery'] and4_x1[2].[_InstanceNet[i1], 'Gallery'] and4_x1[2].[_InstanceNet[i2], 'Gallery'] and4_x1[2].[_InstanceNet[i3], 'Gallery'] and4_x1
Xor4_x1[0] vdd vss or4_x1[0].[_InstanceNet[q], 'Gallery'] or4_x1[0].[_InstanceNet[i0], 'Gallery'] or4_x1[0].[_InstanceNet[i1], 'Gallery'] or4_x1[0].[_InstanceNet[i2], 'Gallery'] or4_x1[0].[_InstanceNet[i3], 'Gallery'] or4_x1
Xtie_poly_w4[1] vdd vss tie_poly_w4
Xinv_x4[2] vdd vss inv_x4[2].[_InstanceNet[i], 'Gallery'] inv_x4[2].[_InstanceNet[nq], 'Gallery'] inv_x4
Xmux2_x1[0] vdd vss mux2_x1[0].[_InstanceNet[i0], 'Gallery'] mux2_x1[0].[_InstanceNet[i1], 'Gallery'] mux2_x1[0].[_InstanceNet[cmd], 'Gallery'] mux2_x1[0].[_InstanceNet[q], 'Gallery'] mux2_x1
Xtie_diff_w4[1] vdd vss tie_diff_w4
Xand3_x1[2] vdd vss and3_x1[2].[_InstanceNet[q], 'Gallery'] and3_x1[2].[_InstanceNet[i0], 'Gallery'] and3_x1[2].[_InstanceNet[i1], 'Gallery'] and3_x1[2].[_InstanceNet[i2], 'Gallery'] and3_x1
Xand21nor_x0[0] vdd vss and21nor_x0[0].[_InstanceNet[nq], 'Gallery'] and21nor_x0[0].[_InstanceNet[i0], 'Gallery'] and21nor_x0[0].[_InstanceNet[i1], 'Gallery'] and21nor_x0[0].[_InstanceNet[i2], 'Gallery'] and21nor_x0
Xtie_w4[1] vdd vss tie_w4
Xbuf_x1[2] vdd vss buf_x1[2].[_InstanceNet[i], 'Gallery'] buf_x1[2].[_InstanceNet[q], 'Gallery'] buf_x1
Xand21nor_x1[0] vdd vss and21nor_x1[0].[_InstanceNet[nq], 'Gallery'] and21nor_x1[0].[_InstanceNet[i0], 'Gallery'] and21nor_x1[0].[_InstanceNet[i1], 'Gallery'] and21nor_x1[0].[_InstanceNet[i2], 'Gallery'] and21nor_x1
Xfill_w4[1] vdd vss fill_w4
Xand2_x1[2] vdd vss and2_x1[2].[_InstanceNet[q], 'Gallery'] and2_x1[2].[_InstanceNet[i0], 'Gallery'] and2_x1[2].[_InstanceNet[i1], 'Gallery'] and2_x1
Xor21nand_x0[0] vdd vss or21nand_x0[0].[_InstanceNet[nq], 'Gallery'] or21nand_x0[0].[_InstanceNet[i0], 'Gallery'] or21nand_x0[0].[_InstanceNet[i1], 'Gallery'] or21nand_x0[0].[_InstanceNet[i2], 'Gallery'] or21nand_x0
Xtie_poly_w2[1] vdd vss tie_poly_w2
Xbuf_x2[2] vdd vss buf_x2[2].[_InstanceNet[i], 'Gallery'] buf_x2[2].[_InstanceNet[q], 'Gallery'] buf_x2
Xor21nand_x1[0] vdd vss or21nand_x1[0].[_InstanceNet[nq], 'Gallery'] or21nand_x1[0].[_InstanceNet[i0], 'Gallery'] or21nand_x1[0].[_InstanceNet[i1], 'Gallery'] or21nand_x1[0].[_InstanceNet[i2], 'Gallery'] or21nand_x1
Xtie_diff_w2[1] vdd vss tie_diff_w2
Xnand4_x1[2] vdd vss nand4_x1[2].[_InstanceNet[nq], 'Gallery'] nand4_x1[2].[_InstanceNet[i0], 'Gallery'] nand4_x1[2].[_InstanceNet[i1], 'Gallery'] nand4_x1[2].[_InstanceNet[i2], 'Gallery'] nand4_x1[2].[_InstanceNet[i3], 'Gallery'] nand4_x1
Xxor2_x0[0] vdd vss xor2_x0[0].[_InstanceNet[i0], 'Gallery'] xor2_x0[0].[_InstanceNet[i1], 'Gallery'] xor2_x0[0].[_InstanceNet[q], 'Gallery'] xor2_x0
Xtie_w2[1] vdd vss tie_w2
Xbuf_x4[2] vdd vss buf_x4[2].[_InstanceNet[i], 'Gallery'] buf_x4[2].[_InstanceNet[q], 'Gallery'] buf_x4
Xnexor2_x0[0] vdd vss nexor2_x0[0].[_InstanceNet[i0], 'Gallery'] nexor2_x0[0].[_InstanceNet[i1], 'Gallery'] nexor2_x0[0].[_InstanceNet[nq], 'Gallery'] nexor2_x0
Xfill_w2[1] vdd vss fill_w2
Xnand4_x0[2] vdd vss nand4_x0[2].[_InstanceNet[nq], 'Gallery'] nand4_x0[2].[_InstanceNet[i0], 'Gallery'] nand4_x0[2].[_InstanceNet[i1], 'Gallery'] nand4_x0[2].[_InstanceNet[i2], 'Gallery'] nand4_x0[2].[_InstanceNet[i3], 'Gallery'] nand4_x0
Xnsnrlatch_x0[0] vdd vss nsnrlatch_x0[0].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x0[0].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x0[0].[_InstanceNet[q], 'Gallery'] nsnrlatch_x0[0].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x0
Xtie_poly[1] vdd vss tie_poly
Xnand2_x0[2] vdd vss nand2_x0[2].[_InstanceNet[nq], 'Gallery'] nand2_x0[2].[_InstanceNet[i0], 'Gallery'] nand2_x0[2].[_InstanceNet[i1], 'Gallery'] nand2_x0
Xnsnrlatch_x1[0] vdd vss nsnrlatch_x1[0].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x1[0].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x1[0].[_InstanceNet[q], 'Gallery'] nsnrlatch_x1[0].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x1
Xtie_diff[1] vdd vss tie_diff
Xnand3_x1[2] vdd vss nand3_x1[2].[_InstanceNet[nq], 'Gallery'] nand3_x1[2].[_InstanceNet[i0], 'Gallery'] nand3_x1[2].[_InstanceNet[i1], 'Gallery'] nand3_x1[2].[_InstanceNet[i2], 'Gallery'] nand3_x1
Xdff_x1[0] vdd vss dff_x1[0].[_InstanceNet[i], 'Gallery'] dff_x1[0].[_InstanceNet[clk], 'Gallery'] dff_x1[0].[_InstanceNet[q], 'Gallery'] dff_x1
Xtie[1] vdd vss tie
Xnand2_x1[2] vdd vss nand2_x1[2].[_InstanceNet[nq], 'Gallery'] nand2_x1[2].[_InstanceNet[i0], 'Gallery'] nand2_x1[2].[_InstanceNet[i1], 'Gallery'] nand2_x1
Xdffnr_x1[0] vdd vss dffnr_x1[0].[_InstanceNet[i], 'Gallery'] dffnr_x1[0].[_InstanceNet[clk], 'Gallery'] dffnr_x1[0].[_InstanceNet[q], 'Gallery'] dffnr_x1[0].[_InstanceNet[nrst], 'Gallery'] dffnr_x1
Xfill[1] vdd vss fill
Xnand3_x0[2] vdd vss nand3_x0[2].[_InstanceNet[nq], 'Gallery'] nand3_x0[2].[_InstanceNet[i0], 'Gallery'] nand3_x0[2].[_InstanceNet[i1], 'Gallery'] nand3_x0[2].[_InstanceNet[i2], 'Gallery'] nand3_x0
.ends Gallery
