* Spice description of mx3_x2
* Spice driver version -455680229
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:46

* INTERF cmd0 cmd1 i0 i1 i2 q vdd vss 


.subckt mx3_x2 9 18 6 8 14 7 5 19 
* NET 5 = vdd
* NET 6 = i0
* NET 7 = q
* NET 8 = i1
* NET 9 = cmd0
* NET 14 = i2
* NET 18 = cmd1
* NET 19 = vss
Mtr_00020 7 15 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00019 5 9 10 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00018 4 14 3 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00017 15 18 4 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00016 2 13 15 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00015 3 8 2 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00014 5 10 3 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00013 1 9 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00012 15 6 1 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00011 13 18 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00010 7 15 19 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.29U AS=0.5496P AD=0.5496P PS=5.07U PD=5.07U 
Mtr_00009 19 9 10 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.51U AS=0.1224P AD=0.1224P PS=1.5U PD=1.5U 
Mtr_00008 11 10 19 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00007 13 18 19 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.68U AS=0.1632P AD=0.1632P PS=1.84U PD=1.84U 
Mtr_00006 15 6 11 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00005 19 9 17 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00004 17 8 12 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00003 15 13 16 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00002 16 14 17 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00001 12 18 15 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
C17 3 19 7.87036e-16
C15 5 19 3.997e-15
C14 6 19 1.98577e-15
C13 7 19 2.20321e-15
C12 8 19 1.39136e-15
C11 9 19 2.17007e-15
C10 10 19 1.82741e-15
C7 13 19 1.78155e-15
C6 14 19 1.08733e-15
C5 15 19 3.70347e-15
C3 17 19 7.71835e-16
C2 18 19 2.10758e-15
C1 19 19 3.81459e-15
.ends mx3_x2

