* Spice description of o4_x2
* Spice driver version 1933877019
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:24

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt o4_x2 7 8 6 9 5 2 10 
* NET 2 = vdd
* NET 5 = q
* NET 6 = i2
* NET 7 = i0
* NET 8 = i1
* NET 9 = i3
* NET 10 = vss
Mtr_00010 5 11 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 2 6 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00008 3 7 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00007 1 8 4 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00006 4 9 11 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00005 5 11 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 10 6 11 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00003 11 7 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 10 8 11 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 11 9 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C10 2 10 1.90796e-15
C7 5 10 2.15173e-15
C6 6 10 1.46564e-15
C5 7 10 1.52471e-15
C4 8 10 1.46995e-15
C3 9 10 1.7831e-15
C2 10 10 2.49738e-15
C1 11 10 2.99555e-15
.ends o4_x2

