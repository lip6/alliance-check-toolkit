sky130_fd_sc_hd__inv_1_3 with slope
*
* inv_1_3_hitas.spi
* sta compatible ngspice
* from simu/ngpice/top_sky130_fd_sc_hd__inv_1_3.spi

*****************

.TEMP 25

******************
******************
* BSIM4 transistor model parameters for ngspice included in db_ng.tcl
*
* nfet_01v8
*.include sky130_fd_pr__nfet_01v8__mismatch.corner.spice
*.include sky130_fd_pr__nfet_01v8__tt.corner.spice
* pfet_01v8_hvt
*.include sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
*.include sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice

*******************************

*******************************
*Simulation conditions

Vground evss 0 0
Vsupply evdd 0 DC 1.8
*gfoncd evdd 0 evdd 0 1.0e-15

******************
* circuit model
* include circuit netlist
.INCLUDE sky130_fd_sc_hd__inv_1_3.spi
*****************

*****************
* Circuit Instantiation
*.subckt sky130_fd_sc_hd__inv_1_3 in out vdd gnd
* 3 inverters loaded

Xinv_1_3 in out evdd evss sky130_fd_sc_hd__inv_1_3

.end

