*
* 

*****************

.TEMP 25

******************
* BSIM4 transistor model parameters for ngspice
*.lib /users/soft/analogdesign/scalable/techno/sky130_models_20220217/C4M.Sky130_all_lib.spice logic_tt 

*******************************
*Simulation conditions

Vground evss 0 0
Vsupply evdd 0 DC 1.8
*gfoncd evdd 0 evdd 0 1.0e-15

******************
* circuit model
* include circuit netlist
.include arlet6502_cts_r.spi
*****************

*****************
* Circuit Instantiation
*.subckt inv_x2 vdd vss i nq

Xc 2245 1706 1923 1547 1583 1361 3141 1351 2443 8237 8211 8186 8159 8133 8106 8082 4100 8118 8155 7383 6857 7083 6371 5620 4773 2365 1671 1370 1365 7309 6520 5614 4868 4312 1718 4160 3862 evdd evss 1424 arlet6502_cts_r
.end

