-- no model for nor3_x1
