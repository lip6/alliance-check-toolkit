* Spice description of gates
* Spice driver version 4677831
* Date ( dd/mm/yyyy hh:mm:ss ): 26/05/2017 at 19:09:16

* INTERF i[0] i[1] i[2] i[3] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] q[8] 
* INTERF q[9] q[10] q[11] q[12] q[13] vdd vss 

.INCLUDE rowend_x0.spi
.INCLUDE tie_x0.spi
.INCLUDE no3_x1.spi
.INCLUDE noa22_x1.spi
.INCLUDE no4_x1.spi
.INCLUDE na3_x1.spi
.INCLUDE na4_x1.spi
.INCLUDE an12_x1.spi
.INCLUDE nao22_x1.spi
.INCLUDE no2_x1.spi
.INCLUDE sff1_x4.spi
.INCLUDE inv_x1.spi
.INCLUDE na2_x1.spi
.INCLUDE xr2_x1.spi
.INCLUDE on12_x1.spi
.INCLUDE nxr2_x1.spi

.subckt gates 19 17 9 3 8 12 14 5 6 7 10 2 4 1 18 16 15 11 20 13 
* NET 1 = q[9]
* NET 2 = q[7]
* NET 3 = i[3]
* NET 4 = q[8]
* NET 5 = q[3]
* NET 6 = q[4]
* NET 7 = q[5]
* NET 8 = q[0]
* NET 9 = i[2]
* NET 10 = q[6]
* NET 11 = q[13]
* NET 12 = q[1]
* NET 13 = vss
* NET 14 = q[2]
* NET 15 = q[12]
* NET 16 = q[11]
* NET 17 = i[1]
* NET 18 = q[10]
* NET 19 = i[0]
* NET 20 = vdd
xtiex0_9 20 13 tie_x0
xtiex0_8 20 13 tie_x0
xtiex0_7 20 13 tie_x0
xtiex0_6 20 13 tie_x0
xtiex0_5 20 13 tie_x0
xtiex0_4 20 13 tie_x0
xrowendx0_3 20 13 rowend_x0
xtiex0_2 20 13 tie_x0
xtiex0_1 20 13 tie_x0
xg7 19 17 9 2 20 13 no3_x1
xg9 19 17 9 1 20 13 noa22_x1
xg8 19 17 9 3 4 20 13 no4_x1
xg3 19 17 9 5 20 13 na3_x1
xg4 19 17 9 3 6 20 13 na4_x1
xg0 19 17 8 20 13 an12_x1
xg5 19 17 9 7 20 13 nao22_x1
xg6 19 17 10 20 13 no2_x1
xg13 19 17 11 20 13 sff1_x4
xg1 19 12 20 13 inv_x1
xg2 19 17 14 20 13 na2_x1
xg12 19 17 15 20 13 xr2_x1
xg11 19 17 16 20 13 on12_x1
xg10 19 17 18 20 13 nxr2_x1
.ends gates

