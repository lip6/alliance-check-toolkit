* NGSPICE file created from picorv32.ext - technology: sky130A
* ouput form OpneLnae, further updated
* libray.spice modified to handle decap_12 cell
* Ali Oudhriri, Mazher Iqbal and Roselyne Chotin, April 2024
* MML April 17, 2024
**

*.include /users/cao/aoudrhiri/coriolis-2.x/src/alliance-check-toolkit/benchs/RISC-V/picorv32/skyWater130/timing/sta/skylibm/library.spice

.subckt picorv32_m VGND VPWR clk eoi[0] eoi[15] eoi[1] eoi[2] eoi[3] eoi[4] eoi[5] irq[0]
+ irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[16] irq[17] irq[18] irq[19]
+ irq[1] irq[20] irq[21] irq[22] irq[23] irq[24] irq[25] irq[26] irq[27] irq[28] irq[29]
+ irq[2] irq[30] irq[31] irq[3] irq[4] irq[5] irq[6] irq[7] irq[8] irq[9] mem_addr[10]
+ mem_addr[11] mem_addr[12] mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[16] mem_addr[17]
+ mem_addr[18] mem_addr[19] mem_addr[20] mem_addr[21] mem_addr[22] mem_addr[23] mem_addr[24]
+ mem_addr[25] mem_addr[26] mem_addr[27] mem_addr[28] mem_addr[29] mem_addr[2] mem_addr[30]
+ mem_addr[31] mem_addr[3] mem_addr[4] mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8]
+ mem_addr[9] mem_instr mem_la_addr[0] mem_la_addr[10] mem_la_addr[11] mem_la_addr[12]
+ mem_la_addr[13] mem_la_addr[14] mem_la_addr[15] mem_la_addr[16] mem_la_addr[17]
+ mem_la_addr[18] mem_la_addr[19] mem_la_addr[1] mem_la_addr[20] mem_la_addr[21] mem_la_addr[22]
+ mem_la_addr[23] mem_la_addr[24] mem_la_addr[25] mem_la_addr[26] mem_la_addr[27]
+ mem_la_addr[28] mem_la_addr[29] mem_la_addr[2] mem_la_addr[30] mem_la_addr[31] mem_la_addr[3]
+ mem_la_addr[4] mem_la_addr[5] mem_la_addr[6] mem_la_addr[7] mem_la_addr[8] mem_la_addr[9]
+ mem_la_read mem_la_wdata[0] mem_la_wdata[10] mem_la_wdata[11] mem_la_wdata[12] mem_la_wdata[13]
+ mem_la_wdata[14] mem_la_wdata[15] mem_la_wdata[16] mem_la_wdata[17] mem_la_wdata[18]
+ mem_la_wdata[19] mem_la_wdata[1] mem_la_wdata[20] mem_la_wdata[21] mem_la_wdata[22]
+ mem_la_wdata[23] mem_la_wdata[24] mem_la_wdata[25] mem_la_wdata[26] mem_la_wdata[27]
+ mem_la_wdata[28] mem_la_wdata[29] mem_la_wdata[2] mem_la_wdata[30] mem_la_wdata[31]
+ mem_la_wdata[3] mem_la_wdata[4] mem_la_wdata[5] mem_la_wdata[6] mem_la_wdata[7]
+ mem_la_wdata[8] mem_la_wdata[9] mem_la_write mem_la_wstrb[0] mem_la_wstrb[1] mem_la_wstrb[2]
+ mem_la_wstrb[3] mem_rdata[0] mem_rdata[10] mem_rdata[11] mem_rdata[12] mem_rdata[13]
+ mem_rdata[14] mem_rdata[15] mem_rdata[16] mem_rdata[17] mem_rdata[18] mem_rdata[19]
+ mem_rdata[1] mem_rdata[20] mem_rdata[21] mem_rdata[22] mem_rdata[23] mem_rdata[24]
+ mem_rdata[25] mem_rdata[26] mem_rdata[27] mem_rdata[28] mem_rdata[29] mem_rdata[2]
+ mem_rdata[30] mem_rdata[31] mem_rdata[3] mem_rdata[4] mem_rdata[5] mem_rdata[6]
+ mem_rdata[7] mem_rdata[8] mem_rdata[9] mem_ready mem_valid mem_wdata[0] mem_wdata[10]
+ mem_wdata[11] mem_wdata[12] mem_wdata[13] mem_wdata[14] mem_wdata[15] mem_wdata[16]
+ mem_wdata[17] mem_wdata[18] mem_wdata[19] mem_wdata[1] mem_wdata[20] mem_wdata[21]
+ mem_wdata[22] mem_wdata[23] mem_wdata[24] mem_wdata[25] mem_wdata[26] mem_wdata[27]
+ mem_wdata[28] mem_wdata[29] mem_wdata[2] mem_wdata[30] mem_wdata[31] mem_wdata[3]
+ mem_wdata[4] mem_wdata[5] mem_wdata[6] mem_wdata[7] mem_wdata[8] mem_wdata[9] mem_wstrb[0]
+ mem_wstrb[1] mem_wstrb[2] mem_wstrb[3] pcpi_insn[0] pcpi_insn[10] pcpi_insn[11]
+ pcpi_insn[12] pcpi_insn[13] pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17]
+ pcpi_insn[18] pcpi_insn[19] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[28]
+ pcpi_insn[29] pcpi_insn[30] pcpi_insn[31] pcpi_insn[9] pcpi_rd[0] pcpi_rd[10] pcpi_rd[11]
+ pcpi_rd[12] pcpi_rd[13] pcpi_rd[14] pcpi_rd[15] pcpi_rd[16] pcpi_rd[17] pcpi_rd[18]
+ pcpi_rd[19] pcpi_rd[1] pcpi_rd[20] pcpi_rd[21] pcpi_rd[22] pcpi_rd[23] pcpi_rd[24]
+ pcpi_rd[25] pcpi_rd[26] pcpi_rd[27] pcpi_rd[28] pcpi_rd[29] pcpi_rd[2] pcpi_rd[30]
+ pcpi_rd[31] pcpi_rd[3] pcpi_rd[4] pcpi_rd[5] pcpi_rd[6] pcpi_rd[7] pcpi_rd[8] pcpi_rd[9]
+ pcpi_ready pcpi_rs1[0] pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14]
+ pcpi_rs1[15] pcpi_rs1[16] pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20]
+ pcpi_rs1[21] pcpi_rs1[22] pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27]
+ pcpi_rs1[28] pcpi_rs1[29] pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4]
+ pcpi_rs1[5] pcpi_rs1[6] pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10]
+ pcpi_rs2[11] pcpi_rs2[12] pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17]
+ pcpi_rs2[18] pcpi_rs2[19] pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23]
+ pcpi_rs2[24] pcpi_rs2[25] pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2]
+ pcpi_rs2[30] pcpi_rs2[31] pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7]
+ pcpi_rs2[8] pcpi_rs2[9] pcpi_wait pcpi_wr resetn trace_data[0] trace_data[15] trace_data[16]
+ trace_data[1] trace_data[20] trace_data[21] trace_data[22] trace_data[23] trace_data[24]
+ trace_data[25] trace_data[26] trace_data[27] trace_data[28] trace_data[29] trace_data[2]
+ trace_data[35] trace_data[3] trace_data[4] trace_data[5] trace_data[6] trace_data[7]
+ trace_data[8] trace_data[9] trace_valid trap pcpi_insn[27] pcpi_insn[26] trace_data[14]
+ pcpi_insn[25] trace_data[13] pcpi_insn[24] trace_data[12] trace_data[34] pcpi_insn[23]
+ trace_data[33] trace_data[11] trace_data[32] trace_data[10] pcpi_valid trace_data[31]
+ trace_data[30] trace_data[19] trace_data[18] trace_data[17] eoi[14] eoi[25] eoi[24]
+ eoi[13] eoi[23] eoi[12] mem_addr[1] pcpi_insn[8] eoi[11] eoi[22] pcpi_insn[7] mem_addr[0]
+ eoi[21] eoi[10] pcpi_insn[6] eoi[31] eoi[9] eoi[20] pcpi_insn[5] eoi[30] eoi[19]
+ eoi[8] eoi[18] eoi[29] pcpi_insn[4] eoi[7] eoi[28] eoi[17] pcpi_insn[3] eoi[6] eoi[27]
+ pcpi_insn[2] eoi[16] pcpi_insn[1] eoi[26]
X_09671_ cpuregs\[20\]\[19\] cpuregs\[21\]\[19\] cpuregs\[22\]\[19\] cpuregs\[23\]\[19\]
+ _03548_ _03449_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__mux4_1
X_08622_ _03113_ _03138_ _03139_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08553_ reg_sh\[3\] reg_sh\[2\] reg_sh\[4\] VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__nor3_1
X_07504_ _02142_ _02143_ _01954_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__o21a_1
X_08484_ net252 _03015_ _01816_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_159_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07435_ _02062_ _02040_ _02077_ _02078_ _02059_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__o311a_1
XFILLER_0_119_235 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07366_ instr_rdcycleh VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_44_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_203 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09105_ cpuregs\[4\]\[3\] cpuregs\[5\]\[3\] cpuregs\[6\]\[3\] cpuregs\[7\]\[3\] _03439_
+ _03576_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__mux4_1
XFILLER_0_134_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07297_ instr_rdinstr VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_150_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_761 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_603 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09036_ _03410_ _03509_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold340 cpuregs\[30\]\[7\] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold351 cpuregs\[20\]\[19\] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold362 cpuregs\[14\]\[22\] VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 cpuregs\[12\]\[30\] VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 cpuregs\[29\]\[24\] VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 cpuregs\[9\]\[15\] VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__dlygate4sd3_1
X_09938_ _04305_ _04337_ _04339_ _02331_ decoded_imm\[26\] VGND VGND VPWR VPWR _04386_
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_148_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09869_ cpuregs\[16\]\[25\] cpuregs\[17\]\[25\] cpuregs\[18\]\[25\] cpuregs\[19\]\[25\]
+ _03548_ _03549_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__mux4_1
Xhold1040 count_cycle\[53\] VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 count_cycle\[28\] VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ _05712_ _05710_ _05714_ _05052_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__a211oi_1
X_12880_ _05041_ _06566_ _06569_ _06529_ net441 VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
*XANTENNA_202 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_213 _03401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11831_ count_cycle\[32\] count_cycle\[33\] count_cycle\[31\] _05661_ VGND VGND VPWR
+ VPWR _05667_ sky130_fd_sc_hd__and4_1
*XANTENNA_224 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_235 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ clknet_leaf_8_clk _00208_ VGND VGND VPWR VPWR cpuregs\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11762_ _05619_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_64_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13501_ _06887_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__buf_4
X_10713_ cpuregs\[26\]\[16\] _04852_ _04840_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14481_ clknet_leaf_35_clk _00139_ VGND VGND VPWR VPWR cpuregs\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11693_ _05560_ _05561_ _05564_ _05565_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13432_ _06873_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__clkbuf_1
X_10644_ _04808_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10575_ net1019 _03334_ _04768_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__mux2_1
X_13363_ net1224 _04858_ _06827_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer7 net387 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15102_ clknet_leaf_104_clk _07126_ VGND VGND VPWR VPWR reg_out\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12314_ _06026_ _06071_ _03081_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__o21a_1
X_16082_ net124 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_2
X_13294_ _06800_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__clkbuf_1
X_15033_ clknet_leaf_122_clk _00691_ VGND VGND VPWR VPWR count_cycle\[16\] sky130_fd_sc_hd__dfxtp_1
X_12245_ cpuregs\[24\]\[9\] cpuregs\[25\]\[9\] cpuregs\[26\]\[9\] cpuregs\[27\]\[9\]
+ _03095_ _05932_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__mux4_1
X_12176_ cpuregs\[0\]\[7\] cpuregs\[1\]\[7\] cpuregs\[2\]\[7\] cpuregs\[3\]\[7\] _05908_
+ _05909_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__mux4_1
X_11127_ net559 _05095_ _05097_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__o21a_1
X_11058_ _05048_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__clkbuf_1
X_15935_ clknet_leaf_132_clk _01507_ VGND VGND VPWR VPWR cpuregs\[0\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10009_ decoded_imm\[30\] _02380_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__or2_1
X_15866_ clknet_leaf_135_clk _01438_ VGND VGND VPWR VPWR cpuregs\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_14817_ clknet_leaf_147_clk _00475_ VGND VGND VPWR VPWR cpuregs\[25\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15797_ clknet_leaf_141_clk _01372_ VGND VGND VPWR VPWR cpuregs\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14748_ clknet_leaf_157_clk _00406_ VGND VGND VPWR VPWR cpuregs\[26\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14679_ clknet_leaf_152_clk _00337_ VGND VGND VPWR VPWR cpuregs\[27\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07220_ _01882_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07151_ _01819_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_1
XFILLER_0_27_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_497 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07984_ _02507_ _02503_ _02509_ _02573_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09723_ decoded_imm\[21\] net184 VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__nand2_1
X_09654_ _03574_ _04102_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08605_ _03054_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_143_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09585_ _03500_ _04043_ _03468_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_49_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08536_ _03035_ _03041_ _03044_ _03049_ _03055_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_46_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08467_ _03004_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_1
XFILLER_0_93_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07418_ _02062_ _02040_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08398_ _02956_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_1
XFILLER_0_46_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07349_ _01996_ _01997_ _01954_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__o21a_2
XFILLER_0_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_912 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10360_ cpuregs\[28\]\[19\] _03307_ _04647_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09019_ _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__inv_2
X_10291_ _04620_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__clkbuf_1
X_12030_ is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__inv_2
Xhold170 instr_lhu VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 cpuregs\[0\]\[28\] VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 instr_slt VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13981_ net1316 _06937_ _01602_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__mux2_1
X_15720_ clknet_leaf_31_clk _01295_ VGND VGND VPWR VPWR cpuregs\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12932_ decoded_imm_j\[10\] _01092_ _03169_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__mux2_1
X_15651_ clknet_leaf_45_clk _01226_ VGND VGND VPWR VPWR cpuregs\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12863_ net672 _06554_ _06556_ net647 VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14602_ clknet_leaf_54_clk _00260_ VGND VGND VPWR VPWR cpuregs\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11814_ net487 _05652_ _05647_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__o21ai_1
X_15582_ clknet_leaf_21_clk _01157_ VGND VGND VPWR VPWR cpuregs\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12794_ _06521_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__buf_1
XFILLER_0_157_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14533_ clknet_leaf_137_clk _00191_ VGND VGND VPWR VPWR cpuregs\[13\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11745_ net542 _05604_ _05169_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_99_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14464_ clknet_leaf_137_clk _00122_ VGND VGND VPWR VPWR cpuregs\[12\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11676_ _05494_ _05251_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_558 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13415_ net1110 _04842_ _06863_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__mux2_1
X_10627_ _04799_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__clkbuf_1
X_14395_ clknet_leaf_135_clk _00058_ VGND VGND VPWR VPWR cpuregs\[11\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13346_ _06828_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_720 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_306 VGND VGND VPWR VPWR picorv32_306/HI pcpi_insn[16] sky130_fd_sc_hd__conb_1
X_10558_ net1103 _03282_ _04757_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__mux2_1
Xpicorv32_317 VGND VGND VPWR VPWR picorv32_317/HI pcpi_insn[27] sky130_fd_sc_hd__conb_1
Xpicorv32_328 VGND VGND VPWR VPWR picorv32_328/HI trace_data[5] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_339 VGND VGND VPWR VPWR picorv32_339/HI trace_data[16] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_94_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13277_ net1175 _04839_ _06791_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10489_ cpuregs\[14\]\[15\] _03282_ _04720_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15016_ clknet_leaf_106_clk _00674_ VGND VGND VPWR VPWR reg_next_pc\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12228_ _02476_ _05989_ _05863_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12159_ cpuregs\[20\]\[6\] cpuregs\[21\]\[6\] cpuregs\[22\]\[6\] cpuregs\[23\]\[6\]
+ _05921_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_35 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_87_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15918_ clknet_leaf_5_clk _01490_ VGND VGND VPWR VPWR cpuregs\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_160_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15849_ clknet_leaf_34_clk _01421_ VGND VGND VPWR VPWR cpuregs\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_125_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09370_ _03795_ _03831_ _03834_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08321_ _02380_ _02909_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_96_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08252_ _02845_ _02846_ _02844_ _02807_ _02847_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_694 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_222 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07203_ instr_lhu instr_lh _01867_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_41_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08183_ net180 _02783_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_160_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput220 net220 VGND VGND VPWR VPWR pcpi_rs2[25] sky130_fd_sc_hd__buf_2
Xoutput231 net231 VGND VGND VPWR VPWR pcpi_rs2[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_145_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07967_ _02584_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__clkbuf_4
X_09706_ cpuregs\[24\]\[20\] cpuregs\[25\]\[20\] cpuregs\[26\]\[20\] cpuregs\[27\]\[20\]
+ _03640_ _03496_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__mux4_1
X_07898_ net249 VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09637_ _03075_ _04091_ _04093_ _01943_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__o211a_1
X_09568_ _04025_ _04026_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08519_ _00008_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__buf_4
X_09499_ _03890_ _03959_ _03075_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11530_ _05193_ reg_next_pc\[14\] _05220_ _05403_ _01905_ VGND VGND VPWR VPWR _05417_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_182 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11461_ _05346_ _05349_ _05351_ _05345_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_156_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13200_ decoded_imm\[24\] _06740_ _06737_ _06748_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__o22a_1
X_10412_ _04685_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__clkbuf_1
X_11392_ _05288_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__clkbuf_4
X_14180_ _01714_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13131_ net148 net110 _06707_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__mux2_1
X_10343_ _04648_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_775 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_131_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10274_ net1395 _03248_ _04611_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__mux2_1
X_13062_ net1082 _04881_ _06635_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__mux2_1
X_12013_ _05793_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13964_ _01599_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__clkbuf_1
X_15703_ clknet_leaf_134_clk _01278_ VGND VGND VPWR VPWR cpuregs\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12915_ _06592_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__clkbuf_1
X_13895_ _01562_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__clkbuf_1
X_15634_ clknet_leaf_155_clk _01209_ VGND VGND VPWR VPWR cpuregs\[23\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12846_ net956 _06554_ _06556_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15565_ clknet_leaf_17_clk _01140_ VGND VGND VPWR VPWR cpuregs\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ instr_lb _01928_ _06509_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_131_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ clknet_leaf_10_clk _00174_ VGND VGND VPWR VPWR cpuregs\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11728_ _05052_ net431 VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_618 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15496_ clknet_leaf_89_clk _01081_ VGND VGND VPWR VPWR mem_rdata_q\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_126_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14447_ clknet_leaf_38_clk _00105_ VGND VGND VPWR VPWR cpuregs\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11659_ _05530_ _05532_ _05533_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__nor3_1
XFILLER_0_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_107_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14378_ clknet_leaf_26_clk _00041_ VGND VGND VPWR VPWR cpuregs\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold906 cpuregs\[13\]\[23\] VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold917 cpuregs\[15\]\[31\] VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ _06819_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__clkbuf_1
Xhold928 cpuregs\[12\]\[0\] VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 cpuregs\[16\]\[25\] VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_110_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08870_ reg_pc\[26\] _03345_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07821_ net192 net224 VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07752_ count_instr\[30\] _02054_ count_cycle\[30\] _02020_ _02373_ VGND VGND VPWR
+ VPWR _02374_ sky130_fd_sc_hd__a221o_2
X_07683_ reg_pc\[25\] decoded_imm\[25\] VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_140_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09422_ _03474_ _03876_ _03885_ _03527_ reg_pc\[11\] VGND VGND VPWR VPWR _03886_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_149_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09353_ cpuregs\[24\]\[9\] cpuregs\[25\]\[9\] cpuregs\[26\]\[9\] cpuregs\[27\]\[9\]
+ _03438_ _03812_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08304_ _02568_ _02618_ _02439_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_916 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09284_ cpuregs\[20\]\[7\] cpuregs\[21\]\[7\] cpuregs\[22\]\[7\] cpuregs\[23\]\[7\]
+ _03598_ _03460_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08235_ _02801_ _02808_ _02818_ _02832_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__o31a_1
XFILLER_0_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_826 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08166_ net247 _02759_ _02656_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08097_ net174 _02703_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08999_ _03473_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10961_ _04991_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__clkbuf_1
X_12700_ cpuregs\[12\]\[29\] cpuregs\[13\]\[29\] cpuregs\[14\]\[29\] cpuregs\[15\]\[29\]
+ _03133_ _03134_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__mux4_1
X_13680_ cpuregs\[23\]\[25\] _06977_ _07014_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__mux2_1
X_10892_ net860 _04879_ _04945_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12631_ _03042_ _06374_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15350_ clknet_leaf_68_clk _00940_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12562_ _06309_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14301_ net577 VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__clkbuf_1
X_11513_ _05394_ _05399_ _05393_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__o21ai_2
X_15281_ clknet_leaf_105_clk _00874_ VGND VGND VPWR VPWR decoded_imm_j\[18\] sky130_fd_sc_hd__dfxtp_1
X_12493_ net213 _06243_ _06052_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14232_ _01741_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__clkbuf_1
X_11444_ _05322_ _05331_ _05335_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14163_ net906 _06983_ _01696_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11375_ _05269_ _05271_ _05272_ _05191_ _05273_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__a32o_1
XFILLER_0_150_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13114_ net139 net101 _06696_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__mux2_1
X_10326_ _04639_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__clkbuf_1
X_14094_ _01668_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__clkbuf_1
X_13045_ _06660_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__clkbuf_1
X_10257_ cpuregs\[2\]\[2\] _03194_ _04600_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__mux2_1
X_10188_ _04566_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__clkbuf_1
X_14996_ clknet_leaf_86_clk _00654_ VGND VGND VPWR VPWR reg_next_pc\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13947_ net1236 _06971_ _01588_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13878_ net1079 _06971_ _01551_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15617_ clknet_leaf_28_clk _01192_ VGND VGND VPWR VPWR cpuregs\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12829_ _06546_ _06542_ _06547_ _06530_ net455 VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__a32o_1
XFILLER_0_158_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15548_ clknet_leaf_81_clk _00021_ VGND VGND VPWR VPWR cpu_state\[4\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_150_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_501 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15479_ clknet_leaf_83_clk _01064_ VGND VGND VPWR VPWR mem_rdata_q\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_651 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08020_ net199 _02632_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold703 cpuregs\[13\]\[25\] VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold714 cpuregs\[25\]\[11\] VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold725 cpuregs\[8\]\[15\] VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_40_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold736 cpuregs\[26\]\[6\] VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 cpuregs\[28\]\[9\] VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 cpuregs\[12\]\[10\] VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _03403_ _04417_ _03420_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__o21a_1
Xhold769 cpuregs\[25\]\[4\] VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__dlygate4sd3_1
X_08922_ _01854_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__clkbuf_4
X_08853_ reg_out\[24\] alu_out_q\[24\] _03176_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07804_ _02290_ net218 VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__or2b_1
X_08784_ _03276_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_28_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ _01943_ net253 _02184_ _02358_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__a22o_1
X_07666_ count_instr\[24\] _01965_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09405_ cpuregs\[4\]\[11\] cpuregs\[5\]\[11\] cpuregs\[6\]\[11\] cpuregs\[7\]\[11\]
+ _03405_ _03409_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07597_ count_instr\[19\] _02054_ count_cycle\[51\] _02055_ VGND VGND VPWR VPWR _02230_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09336_ cpuregs\[4\]\[9\] cpuregs\[5\]\[9\] cpuregs\[6\]\[9\] cpuregs\[7\]\[9\] _03800_
+ _03801_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_510 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_118_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09267_ decoded_imm\[7\] net200 VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_141_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_141_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_62_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08218_ net184 _02815_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_153_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09198_ _03075_ _03667_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08149_ _02706_ _02720_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_56_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11160_ count_instr\[34\] net376 count_instr\[35\] VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__a21o_1
X_10111_ latched_rd\[0\] _01877_ _03181_ latched_rd\[1\] VGND VGND VPWR VPWR _04523_
+ sky130_fd_sc_hd__or4b_1
X_11091_ _05070_ _05068_ _05072_ _05052_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__a211oi_1
X_10042_ _04481_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__nor2_2
X_14850_ clknet_leaf_128_clk _00508_ VGND VGND VPWR VPWR cpuregs\[20\]\[24\] sky130_fd_sc_hd__dfxtp_1
Xhold52 mem_rdata[30] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold63 mem_rdata[10] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 decoded_rd\[1\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 instr_fence VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ net1307 _06962_ _07075_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__mux2_1
Xhold96 instr_bltu VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ clknet_leaf_157_clk _00439_ VGND VGND VPWR VPWR cpuregs\[16\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11993_ net41 net72 _05774_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13732_ _07047_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__clkbuf_1
X_10944_ net788 _04863_ _04981_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13663_ net1238 _06960_ _07003_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10875_ _04946_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15402_ clknet_leaf_85_clk _00992_ VGND VGND VPWR VPWR decoded_imm\[6\] sky130_fd_sc_hd__dfxtp_2
X_12614_ _03132_ _06358_ _05840_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__o21a_1
XFILLER_0_155_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13594_ cpuregs\[31\]\[21\] _06969_ _06967_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15333_ clknet_leaf_75_clk _00923_ VGND VGND VPWR VPWR mem_state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12545_ _05845_ _06290_ _06292_ _03139_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_132_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_132_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15264_ clknet_leaf_85_clk _00857_ VGND VGND VPWR VPWR decoded_imm_j\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12476_ cpuregs\[0\]\[19\] cpuregs\[1\]\[19\] cpuregs\[2\]\[19\] cpuregs\[3\]\[19\]
+ _06055_ _05829_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14215_ net1220 _06966_ _01732_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_5 _01872_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11427_ decoded_imm_j\[7\] _05204_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15195_ clknet_leaf_70_clk alu_out\[8\] VGND VGND VPWR VPWR alu_out_q\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14146_ _01673_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11358_ _01872_ _05259_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10309_ net1359 _03360_ _04622_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__mux2_1
X_14077_ _01659_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__clkbuf_1
X_11289_ _05188_ reg_pc\[10\] VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__or2_1
X_13028_ _06651_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer17 _05116_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer28 net388 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_1
Xrebuffer39 net399 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_1
X_14979_ clknet_leaf_103_clk _00637_ VGND VGND VPWR VPWR reg_pc\[25\] sky130_fd_sc_hd__dfxtp_2
X_07520_ _02019_ _02148_ _02158_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07451_ reg_pc\[9\] decoded_imm\[9\] VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07382_ _02023_ _02027_ _02026_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_510 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09121_ _03446_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_123_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_123_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_576 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09052_ _03525_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_135_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08003_ _02618_ _02568_ _02499_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__mux2_1
Xhold500 cpuregs\[9\]\[13\] VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 cpuregs\[6\]\[28\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold522 cpuregs\[20\]\[31\] VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold533 cpuregs\[15\]\[6\] VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 cpuregs\[29\]\[28\] VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 cpuregs\[13\]\[12\] VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 cpuregs\[17\]\[27\] VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 cpuregs\[25\]\[30\] VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold588 cpuregs\[19\]\[30\] VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ decoded_imm\[28\] net253 VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__nand2_1
Xhold599 cpuregs\[25\]\[21\] VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ net1324 _03381_ _03184_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _02380_ _03619_ _04264_ _03657_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__a211o_1
X_08836_ _03321_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__clkbuf_4
X_08767_ _03257_ _03260_ _03261_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__mux2_4
X_07718_ _01970_ _02339_ _02342_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__a21oi_1
X_08698_ _03201_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_49_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ _01977_ _02277_ _02201_ _02278_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_203 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10660_ _04816_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09319_ cpuregs\[24\]\[8\] cpuregs\[25\]\[8\] cpuregs\[26\]\[8\] cpuregs\[27\]\[8\]
+ _03494_ _03497_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_114_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_114_clk sky130_fd_sc_hd__clkbuf_2
X_10591_ net867 _03386_ _04745_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12330_ cpuregs\[8\]\[13\] cpuregs\[9\]\[13\] cpuregs\[10\]\[13\] cpuregs\[11\]\[13\]
+ _05907_ _03047_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12261_ cpuregs\[20\]\[10\] cpuregs\[21\]\[10\] cpuregs\[22\]\[10\] cpuregs\[23\]\[10\]
+ _05921_ _05922_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__mux4_1
X_14000_ net1304 _06956_ _01613_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__mux2_1
X_11212_ net525 _05155_ _05133_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__o21ai_1
X_12192_ _05947_ _05950_ _05952_ _05954_ _03080_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput42 net42 VGND VGND VPWR VPWR mem_addr[17] sky130_fd_sc_hd__clkbuf_4
X_11143_ _05107_ _05108_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__nor2_1
Xoutput53 net53 VGND VGND VPWR VPWR mem_addr[28] sky130_fd_sc_hd__buf_2
Xoutput64 net64 VGND VGND VPWR VPWR mem_addr[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput75 net75 VGND VGND VPWR VPWR mem_la_addr[19] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 VGND VGND VPWR VPWR mem_la_addr[2] sky130_fd_sc_hd__clkbuf_4
Xoutput97 net97 VGND VGND VPWR VPWR mem_la_wdata[0] sky130_fd_sc_hd__clkbuf_4
X_11074_ net456 VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__inv_2
X_15951_ clknet_leaf_13_clk _01523_ VGND VGND VPWR VPWR cpuregs\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_14902_ clknet_leaf_102_clk _00560_ VGND VGND VPWR VPWR count_instr\[11\] sky130_fd_sc_hd__dfxtp_1
X_10025_ cpuregs\[12\]\[30\] cpuregs\[13\]\[30\] cpuregs\[14\]\[30\] cpuregs\[15\]\[30\]
+ _03680_ _03443_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__mux4_1
X_15882_ clknet_leaf_57_clk _01454_ VGND VGND VPWR VPWR cpuregs\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14833_ clknet_leaf_36_clk _00491_ VGND VGND VPWR VPWR cpuregs\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14764_ clknet_leaf_28_clk _00422_ VGND VGND VPWR VPWR cpuregs\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11976_ _05766_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13715_ _07038_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__clkbuf_1
X_10927_ cpuregs\[20\]\[13\] _04846_ _04970_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__mux2_1
X_14695_ clknet_leaf_127_clk _00353_ VGND VGND VPWR VPWR cpuregs\[27\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13646_ net1127 _06943_ _06992_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__mux2_1
X_10858_ _04937_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_567 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13577_ _03286_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_105_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_105_clk sky130_fd_sc_hd__clkbuf_2
X_10789_ net1380 _04844_ _04898_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15316_ clknet_leaf_145_clk _00906_ VGND VGND VPWR VPWR cpuregs\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12528_ _06026_ _06276_ _06193_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_117_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15247_ clknet_leaf_77_clk _00840_ VGND VGND VPWR VPWR instr_sll sky130_fd_sc_hd__dfxtp_1
X_12459_ cpuregs\[24\]\[18\] cpuregs\[25\]\[18\] cpuregs\[26\]\[18\] cpuregs\[27\]\[18\]
+ _05970_ _03108_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15178_ clknet_leaf_98_clk _00803_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_130_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14129_ _01687_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09670_ _03547_ _04121_ _04123_ _04125_ _03489_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08621_ _00010_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__buf_4
XFILLER_0_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08552_ _03071_ decoded_imm_j\[2\] is_slli_srli_srai VGND VGND VPWR VPWR _03072_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07503_ count_instr\[12\] instr_rdinstr count_cycle\[12\] _01950_ VGND VGND VPWR
+ VPWR _02143_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08483_ reg_next_pc\[31\] reg_out\[31\] _02991_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_605 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_76_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07434_ _02075_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_478 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07365_ _01946_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_44_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09104_ _03549_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07296_ count_instr\[32\] _01946_ _01947_ count_cycle\[32\] VGND VGND VPWR VPWR _01948_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09035_ cpuregs\[4\]\[1\] cpuregs\[5\]\[1\] _03494_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold330 decoded_imm\[3\] VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 cpuregs\[0\]\[19\] VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold352 cpuregs\[1\]\[26\] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 cpuregs\[18\]\[4\] VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold374 mem_do_rdata VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 cpuregs\[4\]\[24\] VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 cpuregs\[19\]\[26\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09937_ decoded_imm\[27\] net190 VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _03807_ _04317_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__or2_1
Xhold1030 cpuregs\[8\]\[3\] VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 count_instr\[44\] VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 count_instr\[21\] VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__clkbuf_4
X_09799_ _03647_ _04250_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__or2_1
*XANTENNA_203 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11830_ _05666_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__clkbuf_1
*XANTENNA_214 _03401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_225 _03108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_236 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _05617_ _05113_ _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_37_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _06909_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__clkbuf_1
X_10712_ _03286_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14480_ clknet_leaf_33_clk _00138_ VGND VGND VPWR VPWR cpuregs\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11692_ _05549_ _05562_ _05563_ _05288_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__o31a_1
X_13431_ net1228 _04858_ _06863_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__mux2_1
X_10643_ net1364 _03334_ _04804_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13362_ _06836_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__clkbuf_1
X_10574_ _04771_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer8 _05667_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_1
X_15101_ clknet_leaf_100_clk _07124_ VGND VGND VPWR VPWR reg_out\[19\] sky130_fd_sc_hd__dfxtp_1
X_12313_ cpuregs\[28\]\[12\] cpuregs\[29\]\[12\] cpuregs\[30\]\[12\] cpuregs\[31\]\[12\]
+ _05895_ _05929_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16081_ net123 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_2
X_13293_ net1130 _04856_ _06791_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_125_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_760 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15032_ clknet_leaf_132_clk _00690_ VGND VGND VPWR VPWR count_cycle\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_911 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12244_ _03083_ _06004_ _03081_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ cpuregs\[4\]\[7\] cpuregs\[5\]\[7\] cpuregs\[6\]\[7\] cpuregs\[7\]\[7\] _05834_
+ _03097_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__mux4_1
X_11126_ net1414 _05095_ _05052_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__a21oi_1
X_15934_ clknet_leaf_134_clk _01506_ VGND VGND VPWR VPWR cpuregs\[0\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11057_ _01905_ _05046_ _05047_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10008_ decoded_imm\[30\] _02380_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_134_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15865_ clknet_leaf_140_clk _01437_ VGND VGND VPWR VPWR cpuregs\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_14816_ clknet_leaf_149_clk _00474_ VGND VGND VPWR VPWR cpuregs\[25\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15796_ clknet_leaf_102_clk _01371_ VGND VGND VPWR VPWR cpuregs\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14747_ clknet_leaf_160_clk _00405_ VGND VGND VPWR VPWR cpuregs\[26\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_512 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11959_ _05762_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__buf_2
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14678_ clknet_leaf_155_clk _00336_ VGND VGND VPWR VPWR cpuregs\[27\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_690 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_129_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13629_ _06993_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07150_ net34 _01818_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07983_ _02514_ _02581_ _02599_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__a21o_1
X_09722_ _02250_ _03624_ _04176_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09653_ _04104_ _04106_ _04109_ _03433_ _03591_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a221o_1
X_08604_ reg_sh\[3\] reg_sh\[2\] reg_sh\[4\] VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__o21a_1
X_09584_ cpuregs\[8\]\[16\] cpuregs\[9\]\[16\] cpuregs\[10\]\[16\] cpuregs\[11\]\[16\]
+ _03680_ _03461_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_143_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08535_ _03050_ _03053_ _03054_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08466_ _02316_ _03003_ _02993_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07417_ reg_pc\[6\] decoded_imm\[6\] VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08397_ _02008_ _02955_ _02951_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_811 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07348_ count_instr\[3\] instr_rdinstr count_cycle\[3\] _01950_ VGND VGND VPWR VPWR
+ _01997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07279_ mem_wordsize\[2\] mem_wordsize\[1\] VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__nor2_4
XFILLER_0_5_481 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09018_ _03408_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__buf_6
X_10290_ cpuregs\[2\]\[18\] _03302_ _04611_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold160 net44 VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 cpuregs\[0\]\[24\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 mem_rdata_q\[19\] VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 cpuregs\[0\]\[23\] VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
X_13980_ _01608_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__clkbuf_1
X_12931_ _06600_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__clkbuf_1
X_15650_ clknet_leaf_37_clk _01225_ VGND VGND VPWR VPWR cpuregs\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12862_ _06546_ _06548_ _06559_ _06562_ net453 VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11813_ count_cycle\[25\] count_cycle\[26\] count_cycle\[27\] _05649_ VGND VGND VPWR
+ VPWR _05655_ sky130_fd_sc_hd__and4_4
X_14601_ clknet_leaf_20_clk _00259_ VGND VGND VPWR VPWR cpuregs\[28\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15581_ clknet_leaf_22_clk _01156_ VGND VGND VPWR VPWR cpuregs\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12793_ mem_rdata_q\[4\] net27 _03017_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__mux2_1
X_14532_ clknet_leaf_137_clk _00190_ VGND VGND VPWR VPWR cpuregs\[13\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11744_ count_cycle\[4\] count_cycle\[5\] count_cycle\[6\] _05601_ VGND VGND VPWR
+ VPWR _05607_ sky130_fd_sc_hd__and4_1
XFILLER_0_154_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14463_ clknet_leaf_97_clk _00121_ VGND VGND VPWR VPWR cpuregs\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11675_ _05494_ _05251_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__and2_1
X_13414_ _06864_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10626_ cpuregs\[15\]\[15\] _03282_ _04793_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__mux2_1
X_14394_ clknet_leaf_139_clk _00057_ VGND VGND VPWR VPWR cpuregs\[11\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13345_ cpuregs\[19\]\[10\] _04839_ _06827_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_106_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10557_ _04762_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpicorv32_307 VGND VGND VPWR VPWR picorv32_307/HI pcpi_insn[17] sky130_fd_sc_hd__conb_1
Xpicorv32_318 VGND VGND VPWR VPWR picorv32_318/HI pcpi_insn[28] sky130_fd_sc_hd__conb_1
XFILLER_0_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_329 VGND VGND VPWR VPWR picorv32_329/HI trace_data[6] sky130_fd_sc_hd__conb_1
X_13276_ _06779_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_94_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10488_ _04725_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_94_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15015_ clknet_leaf_108_clk _00673_ VGND VGND VPWR VPWR reg_next_pc\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_110_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_264 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12227_ _05901_ _05968_ _05988_ _05904_ decoded_imm\[8\] VGND VGND VPWR VPWR _05989_
+ sky130_fd_sc_hd__a32o_1
X_12158_ _03052_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__clkbuf_8
X_11109_ net478 count_instr\[18\] _05082_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_142_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12089_ _03124_ _05857_ _03054_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__o21ai_1
X_15917_ clknet_leaf_7_clk _01489_ VGND VGND VPWR VPWR cpuregs\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_160_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ clknet_leaf_34_clk _01420_ VGND VGND VPWR VPWR cpuregs\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_125_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_903 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15779_ clknet_leaf_47_clk _01354_ VGND VGND VPWR VPWR cpuregs\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08320_ _02380_ _02909_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_515 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08251_ _02831_ _02832_ _02838_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_151_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07202_ instr_lbu instr_lw instr_lb VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_234 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08182_ net180 _02783_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_41_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput210 net210 VGND VGND VPWR VPWR pcpi_rs2[16] sky130_fd_sc_hd__buf_2
Xoutput221 net221 VGND VGND VPWR VPWR pcpi_rs2[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput232 net232 VGND VGND VPWR VPWR pcpi_rs2[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_160_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07966_ net240 VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__clkbuf_4
X_09705_ _04158_ _04159_ _03413_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07897_ _01992_ _02502_ _02516_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_94_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_2
X_09636_ _02237_ _03481_ _04092_ _03616_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09567_ _04022_ _04023_ _04024_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_139_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08518_ _00007_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__buf_4
X_09498_ _02154_ _03619_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_19_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08449_ _02948_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11460_ _05345_ _05346_ _05349_ _05351_ _01889_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__a41o_1
XFILLER_0_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10411_ net1093 _03248_ _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11391_ instr_jal VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13130_ _06708_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10342_ net1353 _03248_ _04647_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_787 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13061_ _06668_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__clkbuf_1
X_10273_ _04599_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__clkbuf_8
X_12012_ net50 net81 _05785_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13963_ net931 _06987_ _01565_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_85_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_2
X_15702_ clknet_leaf_145_clk _01277_ VGND VGND VPWR VPWR cpuregs\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12914_ mem_rdata_q\[26\] net19 _06589_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__mux2_1
X_13894_ net1111 _06987_ _07099_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15633_ clknet_leaf_154_clk _01208_ VGND VGND VPWR VPWR cpuregs\[23\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12845_ _06553_ _06555_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15564_ clknet_leaf_18_clk _01139_ VGND VGND VPWR VPWR cpuregs\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12776_ latched_is_lh _06509_ _06510_ _05257_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_802 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11727_ _05185_ _05595_ _05596_ _05257_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__o211a_1
X_14515_ clknet_leaf_31_clk _00173_ VGND VGND VPWR VPWR cpuregs\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15495_ clknet_leaf_89_clk _01080_ VGND VGND VPWR VPWR mem_rdata_q\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11658_ _05530_ _05532_ _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__o21a_1
X_14446_ clknet_leaf_54_clk _00104_ VGND VGND VPWR VPWR cpuregs\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10609_ net1171 _03228_ _04782_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14377_ clknet_leaf_38_clk _00040_ VGND VGND VPWR VPWR cpuregs\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11589_ _05230_ _05233_ _05448_ _05235_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold907 cpuregs\[26\]\[4\] VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold918 cpuregs\[8\]\[31\] VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ net895 _04823_ _06816_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_540 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold929 cpuregs\[22\]\[13\] VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_110_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13259_ _06782_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_20_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07820_ net192 net224 VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07751_ count_instr\[62\] _01946_ _02014_ count_cycle\[62\] VGND VGND VPWR VPWR _02373_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_76_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_2
X_07682_ _02019_ _02296_ _02309_ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_140_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09421_ _03878_ _03880_ _03882_ _03884_ _03760_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__a221o_4
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09352_ _03446_ _03817_ _03418_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08303_ _02892_ _02893_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09283_ _03575_ _03745_ _03748_ _03750_ _03591_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08234_ _02799_ _02816_ _02817_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08165_ _02584_ _02765_ _02766_ _02768_ _02538_ VGND VGND VPWR VPWR alu_out\[16\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_31_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08096_ net174 _02703_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_54_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__buf_4
X_07949_ _02568_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_67_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_2
X_10960_ net1366 _04879_ _04981_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09619_ _02200_ _03660_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__and2_1
X_10891_ _04954_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__clkbuf_1
X_12630_ cpuregs\[8\]\[26\] cpuregs\[9\]\[26\] cpuregs\[10\]\[26\] cpuregs\[11\]\[26\]
+ _05907_ _03039_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12561_ net217 _06308_ _06282_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11512_ _05393_ _05394_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__or3_1
X_14300_ _01775_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__clkbuf_1
X_15280_ clknet_leaf_99_clk _00873_ VGND VGND VPWR VPWR decoded_imm_j\[17\] sky130_fd_sc_hd__dfxtp_2
X_12492_ _06132_ _06233_ _06242_ _06153_ decoded_imm\[19\] VGND VGND VPWR VPWR _06243_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14231_ net1206 _06983_ _01732_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11443_ _05322_ _05331_ _05335_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14162_ _01704_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__clkbuf_1
X_11374_ _01901_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13113_ _06699_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10325_ cpuregs\[28\]\[2\] _03194_ _04636_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14093_ cpuregs\[6\]\[27\] _06981_ _01660_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__mux2_1
X_13044_ net1360 _04863_ _06658_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__mux2_1
X_10256_ _04602_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10187_ net1242 _03189_ _04564_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14995_ clknet_leaf_86_clk _00653_ VGND VGND VPWR VPWR reg_next_pc\[10\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_58_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_89_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13946_ _01590_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_105_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13877_ _01553_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15616_ clknet_leaf_53_clk _01191_ VGND VGND VPWR VPWR cpuregs\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12828_ _06533_ mem_rdata_q\[13\] _06532_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15547_ clknet_leaf_81_clk _00020_ VGND VGND VPWR VPWR cpu_state\[3\] sky130_fd_sc_hd__dfxtp_4
X_12759_ _03106_ _06497_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15478_ clknet_leaf_82_clk _01063_ VGND VGND VPWR VPWR mem_rdata_q\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_513 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14429_ clknet_leaf_60_clk _00087_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_142_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold704 cpuregs\[1\]\[24\] VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold715 cpuregs\[14\]\[20\] VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold726 cpuregs\[6\]\[15\] VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 cpuregs\[29\]\[4\] VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_666 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_189 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09970_ cpuregs\[28\]\[28\] cpuregs\[29\]\[28\] cpuregs\[30\]\[28\] cpuregs\[31\]\[28\]
+ _03494_ _03497_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__mux4_1
Xhold748 cpuregs\[18\]\[14\] VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 cpuregs\[20\]\[15\] VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08921_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08852_ _03335_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__clkbuf_1
X_07803_ _02237_ _02409_ _02422_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__o21a_1
X_08783_ net1384 _03275_ _03249_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_49_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07734_ net21 _02251_ _02179_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__a21o_1
X_07665_ _02019_ _02284_ _02293_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09404_ _03866_ _03867_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__and2b_1
X_07596_ count_instr\[51\] _02052_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09335_ _00013_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_610 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09266_ decoded_imm\[7\] net200 VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_630 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_133_602 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_63_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08217_ net184 _02815_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_153_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09197_ _01845_ _02099_ _03619_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_646 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_31_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08148_ _02745_ _02749_ _02750_ _02751_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08079_ _02480_ _02569_ _02688_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__a21o_1
X_10110_ latched_rd\[3\] latched_rd\[4\] latched_rd\[2\] VGND VGND VPWR VPWR _04522_
+ sky130_fd_sc_hd__nand3_4
X_11090_ count_instr\[11\] count_instr\[10\] _05062_ _05071_ VGND VGND VPWR VPWR _05072_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_101_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10041_ _04484_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__buf_4
Xhold53 mem_rdata[0] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 mem_rdata[28] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 reg_sh\[0\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _07083_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__clkbuf_1
Xhold86 mem_rdata_q\[7\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 count_instr\[9\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_622 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14780_ clknet_leaf_152_clk _00438_ VGND VGND VPWR VPWR cpuregs\[16\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11992_ _05782_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13731_ net1212 _06960_ _07039_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__mux2_1
X_10943_ _04982_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_210 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13662_ _07010_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__clkbuf_1
X_10874_ net1007 _04860_ _04945_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15401_ clknet_leaf_85_clk _00991_ VGND VGND VPWR VPWR decoded_imm\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12613_ cpuregs\[16\]\[25\] cpuregs\[17\]\[25\] cpuregs\[18\]\[25\] cpuregs\[19\]\[25\]
+ _05984_ _06068_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13593_ _03321_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_574 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_155_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_93_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12544_ _03042_ _06291_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__or2_1
X_15332_ clknet_leaf_75_clk _00922_ VGND VGND VPWR VPWR mem_state\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12475_ cpuregs\[4\]\[19\] cpuregs\[5\]\[19\] cpuregs\[6\]\[19\] cpuregs\[7\]\[19\]
+ _06011_ _06156_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__mux4_1
X_15263_ clknet_leaf_85_clk _00856_ VGND VGND VPWR VPWR decoded_imm_j\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14214_ _01709_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__buf_4
X_11426_ _05258_ net533 _05239_ _05320_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_6 _01884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15194_ clknet_leaf_74_clk alu_out\[7\] VGND VGND VPWR VPWR alu_out_q\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14145_ _01695_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__clkbuf_1
X_11357_ reg_next_pc\[30\] _03378_ _02948_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10308_ _04629_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__clkbuf_1
X_14076_ cpuregs\[6\]\[19\] _06964_ _01649_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__mux2_1
X_11288_ reg_next_pc\[10\] _03243_ _02946_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13027_ net866 _04846_ _06647_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__mux2_1
X_10239_ net1077 _03355_ _04586_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__mux2_1
Xrebuffer18 _05109_ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_1
Xrebuffer29 net389 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_1
X_14978_ clknet_leaf_112_clk _00636_ VGND VGND VPWR VPWR reg_pc\[24\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_159_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13929_ _01581_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_157_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07450_ count_instr\[9\] _02054_ count_cycle\[9\] _02020_ _02092_ VGND VGND VPWR
+ VPWR _02093_ sky130_fd_sc_hd__a221o_2
XFILLER_0_9_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07381_ _02023_ _02026_ _02027_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__or3_1
XFILLER_0_123_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_714 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09120_ _03575_ _03580_ _03585_ _03590_ _03591_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__a221o_2
XFILLER_0_29_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09051_ instr_lui is_lui_auipc_jal VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__and2b_2
XFILLER_0_4_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08002_ _02560_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold501 cpuregs\[25\]\[29\] VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold512 cpuregs\[9\]\[31\] VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold523 count_instr\[28\] VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold534 cpuregs\[13\]\[6\] VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold545 cpuregs\[10\]\[13\] VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 cpuregs\[24\]\[18\] VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold567 cpuregs\[7\]\[12\] VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 cpuregs\[21\]\[9\] VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ decoded_imm\[28\] net253 VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__nor2_1
Xhold589 cpuregs\[17\]\[9\] VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08904_ _03380_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_51_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _04333_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08835_ _03317_ _03320_ _03293_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__mux2_1
X_08766_ _03199_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__clkbuf_4
X_07717_ _02007_ _02340_ _02201_ _02341_ _01955_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__a221o_1
X_08697_ _03173_ _03196_ _03197_ _03200_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_49_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ net15 _02252_ _02180_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_49_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07579_ net9 _02202_ _02179_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09318_ _03783_ _03784_ _03437_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10590_ _04779_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09249_ _03581_ _03717_ _03467_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12260_ _05879_ _06015_ _06017_ _06019_ _03104_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__a221o_2
XFILLER_0_105_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11211_ count_instr\[50\] count_instr\[47\] _05146_ _05154_ VGND VGND VPWR VPWR _05156_
+ sky130_fd_sc_hd__and4_1
X_12191_ _03149_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__or2_1
Xoutput43 net43 VGND VGND VPWR VPWR mem_addr[18] sky130_fd_sc_hd__buf_2
X_11142_ net604 _05105_ _05090_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__o21ai_1
Xoutput54 net54 VGND VGND VPWR VPWR mem_addr[29] sky130_fd_sc_hd__clkbuf_4
Xoutput65 net65 VGND VGND VPWR VPWR mem_instr sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput76 net76 VGND VGND VPWR VPWR mem_la_addr[20] sky130_fd_sc_hd__buf_2
Xoutput87 net87 VGND VGND VPWR VPWR mem_la_addr[30] sky130_fd_sc_hd__buf_2
X_11073_ _05059_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__clkbuf_1
X_15950_ clknet_leaf_15_clk _01522_ VGND VGND VPWR VPWR cpuregs\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
Xoutput98 net98 VGND VGND VPWR VPWR mem_la_wdata[10] sky130_fd_sc_hd__clkbuf_4
X_14901_ clknet_leaf_102_clk _00559_ VGND VGND VPWR VPWR count_instr\[10\] sky130_fd_sc_hd__dfxtp_1
X_10024_ _03427_ _04464_ _04466_ _04468_ _03431_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__a221o_1
X_15881_ clknet_leaf_36_clk _01453_ VGND VGND VPWR VPWR cpuregs\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ clknet_leaf_30_clk _00490_ VGND VGND VPWR VPWR cpuregs\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_463 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14763_ clknet_leaf_48_clk _00421_ VGND VGND VPWR VPWR cpuregs\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11975_ _05773_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13714_ net943 _06943_ _07028_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__mux2_1
X_10926_ _04973_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__clkbuf_1
X_14694_ clknet_leaf_126_clk _00352_ VGND VGND VPWR VPWR cpuregs\[27\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10857_ net675 _04844_ _04934_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__mux2_1
X_13645_ _07001_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13576_ _06957_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__clkbuf_1
X_10788_ _04900_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15315_ clknet_leaf_3_clk _00905_ VGND VGND VPWR VPWR cpuregs\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12527_ cpuregs\[28\]\[21\] cpuregs\[29\]\[21\] cpuregs\[30\]\[21\] cpuregs\[31\]\[21\]
+ _06191_ _05914_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15246_ clknet_leaf_76_clk _00839_ VGND VGND VPWR VPWR instr_sub sky130_fd_sc_hd__dfxtp_2
XFILLER_0_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12458_ _03142_ _06205_ _06209_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_111_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11409_ _05290_ _05293_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__nand2_1
X_12389_ _06142_ _06143_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15177_ clknet_leaf_98_clk _00802_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_130_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14128_ net902 _06948_ _01685_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14059_ _01650_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08620_ cpuregs\[12\]\[4\] cpuregs\[13\]\[4\] cpuregs\[14\]\[4\] cpuregs\[15\]\[4\]
+ _03107_ _03137_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__mux4_1
X_08551_ _03033_ _03056_ _03058_ _03070_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__o211a_2
X_07502_ count_instr\[44\] instr_rdinstrh instr_rdcycleh count_cycle\[44\] VGND VGND
+ VPWR VPWR _02142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08482_ _03014_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_18_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_134_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_513 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07433_ _02060_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_628 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07364_ _02007_ _02008_ _02011_ _01927_ _01968_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__a221o_1
X_09103_ _03426_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_44_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07295_ instr_rdcycleh VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_641 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09034_ _03403_ _03503_ _03507_ _03434_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_131_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold320 count_instr\[11\] VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 cpu_state\[0\] VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 cpuregs\[31\]\[7\] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 net168 VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 cpuregs\[20\]\[24\] VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 cpuregs\[0\]\[29\] VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_660 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_159_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold386 cpuregs\[8\]\[10\] VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold397 cpuregs\[28\]\[30\] VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__dlygate4sd3_1
X_09936_ decoded_imm\[27\] net190 VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_148_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ cpuregs\[20\]\[25\] cpuregs\[21\]\[25\] cpuregs\[22\]\[25\] cpuregs\[23\]\[25\]
+ _03438_ _03812_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__mux4_1
Xhold1020 _02504_ VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 cpuregs\[14\]\[5\] VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 count_instr\[48\] VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 count_instr\[24\] VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ _03304_ _03305_ _03293_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__mux2_4
X_09798_ cpuregs\[12\]\[23\] cpuregs\[13\]\[23\] cpuregs\[14\]\[23\] cpuregs\[15\]\[23\]
+ _03516_ _03409_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__mux4_1
*XANTENNA_204 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08749_ _03172_ _03245_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__nor2_1
*XANTENNA_215 _03496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_226 _03581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_237 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11760_ net1402 _05613_ count_cycle\[11\] VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_37_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _04851_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11691_ _05549_ _05562_ _05563_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__o21ai_1
X_13430_ _06872_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__clkbuf_1
X_10642_ _04807_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13361_ net1151 _04856_ _06827_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10573_ net1014 _03329_ _04768_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15100_ clknet_leaf_104_clk _07123_ VGND VGND VPWR VPWR reg_out\[18\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer9 net367 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_1
X_12312_ _06023_ _06069_ _05927_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__o21a_1
X_16080_ net122 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_2
X_13292_ _06799_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15031_ clknet_leaf_132_clk _00689_ VGND VGND VPWR VPWR count_cycle\[14\] sky130_fd_sc_hd__dfxtp_1
X_12243_ cpuregs\[28\]\[9\] cpuregs\[29\]\[9\] cpuregs\[30\]\[9\] cpuregs\[31\]\[9\]
+ _05895_ _05929_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__mux4_1
XFILLER_0_122_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12174_ _05937_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__clkbuf_1
X_11125_ _05095_ _05096_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11056_ count_instr\[4\] _05043_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__nand2_1
X_15933_ clknet_leaf_20_clk _01505_ VGND VGND VPWR VPWR cpuregs\[0\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10007_ _04452_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_1
X_15864_ clknet_leaf_142_clk _01436_ VGND VGND VPWR VPWR cpuregs\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14815_ clknet_leaf_124_clk _00473_ VGND VGND VPWR VPWR cpuregs\[25\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15795_ clknet_leaf_140_clk _01370_ VGND VGND VPWR VPWR cpuregs\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_98_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14746_ clknet_leaf_159_clk _00404_ VGND VGND VPWR VPWR cpuregs\[26\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11958_ _01820_ net235 VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_524 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10909_ _04964_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__clkbuf_1
X_14677_ clknet_leaf_160_clk _00335_ VGND VGND VPWR VPWR cpuregs\[27\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11889_ count_cycle\[50\] net686 count_cycle\[52\] _05700_ VGND VGND VPWR VPWR _05706_
+ sky130_fd_sc_hd__and4_4
XFILLER_0_157_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13628_ net1264 _06923_ _06992_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13559_ _06924_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15229_ clknet_leaf_77_clk _00822_ VGND VGND VPWR VPWR instr_lb sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07982_ _01992_ net251 _02598_ _02563_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__a31o_1
X_09721_ _03672_ _04157_ _04175_ _03665_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09652_ _04107_ _04108_ _03447_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__mux2_1
X_08603_ net522 _03079_ _03121_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__a21oi_1
X_09583_ _03448_ _04041_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_143_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_143_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ _00010_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08465_ reg_next_pc\[25\] reg_out\[25\] _02991_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07416_ _02059_ _02060_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08396_ reg_next_pc\[4\] reg_out\[4\] _02949_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07347_ count_instr\[35\] instr_rdinstrh instr_rdcycleh count_cycle\[35\] VGND VGND
+ VPWR VPWR _01996_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_396 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_547 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07278_ net171 VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_878 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_130_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09017_ cpuregs\[16\]\[1\] cpuregs\[17\]\[1\] cpuregs\[18\]\[1\] cpuregs\[19\]\[1\]
+ _03406_ _03410_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_457 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_14_794 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold150 count_cycle\[28\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 count_cycle\[36\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 count_cycle\[10\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 count_cycle\[6\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold194 cpuregs\[5\]\[3\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
X_09919_ cpuregs\[12\]\[27\] cpuregs\[13\]\[27\] cpuregs\[14\]\[27\] cpuregs\[15\]\[27\]
+ _03719_ _03588_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__mux4_1
X_12930_ mem_rdata_q\[30\] net24 _06589_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__mux2_1
X_12861_ _06546_ _06547_ _06559_ _06562_ net472 VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__a32o_1
X_14600_ clknet_leaf_24_clk _00258_ VGND VGND VPWR VPWR cpuregs\[28\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11812_ _05654_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ clknet_leaf_136_clk _01155_ VGND VGND VPWR VPWR cpuregs\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12792_ _06520_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__buf_1
XFILLER_0_95_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14531_ clknet_leaf_98_clk _00189_ VGND VGND VPWR VPWR cpuregs\[13\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11743_ _05606_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14462_ clknet_leaf_137_clk _00120_ VGND VGND VPWR VPWR cpuregs\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11674_ _05251_ _05540_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13413_ net998 _04839_ _06863_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10625_ _04798_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14393_ clknet_leaf_14_clk _00056_ VGND VGND VPWR VPWR cpuregs\[11\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10556_ cpuregs\[27\]\[14\] _03275_ _04757_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__mux2_1
X_13344_ _06815_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__buf_4
XFILLER_0_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpicorv32_308 VGND VGND VPWR VPWR picorv32_308/HI pcpi_insn[18] sky130_fd_sc_hd__conb_1
Xpicorv32_319 VGND VGND VPWR VPWR picorv32_319/HI pcpi_insn[29] sky130_fd_sc_hd__conb_1
X_10487_ net1270 _03275_ _04720_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__mux2_1
X_13275_ _06790_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15014_ clknet_leaf_106_clk _00672_ VGND VGND VPWR VPWR reg_next_pc\[29\] sky130_fd_sc_hd__dfxtp_1
X_12226_ _05886_ _05972_ _05977_ _05978_ _05987_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__a311o_1
XFILLER_0_121_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12157_ _03051_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__buf_8
X_11108_ _05083_ _05084_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__nor2_1
X_12088_ cpuregs\[28\]\[1\] cpuregs\[29\]\[1\] cpuregs\[30\]\[1\] cpuregs\[31\]\[1\]
+ _05816_ _03086_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__mux4_1
X_11039_ _05031_ _05032_ count_instr\[0\] VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__a21o_1
X_15916_ clknet_leaf_11_clk _01488_ VGND VGND VPWR VPWR cpuregs\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_160_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ clknet_leaf_41_clk _01419_ VGND VGND VPWR VPWR cpuregs\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_125_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ clknet_leaf_40_clk _01353_ VGND VGND VPWR VPWR cpuregs\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14729_ clknet_leaf_21_clk _00387_ VGND VGND VPWR VPWR cpuregs\[15\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08250_ net186 _02837_ _02829_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_129_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07201_ mem_do_rdata net34 cpu_state\[6\] _01862_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__and4b_2
XFILLER_0_28_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08181_ net212 _02782_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput200 net200 VGND VGND VPWR VPWR pcpi_rs1[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput211 net211 VGND VGND VPWR VPWR pcpi_rs2[17] sky130_fd_sc_hd__clkbuf_4
Xoutput222 net222 VGND VGND VPWR VPWR pcpi_rs2[27] sky130_fd_sc_hd__clkbuf_4
Xoutput233 net233 VGND VGND VPWR VPWR pcpi_rs2[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07965_ _02579_ _02580_ _02583_ net1379 VGND VGND VPWR VPWR alu_out\[1\] sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_145_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09704_ cpuregs\[20\]\[20\] cpuregs\[21\]\[20\] cpuregs\[22\]\[20\] cpuregs\[23\]\[20\]
+ _03719_ _03450_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07896_ _02511_ _02513_ _02514_ _02515_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__a2bb2o_1
X_09635_ _02213_ net243 VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09566_ _04022_ _04023_ _04024_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08517_ _03036_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09497_ _02222_ _03481_ _03888_ _03075_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08448_ _02990_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_148_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08379_ net223 _02252_ _02932_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__a21o_1
XFILLER_0_46_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_817 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10410_ _04672_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11390_ _05258_ net1138 _05239_ _05287_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10341_ _04635_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_59_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13060_ net1121 _04879_ _06658_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10272_ _04610_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_596 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12011_ _05792_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13962_ _01598_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__clkbuf_1
X_15701_ clknet_leaf_142_clk _01276_ VGND VGND VPWR VPWR cpuregs\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_12913_ _06591_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
X_13893_ _01561_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ clknet_leaf_0_clk _01207_ VGND VGND VPWR VPWR cpuregs\[23\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12844_ mem_rdata_q\[14\] _06536_ mem_rdata_q\[12\] VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__or3_2
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15563_ clknet_leaf_4_clk _01138_ VGND VGND VPWR VPWR cpuregs\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12775_ instr_lh _01928_ _06509_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__a21bo_1
X_14514_ clknet_leaf_56_clk _00172_ VGND VGND VPWR VPWR cpuregs\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ reg_next_pc\[31\] _05031_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ clknet_leaf_94_clk _01079_ VGND VGND VPWR VPWR mem_rdata_q\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14445_ clknet_leaf_39_clk _00103_ VGND VGND VPWR VPWR cpuregs\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11657_ _05494_ _05246_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10608_ _04789_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14376_ clknet_leaf_26_clk _00039_ VGND VGND VPWR VPWR cpuregs\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11588_ _05418_ net517 _05343_ _05469_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold908 cpuregs\[5\]\[27\] VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13327_ _06818_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__clkbuf_1
Xhold919 cpuregs\[30\]\[17\] VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10539_ net981 _03221_ _04746_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_122_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13258_ net842 _04821_ _06780_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__mux2_1
X_12209_ cpuregs\[24\]\[8\] cpuregs\[25\]\[8\] cpuregs\[26\]\[8\] cpuregs\[27\]\[8\]
+ _05970_ _03137_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__mux4_1
X_13189_ mem_rdata_q\[29\] _06742_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_127_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07750_ _02018_ _02363_ _02372_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__o21a_1
X_07681_ _02304_ _02305_ _02308_ _02018_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_140_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09420_ _03414_ _03883_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09351_ cpuregs\[28\]\[9\] cpuregs\[29\]\[9\] cpuregs\[30\]\[9\] cpuregs\[31\]\[9\]
+ _03456_ _03441_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08302_ _02892_ _02893_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09282_ _03593_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08233_ _02829_ _02830_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_51_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08164_ _02539_ _02569_ _02767_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_138_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_889 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08095_ _02463_ _02702_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_703 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08997_ decoded_imm_j\[19\] _03471_ is_lui_auipc_jal VGND VGND VPWR VPWR _03472_
+ sky130_fd_sc_hd__o21ba_2
X_07948_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07879_ _02008_ net250 VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__nand2_1
X_09618_ _03488_ _04075_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10890_ net730 _04877_ _04945_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09549_ _03616_ _04007_ _04008_ _01942_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12560_ _06132_ _06294_ _06307_ _06153_ decoded_imm\[22\] VGND VGND VPWR VPWR _06308_
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_102_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_650 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11511_ decoded_imm_j\[12\] _05395_ _05397_ _05398_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__a211o_1
X_12491_ _06235_ _06237_ _06239_ _06241_ _06151_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__a221o_2
XFILLER_0_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14230_ _01740_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11442_ _05333_ _05334_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_839 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14161_ cpuregs\[7\]\[27\] _06981_ _01696_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__mux2_1
X_11373_ decoded_imm_j\[1\] _05187_ _05270_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__nand3_2
XFILLER_0_132_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13112_ net138 net100 _06696_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__mux2_1
X_10324_ _04638_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14092_ _01667_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13043_ _06659_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__clkbuf_1
X_10255_ cpuregs\[2\]\[1\] _03189_ _04600_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_780 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10186_ _04565_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14994_ clknet_leaf_86_clk _00652_ VGND VGND VPWR VPWR reg_next_pc\[9\] sky130_fd_sc_hd__dfxtp_1
X_13945_ cpuregs\[4\]\[21\] _06969_ _01588_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13876_ net593 _06969_ _01551_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__mux2_1
X_15615_ clknet_leaf_54_clk _01190_ VGND VGND VPWR VPWR cpuregs\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12827_ _05040_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15546_ clknet_leaf_80_clk _00019_ VGND VGND VPWR VPWR cpu_state\[2\] sky130_fd_sc_hd__dfxtp_1
X_12758_ cpuregs\[24\]\[31\] cpuregs\[25\]\[31\] cpuregs\[26\]\[31\] cpuregs\[27\]\[31\]
+ _03150_ _03151_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11709_ _05495_ _05259_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nand2_1
X_15477_ clknet_leaf_78_clk _01062_ VGND VGND VPWR VPWR mem_rdata_q\[0\] sky130_fd_sc_hd__dfxtp_1
X_12689_ cpuregs\[28\]\[28\] cpuregs\[29\]\[28\] cpuregs\[30\]\[28\] cpuregs\[31\]\[28\]
+ _06191_ _05914_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14428_ clknet_leaf_59_clk _00086_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14359_ net750 _03354_ _01800_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__mux2_1
Xhold705 cpuregs\[13\]\[2\] VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold716 cpuregs\[26\]\[13\] VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 cpuregs\[28\]\[24\] VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold738 cpuregs\[14\]\[1\] VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 cpuregs\[23\]\[16\] VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08920_ _03394_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08851_ net607 _03334_ _03315_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__mux2_1
X_07802_ _02410_ _02411_ _02412_ _02421_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__a22o_1
X_08782_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__clkbuf_4
X_07733_ _02353_ _02356_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__xor2_1
X_07664_ _02058_ _02289_ _02292_ _01968_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09403_ _03833_ _03836_ _03865_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07595_ _02225_ _02228_ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09334_ _00012_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__buf_6
XFILLER_0_118_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09265_ _02044_ _03624_ _03733_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__a21o_1
XFILLER_0_161_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_688 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08216_ net216 _02814_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_474 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09196_ _02008_ _03624_ _03666_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_658 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08147_ _02704_ _02718_ _02733_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08078_ _02112_ net248 _02618_ _02641_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10040_ _01877_ _04482_ _03181_ _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__or4b_1
Xhold54 mem_rdata[29] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 mem_rdata[9] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 count_cycle\[1\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 mem_rdata_q\[31\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _00558_ VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11991_ net40 net71 _05774_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13730_ _07046_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__clkbuf_1
X_10942_ cpuregs\[20\]\[20\] _04860_ _04981_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13661_ net1108 _06958_ _07003_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__mux2_1
X_10873_ _04922_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15400_ clknet_leaf_90_clk _00990_ VGND VGND VPWR VPWR decoded_imm\[8\] sky130_fd_sc_hd__dfxtp_2
X_12612_ _06142_ _06356_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13592_ _06968_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15331_ clknet_leaf_73_clk _00921_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12543_ cpuregs\[8\]\[22\] cpuregs\[9\]\[22\] cpuregs\[10\]\[22\] cpuregs\[11\]\[22\]
+ _05907_ _03039_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15262_ clknet_leaf_85_clk _00855_ VGND VGND VPWR VPWR decoded_imm_j\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_409 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12474_ _06225_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_910 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14213_ _01731_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__clkbuf_1
X_11425_ _05263_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15193_ clknet_leaf_70_clk alu_out\[6\] VGND VGND VPWR VPWR alu_out_q\[6\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_7 _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14144_ net1362 _06964_ _01685_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__mux2_1
X_11356_ _05193_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_120_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10307_ net1207 _03355_ _04622_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__mux2_1
X_14075_ _01658_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__clkbuf_1
X_11287_ _05186_ _05208_ _05209_ _01885_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__o211a_1
X_13026_ _06650_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__clkbuf_1
X_10238_ _04592_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__clkbuf_1
X_10169_ cpuregs\[30\]\[26\] _03355_ _04548_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__mux2_1
X_14977_ clknet_leaf_112_clk _00635_ VGND VGND VPWR VPWR reg_pc\[23\] sky130_fd_sc_hd__dfxtp_2
Xrebuffer19 _05655_ VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13928_ cpuregs\[4\]\[13\] _06952_ _01577_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13859_ net1288 _06952_ _07111_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07380_ _01988_ _01975_ _01986_ _02000_ _02002_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__o311a_1
XFILLER_0_45_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15529_ clknet_leaf_147_clk _01114_ VGND VGND VPWR VPWR cpuregs\[24\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09050_ _03474_ _03488_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08001_ _02614_ _02615_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold502 cpuregs\[10\]\[8\] VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold513 cpuregs\[21\]\[15\] VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold524 instr_bne VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold535 cpuregs\[11\]\[29\] VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold546 cpuregs\[11\]\[19\] VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 cpuregs\[15\]\[8\] VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold568 cpuregs\[15\]\[24\] VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 cpuregs\[2\]\[13\] VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ decoded_imm\[26\] _02331_ _04384_ _04398_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_0_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08903_ _03261_ _03376_ _03377_ _03379_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_51_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _02316_ _04332_ _03395_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__mux2_1
X_08834_ _03318_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__nor2_1
X_08765_ _03258_ _03259_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__nor2_1
X_07716_ net20 _02202_ _02180_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__a21o_1
X_08696_ reg_pc\[3\] _01971_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_637 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07647_ net185 VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_49_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_542 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_94_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07578_ net179 VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09317_ cpuregs\[20\]\[8\] cpuregs\[21\]\[8\] cpuregs\[22\]\[8\] cpuregs\[23\]\[8\]
+ _03636_ _03637_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09248_ cpuregs\[24\]\[6\] cpuregs\[25\]\[6\] cpuregs\[26\]\[6\] cpuregs\[27\]\[6\]
+ _03582_ _03716_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_145_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
X_09179_ _03474_ _03635_ _03649_ _03527_ reg_pc\[4\] VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11210_ _05153_ _05151_ _05155_ _05052_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_120_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12190_ cpuregs\[24\]\[7\] cpuregs\[25\]\[7\] cpuregs\[26\]\[7\] cpuregs\[27\]\[7\]
+ _03095_ _05932_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11141_ count_instr\[29\] count_instr\[28\] _05103_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__and3_1
Xoutput44 net44 VGND VGND VPWR VPWR mem_addr[19] sky130_fd_sc_hd__buf_2
Xoutput55 net55 VGND VGND VPWR VPWR mem_addr[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput66 net66 VGND VGND VPWR VPWR mem_la_addr[10] sky130_fd_sc_hd__clkbuf_4
Xoutput77 net77 VGND VGND VPWR VPWR mem_la_addr[21] sky130_fd_sc_hd__buf_2
X_11072_ _01905_ _05057_ _05058_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__and3_1
Xoutput88 net88 VGND VGND VPWR VPWR mem_la_addr[31] sky130_fd_sc_hd__buf_2
Xoutput99 net99 VGND VGND VPWR VPWR mem_la_wdata[11] sky130_fd_sc_hd__clkbuf_4
X_14900_ clknet_leaf_113_clk net457 VGND VGND VPWR VPWR count_instr\[9\] sky130_fd_sc_hd__dfxtp_1
X_10023_ _03448_ _04467_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__or2_1
X_15880_ clknet_leaf_33_clk _01452_ VGND VGND VPWR VPWR cpuregs\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_14831_ clknet_leaf_38_clk _00489_ VGND VGND VPWR VPWR cpuregs\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ clknet_leaf_46_clk _00420_ VGND VGND VPWR VPWR cpuregs\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11974_ net919 net93 _05767_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13713_ _07037_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__clkbuf_1
X_10925_ cpuregs\[20\]\[12\] _04844_ _04970_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__mux2_1
X_14693_ clknet_leaf_153_clk _00351_ VGND VGND VPWR VPWR cpuregs\[27\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_542 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13644_ net680 _06941_ _06992_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__mux2_1
X_10856_ _04936_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13575_ net1114 _06956_ _06946_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10787_ net1249 _04842_ _04898_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_463 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_143_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15314_ clknet_leaf_16_clk _00904_ VGND VGND VPWR VPWR cpuregs\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12526_ _06023_ _06274_ _05840_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_720 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15245_ clknet_leaf_80_clk _00838_ VGND VGND VPWR VPWR instr_add sky130_fd_sc_hd__dfxtp_1
X_12457_ _05845_ _06206_ _06208_ _03139_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_280 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_124_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11408_ _05302_ _05303_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__and2_1
X_15176_ clknet_leaf_98_clk _00801_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_97_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12388_ cpuregs\[20\]\[15\] cpuregs\[21\]\[15\] cpuregs\[22\]\[15\] cpuregs\[23\]\[15\]
+ _06065_ _05922_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__mux4_1
X_14127_ _01686_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11339_ reg_next_pc\[25\] _03343_ _02948_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_130_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14058_ cpuregs\[6\]\[10\] _06945_ _01649_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__mux2_1
X_13009_ _06641_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08550_ _03060_ _03065_ _03069_ _00011_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__a211o_1
X_07501_ _02083_ _02140_ _02085_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_18_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08481_ _02380_ _03013_ _02993_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_648 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_134_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07432_ _02060_ _02063_ _02059_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_147_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_726 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07363_ net27 net130 _02010_ _01940_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09102_ _03473_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07294_ instr_rdinstrh VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_44_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_150_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09033_ _03410_ _03504_ _03506_ _03415_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold310 instr_srl VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 cpuregs\[23\]\[8\] VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold332 count_cycle\[61\] VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold343 cpuregs\[0\]\[2\] VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold354 cpuregs\[2\]\[31\] VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 cpuregs\[15\]\[26\] VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 cpuregs\[31\]\[28\] VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 cpuregs\[0\]\[25\] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 cpuregs\[8\]\[13\] VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ _03657_ _04269_ _04380_ _04382_ _01942_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_148_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _03547_ _04311_ _04313_ _04315_ _00016_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__a221o_1
Xhold1010 cpuregs\[18\]\[28\] VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 cpuregs\[16\]\[12\] VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1032 cpuregs\[23\]\[18\] VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ reg_pc\[19\] _03299_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__xor2_1
Xhold1043 count_cycle\[10\] VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 count_instr\[37\] VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _03437_ _04248_ _03419_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__o21a_1
X_08748_ reg_pc\[10\] reg_pc\[9\] _03232_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__and3_1
*XANTENNA_205 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_216 _03547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_227 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_238 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08679_ net816 _03179_ _03185_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_503 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ cpuregs\[26\]\[15\] _04850_ _04840_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _05494_ _05253_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_81_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10641_ net684 _03329_ _04804_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13360_ _06835_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__clkbuf_1
X_10572_ _04770_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_742 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12311_ cpuregs\[16\]\[12\] cpuregs\[17\]\[12\] cpuregs\[18\]\[12\] cpuregs\[19\]\[12\]
+ _05948_ _06068_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_792 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13291_ net1315 _04854_ _06791_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15030_ clknet_leaf_132_clk _00688_ VGND VGND VPWR VPWR count_cycle\[13\] sky130_fd_sc_hd__dfxtp_1
X_12242_ _03090_ _06002_ _05927_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_79_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12173_ _02492_ _05936_ _05863_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11124_ net518 _05092_ _05090_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__o21ai_1
X_11055_ count_instr\[4\] _05043_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__or2_1
X_15932_ clknet_leaf_17_clk _01504_ VGND VGND VPWR VPWR cpuregs\[0\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_10006_ _02369_ _04451_ _03394_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__mux2_1
X_15863_ clknet_leaf_133_clk _01435_ VGND VGND VPWR VPWR cpuregs\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14814_ clknet_leaf_147_clk _00472_ VGND VGND VPWR VPWR cpuregs\[25\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15794_ clknet_leaf_16_clk _01369_ VGND VGND VPWR VPWR cpuregs\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14745_ clknet_leaf_160_clk _00403_ VGND VGND VPWR VPWR cpuregs\[26\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11957_ _05761_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_58_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10908_ cpuregs\[20\]\[4\] _04827_ _04959_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__mux2_1
X_14676_ clknet_leaf_2_clk _00334_ VGND VGND VPWR VPWR cpuregs\[27\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11888_ net447 _05703_ _05705_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_67_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13627_ _06991_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10839_ _04927_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13558_ _03247_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_81_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12509_ cpuregs\[24\]\[20\] cpuregs\[25\]\[20\] cpuregs\[26\]\[20\] cpuregs\[27\]\[20\]
+ _06074_ _03151_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_764 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13489_ cpuregs\[9\]\[14\] _04848_ _06899_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__mux2_1
X_15228_ clknet_leaf_78_clk _00821_ VGND VGND VPWR VPWR instr_jalr sky130_fd_sc_hd__dfxtp_2
XFILLER_0_23_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_50_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15159_ clknet_leaf_49_clk _00784_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dfxtp_2
X_07981_ _02560_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__clkbuf_4
X_09720_ reg_pc\[20\] _03528_ _04174_ _03626_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__a211o_1
X_09651_ cpuregs\[0\]\[18\] cpuregs\[1\]\[18\] cpuregs\[2\]\[18\] cpuregs\[3\]\[18\]
+ _03463_ _03464_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__mux4_1
X_08602_ is_slli_srli_srai _03119_ _03120_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__o21a_1
X_09582_ cpuregs\[12\]\[16\] cpuregs\[13\]\[16\] cpuregs\[14\]\[16\] cpuregs\[15\]\[16\]
+ _03680_ _03443_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_89_250 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08533_ cpuregs\[28\]\[2\] cpuregs\[29\]\[2\] cpuregs\[30\]\[2\] cpuregs\[31\]\[2\]
+ _03051_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ _03002_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_46_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07415_ reg_pc\[7\] decoded_imm\[7\] VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_843 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08395_ _02954_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_1
XFILLER_0_18_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07346_ net26 net130 _01994_ _01940_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07277_ _01844_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_263 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_131_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09016_ _03489_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__buf_6
XFILLER_0_115_285 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_131_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_469 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold140 count_instr\[57\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 decoded_imm_j\[17\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 reg_sh\[4\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _00685_ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 reg_next_pc\[16\] VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 count_instr\[46\] VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ _03581_ _04365_ _03467_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__o21a_1
X_09849_ _03434_ _04295_ _04297_ _04299_ _03431_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__a221o_1
X_12860_ _06546_ _06543_ _06559_ _06562_ net624 VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_913 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11811_ _05652_ _05625_ _05653_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_1_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12791_ mem_rdata_q\[6\] net29 _01857_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14530_ clknet_leaf_137_clk _00188_ VGND VGND VPWR VPWR cpuregs\[13\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11742_ _05604_ _05113_ _05605_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__and3b_1
XFILLER_0_96_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14461_ clknet_leaf_13_clk _00119_ VGND VGND VPWR VPWR cpuregs\[12\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11673_ _05418_ net813 _05358_ _05547_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13412_ _06851_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__buf_4
X_10624_ cpuregs\[15\]\[14\] _03275_ _04793_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14392_ clknet_leaf_15_clk _00055_ VGND VGND VPWR VPWR cpuregs\[11\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13343_ _06826_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__clkbuf_1
X_10555_ _04761_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xpicorv32_309 VGND VGND VPWR VPWR picorv32_309/HI pcpi_insn[19] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_20_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13274_ cpuregs\[18\]\[9\] _04837_ _06780_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__mux2_1
X_10486_ _04724_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_94_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_907 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15013_ clknet_leaf_109_clk _00671_ VGND VGND VPWR VPWR reg_next_pc\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12225_ _05981_ _05983_ _05986_ _03132_ _05815_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__o221a_1
X_12156_ _05879_ _05911_ _05916_ _05919_ _03104_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__a221o_2
X_11107_ net1178 _05082_ _05044_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__o21ai_1
X_12087_ _03128_ _05855_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__nor2_1
X_11038_ _05031_ count_instr\[0\] _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__and3_1
X_15915_ clknet_leaf_31_clk _01487_ VGND VGND VPWR VPWR cpuregs\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_160_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15846_ clknet_leaf_47_clk _01418_ VGND VGND VPWR VPWR cpuregs\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_125_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15777_ clknet_leaf_26_clk _01352_ VGND VGND VPWR VPWR cpuregs\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12989_ _01067_ _06631_ is_lb_lh_lw_lbu_lhu _06513_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_87_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14728_ clknet_leaf_59_clk _00386_ VGND VGND VPWR VPWR cpuregs\[15\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14659_ clknet_leaf_97_clk _00317_ VGND VGND VPWR VPWR cpuregs\[14\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07200_ mem_do_prefetch _01854_ _01860_ _01864_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08180_ net211 net247 _02759_ _02656_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__o31a_1
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_65_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_518 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput201 net201 VGND VGND VPWR VPWR pcpi_rs1[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput212 net212 VGND VGND VPWR VPWR pcpi_rs2[18] sky130_fd_sc_hd__buf_2
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput223 net223 VGND VGND VPWR VPWR pcpi_rs2[28] sky130_fd_sc_hd__buf_2
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput234 net234 VGND VGND VPWR VPWR pcpi_rs2[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07964_ _02505_ _02581_ _02582_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_145_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09703_ cpuregs\[16\]\[20\] cpuregs\[17\]\[20\] cpuregs\[18\]\[20\] cpuregs\[19\]\[20\]
+ _03587_ _03588_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_74_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07895_ _01992_ net251 VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09634_ _02165_ _02277_ _03619_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__mux2_1
X_09565_ decoded_imm\[16\] _02200_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08516_ _00009_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09496_ _03957_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__clkbuf_1
X_08447_ _02250_ _02989_ _02971_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_768 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_83_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08378_ net222 _02252_ _02931_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__a21o_2
XFILLER_0_73_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07329_ net2 net19 _01845_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10340_ _04646_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10271_ net993 _03241_ _04600_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__mux2_1
X_12010_ net49 net80 _05785_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13961_ cpuregs\[4\]\[29\] _06985_ _01588_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__mux2_1
X_15700_ clknet_leaf_133_clk _01275_ VGND VGND VPWR VPWR cpuregs\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12912_ decoded_imm_j\[5\] _01087_ _03169_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__mux2_1
X_13892_ net1177 _06985_ _01551_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ clknet_leaf_0_clk _01206_ VGND VGND VPWR VPWR cpuregs\[23\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12843_ instr_lh _06554_ _06539_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _00823_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_551 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15562_ clknet_leaf_5_clk _01137_ VGND VGND VPWR VPWR cpuregs\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12774_ mem_do_rdata _01927_ _06508_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_139_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14513_ clknet_leaf_34_clk _00171_ VGND VGND VPWR VPWR cpuregs\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11725_ _05261_ _05594_ _05032_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15493_ clknet_leaf_94_clk _01078_ VGND VGND VPWR VPWR mem_rdata_q\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_120_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ clknet_leaf_24_clk _00102_ VGND VGND VPWR VPWR cpuregs\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11656_ _05486_ _05518_ _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__and3b_1
XFILLER_0_154_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_695 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10607_ net892 _03221_ _04782_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14375_ clknet_leaf_51_clk _00038_ VGND VGND VPWR VPWR cpuregs\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11587_ _05269_ _05466_ _05468_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13326_ net681 _04821_ _06816_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__mux2_1
X_10538_ _04752_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__clkbuf_1
Xhold909 cpuregs\[26\]\[1\] VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13257_ _06781_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10469_ _04715_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__clkbuf_1
X_12208_ _03046_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__buf_8
X_13188_ _01823_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__buf_2
X_12139_ _01918_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_127_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07680_ _02007_ _02306_ _02183_ _02307_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_140_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15829_ clknet_leaf_3_clk _01401_ VGND VGND VPWR VPWR cpuregs\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_140_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_59_242 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09350_ _03557_ _03815_ _03425_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08301_ _02869_ _02876_ _02884_ _02886_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__a31o_1
XFILLER_0_157_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09281_ cpuregs\[12\]\[7\] cpuregs\[13\]\[7\] cpuregs\[14\]\[7\] cpuregs\[15\]\[7\]
+ _03594_ _03595_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_153_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_153_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_129_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08232_ net185 _02828_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_684 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08163_ _02200_ net247 _02618_ _02641_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_138_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08094_ _02656_ _02701_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08996_ decoded_imm_j\[18\] decoded_imm_j\[17\] decoded_imm_j\[16\] decoded_imm_j\[15\]
+ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_3_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ instr_xor instr_xori VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__or2_1
X_07878_ _02008_ net250 VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__or2_1
X_09617_ _03574_ _04065_ _04074_ _03527_ reg_pc\[17\] VGND VGND VPWR VPWR _04075_
+ sky130_fd_sc_hd__a32o_1
X_09548_ _02237_ _03480_ _03904_ _03074_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_144_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_144_clk sky130_fd_sc_hd__clkbuf_2
X_09479_ cpuregs\[20\]\[13\] cpuregs\[21\]\[13\] cpuregs\[22\]\[13\] cpuregs\[23\]\[13\]
+ _03438_ _03812_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11510_ decoded_imm_j\[12\] _05395_ _05372_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_22_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_336 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12490_ _06073_ _06240_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11441_ decoded_imm_j\[8\] _05206_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14160_ _01703_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__clkbuf_1
X_11372_ decoded_imm_j\[1\] _05187_ _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13111_ _06698_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10323_ net876 _03189_ _04636_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__mux2_1
X_14091_ cpuregs\[6\]\[26\] _06979_ _01660_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13042_ net1386 _04860_ _06658_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__mux2_1
X_10254_ _04601_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10185_ net1020 _03179_ _04564_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14993_ clknet_leaf_84_clk _00651_ VGND VGND VPWR VPWR reg_next_pc\[8\] sky130_fd_sc_hd__dfxtp_1
X_13944_ _01589_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13875_ _01552_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15614_ clknet_leaf_17_clk _01189_ VGND VGND VPWR VPWR cpuregs\[31\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12826_ net500 _06530_ _06545_ _05804_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12757_ _05912_ _06495_ _06193_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__o21a_1
X_15545_ clknet_leaf_79_clk _00018_ VGND VGND VPWR VPWR cpu_state\[1\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_135_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_135_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_155_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_139_483 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_84_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11708_ _05571_ _05574_ _05572_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__o21ai_1
X_15476_ clknet_leaf_98_clk _00036_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__dfxtp_2
X_12688_ _03132_ _06429_ _05840_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14427_ clknet_leaf_60_clk _00085_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dfxtp_2
X_11639_ _05263_ net933 _05514_ _05516_ _01843_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__o221a_1
XFILLER_0_108_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14358_ _01806_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_613 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold706 cpuregs\[1\]\[8\] VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold717 cpuregs\[3\]\[9\] VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold728 cpuregs\[26\]\[18\] VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ _06808_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_139_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14289_ net746 VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__clkbuf_1
Xhold739 cpuregs\[8\]\[6\] VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08850_ _03333_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07801_ _02415_ _02420_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__or2_1
X_08781_ _03270_ _03273_ _03261_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__mux2_4
XFILLER_0_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07732_ _02354_ _02355_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07663_ _01943_ _02290_ _02184_ _02291_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_148_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09402_ _03833_ _03836_ _03865_ _01870_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07594_ count_cycle\[18\] _02051_ _02227_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09333_ _03796_ _03797_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_126_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_126_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09264_ _03665_ _03712_ _03732_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_749 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08215_ instr_sub net383 VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_401 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09195_ _03626_ _03650_ _03664_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08146_ _02732_ _02746_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08077_ _02682_ _02685_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_567 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08979_ _03401_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__clkbuf_8
Xhold55 net34 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 mem_rdata[22] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 decoded_rd\[4\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 count_cycle\[51\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11990_ _05781_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__clkbuf_1
Xhold99 count_instr\[49\] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _04958_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_27_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13660_ _07009_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10872_ _04944_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_735 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12611_ cpuregs\[20\]\[25\] cpuregs\[21\]\[25\] cpuregs\[22\]\[25\] cpuregs\[23\]\[25\]
+ _06065_ _03144_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_84_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13591_ net1092 _06966_ _06967_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_117_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_117_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15330_ clknet_leaf_73_clk _00920_ VGND VGND VPWR VPWR is_compare sky130_fd_sc_hd__dfxtp_1
X_12542_ cpuregs\[12\]\[22\] cpuregs\[13\]\[22\] cpuregs\[14\]\[22\] cpuregs\[15\]\[22\]
+ _05834_ _03129_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15261_ clknet_leaf_90_clk _00854_ VGND VGND VPWR VPWR decoded_imm_j\[4\] sky130_fd_sc_hd__dfxtp_2
X_12473_ net212 _06224_ _06052_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__mux2_1
X_14212_ net1187 _06964_ _01721_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__mux2_1
X_11424_ _05201_ _05308_ _05318_ _05032_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_50_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15192_ clknet_leaf_73_clk alu_out\[5\] VGND VGND VPWR VPWR alu_out_q\[5\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_8 _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14143_ _01694_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_529 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11355_ _05227_ _05255_ _05256_ _05257_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10306_ _04628_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__clkbuf_1
X_14074_ net1168 _06962_ _01649_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__mux2_1
X_11286_ _05188_ reg_pc\[9\] VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__or2_1
X_13025_ net1312 _04844_ _06647_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__mux2_1
X_10237_ net1062 _03348_ _04586_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__mux2_1
X_10168_ _04554_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__clkbuf_1
X_14976_ clknet_leaf_109_clk _00634_ VGND VGND VPWR VPWR reg_pc\[22\] sky130_fd_sc_hd__dfxtp_2
X_10099_ _04516_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__clkbuf_1
X_13927_ _01580_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__clkbuf_1
X_13858_ _01543_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_157_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12809_ mem_rdata_q\[14\] VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_108_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_108_clk sky130_fd_sc_hd__clkbuf_2
X_13789_ cpuregs\[3\]\[12\] _06950_ _07075_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15528_ clknet_leaf_157_clk _01113_ VGND VGND VPWR VPWR cpuregs\[24\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_913 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15459_ clknet_leaf_157_clk _01049_ VGND VGND VPWR VPWR cpuregs\[19\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08000_ _02614_ _02615_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_618 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold503 cpuregs\[12\]\[1\] VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 cpuregs\[25\]\[26\] VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 cpuregs\[25\]\[22\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 cpuregs\[19\]\[2\] VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 cpuregs\[7\]\[28\] VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09951_ decoded_imm\[27\] _02340_ _04282_ _04396_ _04397_ VGND VGND VPWR VPWR _04398_
+ sky130_fd_sc_hd__a221o_1
Xhold558 cpuregs\[17\]\[30\] VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 cpuregs\[13\]\[19\] VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08902_ _03172_ _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_148_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09882_ _03651_ _04307_ _04308_ _04327_ _04331_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_51_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ reg_pc\[21\] _03311_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08764_ reg_pc\[12\] reg_pc\[11\] _03245_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__and3_1
X_07715_ net190 VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__buf_4
X_08695_ _03198_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__buf_2
X_07646_ _01945_ _02274_ _02275_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07577_ _02210_ _02211_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09316_ cpuregs\[16\]\[8\] cpuregs\[17\]\[8\] cpuregs\[18\]\[8\] cpuregs\[19\]\[8\]
+ _03636_ _03642_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09247_ _03408_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__buf_4
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_911 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09178_ _03639_ _03644_ _03648_ _03434_ _03431_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08129_ _02732_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11140_ _05105_ _05106_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput45 net45 VGND VGND VPWR VPWR mem_addr[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput56 net56 VGND VGND VPWR VPWR mem_addr[30] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VGND VGND VPWR VPWR mem_la_addr[11] sky130_fd_sc_hd__clkbuf_4
Xoutput78 net78 VGND VGND VPWR VPWR mem_la_addr[22] sky130_fd_sc_hd__clkbuf_4
X_11071_ count_instr\[8\] _05055_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__nand2_1
Xoutput89 net89 VGND VGND VPWR VPWR mem_la_addr[3] sky130_fd_sc_hd__clkbuf_4
X_10022_ cpuregs\[28\]\[30\] cpuregs\[29\]\[30\] cpuregs\[30\]\[30\] cpuregs\[31\]\[30\]
+ _03440_ _03451_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__mux4_1
X_14830_ clknet_leaf_44_clk _00488_ VGND VGND VPWR VPWR cpuregs\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ clknet_leaf_18_clk _00419_ VGND VGND VPWR VPWR cpuregs\[26\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_11973_ _05772_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10924_ _04972_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__clkbuf_1
X_13712_ cpuregs\[29\]\[8\] _06941_ _07028_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__mux2_1
X_14692_ clknet_leaf_150_clk _00350_ VGND VGND VPWR VPWR cpuregs\[27\]\[26\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10855_ net1073 _04842_ _04934_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13643_ _07000_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13574_ _03281_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10786_ _04899_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__clkbuf_1
X_12525_ cpuregs\[16\]\[21\] cpuregs\[17\]\[21\] cpuregs\[18\]\[21\] cpuregs\[19\]\[21\]
+ _05984_ _06068_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__mux4_1
X_15313_ clknet_leaf_6_clk _00903_ VGND VGND VPWR VPWR cpuregs\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_732 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_35_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12456_ _03042_ _06207_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__or2_1
X_15244_ clknet_leaf_79_clk _00837_ VGND VGND VPWR VPWR instr_srli sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_292 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11407_ decoded_imm_j\[5\] _05199_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15175_ clknet_leaf_98_clk _00800_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_140_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12387_ _03050_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14126_ cpuregs\[7\]\[10\] _06945_ _01685_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11338_ _05194_ reg_pc\[24\] _05239_ _05245_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_130_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14057_ _01637_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__buf_4
X_11269_ reg_next_pc\[4\] _03204_ _02945_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__mux2_2
XFILLER_0_94_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13008_ net807 _04827_ _06636_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14959_ clknet_leaf_82_clk _00617_ VGND VGND VPWR VPWR reg_pc\[5\] sky130_fd_sc_hd__dfxtp_2
X_07500_ _01846_ _01848_ net21 _01933_ net4 VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__a32o_1
X_08480_ reg_next_pc\[30\] reg_out\[30\] _02991_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07431_ _02073_ _02074_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_885 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_91_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07362_ net13 _01937_ _02009_ _01935_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09101_ _03573_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07293_ cpu_state\[3\] VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09032_ _03493_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold300 cpuregs\[29\]\[14\] VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_798 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold311 cpuregs\[3\]\[28\] VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 cpuregs\[19\]\[1\] VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 cpuregs\[26\]\[19\] VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold344 count_instr\[42\] VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 cpuregs\[9\]\[12\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold366 cpuregs\[29\]\[30\] VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 cpuregs\[31\]\[30\] VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold388 cpuregs\[12\]\[24\] VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 count_instr\[51\] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ _04271_ _04381_ _03657_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09865_ _03552_ _04314_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__or2_1
Xhold1000 cpuregs\[2\]\[27\] VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1011 cpuregs\[17\]\[11\] VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 cpuregs\[16\]\[7\] VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ reg_out\[19\] alu_out_q\[19\] _03175_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__mux2_1
Xhold1033 cpuregs\[20\]\[7\] VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ cpuregs\[8\]\[23\] cpuregs\[9\]\[23\] cpuregs\[10\]\[23\] cpuregs\[11\]\[23\]
+ _03440_ _03451_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__mux4_1
Xhold1044 is_alu_reg_reg VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1055 count_instr\[24\] VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ reg_pc\[9\] reg_pc\[8\] _03223_ reg_pc\[10\] VGND VGND VPWR VPWR _03244_
+ sky130_fd_sc_hd__a31o_1
*XANTENNA_206 net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_217 _04564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_228 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_239 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08678_ _03184_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_37_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07629_ reg_pc\[21\] decoded_imm\[21\] VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10640_ _04806_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10571_ net727 _03322_ _04768_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12310_ _03063_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__buf_4
XFILLER_0_90_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13290_ _06798_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12241_ cpuregs\[16\]\[9\] cpuregs\[17\]\[9\] cpuregs\[18\]\[9\] cpuregs\[19\]\[9\]
+ _05948_ _05925_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_79_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12172_ _05901_ _05920_ _05935_ _05904_ decoded_imm\[6\] VGND VGND VPWR VPWR _05936_
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_112_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11123_ _05094_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__buf_6
XFILLER_0_101_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15931_ clknet_leaf_132_clk _01503_ VGND VGND VPWR VPWR cpuregs\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11054_ _05043_ _05045_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__nor2_1
X_10005_ _01854_ _04427_ _04428_ _04447_ _04450_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__a311o_1
X_15862_ clknet_leaf_141_clk _01434_ VGND VGND VPWR VPWR cpuregs\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14813_ clknet_leaf_157_clk _00471_ VGND VGND VPWR VPWR cpuregs\[25\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15793_ clknet_leaf_16_clk _01368_ VGND VGND VPWR VPWR cpuregs\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14744_ clknet_leaf_152_clk _00402_ VGND VGND VPWR VPWR cpuregs\[26\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11956_ net839 _05757_ _05760_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10907_ _04963_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__clkbuf_1
X_11887_ net447 _05703_ _01905_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__o21ai_1
X_14675_ clknet_leaf_30_clk _00333_ VGND VGND VPWR VPWR cpuregs\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_104_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13626_ _03183_ _04671_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__nor2_2
X_10838_ net1272 _04825_ _04923_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_389 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10769_ _04890_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__clkbuf_1
X_13557_ _06944_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12508_ _06026_ _06257_ _06193_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13488_ _06903_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_613 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12439_ cpuregs\[28\]\[17\] cpuregs\[29\]\[17\] cpuregs\[30\]\[17\] cpuregs\[31\]\[17\]
+ _06191_ _05929_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15227_ clknet_leaf_76_clk _00820_ VGND VGND VPWR VPWR instr_bgeu sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_23_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_112_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15158_ clknet_leaf_50_clk _00783_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14109_ cpuregs\[7\]\[2\] _06929_ _01674_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__mux2_1
X_15089_ clknet_leaf_91_clk _07143_ VGND VGND VPWR VPWR reg_out\[7\] sky130_fd_sc_hd__dfxtp_1
X_07980_ _02585_ _02592_ _02597_ VGND VGND VPWR VPWR alu_out\[2\] sky130_fd_sc_hd__a21o_1
XFILLER_0_129_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09650_ cpuregs\[4\]\[18\] cpuregs\[5\]\[18\] cpuregs\[6\]\[18\] cpuregs\[7\]\[18\]
+ _03463_ _03464_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__mux4_1
X_08601_ is_slli_srli_srai decoded_imm_j\[3\] _02007_ VGND VGND VPWR VPWR _03120_
+ sky130_fd_sc_hd__a21oi_1
X_09581_ _03427_ _04035_ _04037_ _04039_ _03431_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08532_ _00008_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_121_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08463_ _02306_ _03001_ _02993_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07414_ reg_pc\[7\] decoded_imm\[7\] VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__or2_1
X_08394_ _01992_ _02953_ _02951_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_267 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_855 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_529 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07345_ net11 _01937_ _01993_ _01935_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_570 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_18_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_696 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07276_ _01926_ _01929_ _01922_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__a21oi_1
X_09015_ _00016_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_130_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold130 reg_next_pc\[25\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 instr_bge VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 count_instr\[53\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _03078_ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 reg_next_pc\[6\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 reg_sh\[1\] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 mem_rdata_q\[18\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ cpuregs\[8\]\[27\] cpuregs\[9\]\[27\] cpuregs\[10\]\[27\] cpuregs\[11\]\[27\]
+ _03582_ _03716_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_97_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_2
X_09848_ _03455_ _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__or2_1
X_09779_ cpuregs\[0\]\[22\] cpuregs\[1\]\[22\] cpuregs\[2\]\[22\] cpuregs\[3\]\[22\]
+ _03457_ _03595_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11810_ count_cycle\[25\] _05649_ count_cycle\[26\] VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _01065_ _01064_ _06518_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_1_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ count_cycle\[4\] _05601_ count_cycle\[5\] VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14460_ clknet_leaf_15_clk _00118_ VGND VGND VPWR VPWR cpuregs\[12\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11672_ _05285_ _05250_ _05546_ _05300_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10623_ _04797_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__clkbuf_1
X_13411_ _06862_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__clkbuf_1
X_14391_ clknet_leaf_8_clk _00054_ VGND VGND VPWR VPWR cpuregs\[11\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_21_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13342_ net1044 _04837_ _06816_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10554_ net985 _03268_ _04757_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13273_ _06789_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__clkbuf_1
X_10485_ cpuregs\[14\]\[13\] _03268_ _04720_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15012_ clknet_leaf_109_clk _00670_ VGND VGND VPWR VPWR reg_next_pc\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12224_ cpuregs\[16\]\[8\] cpuregs\[17\]\[8\] cpuregs\[18\]\[8\] cpuregs\[19\]\[8\]
+ _05984_ _05985_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_94_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12155_ _03106_ _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11106_ count_instr\[18\] _05082_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12086_ cpuregs\[24\]\[1\] cpuregs\[25\]\[1\] cpuregs\[26\]\[1\] cpuregs\[27\]\[1\]
+ _05834_ _03097_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_88_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_2
X_11037_ decoder_trigger VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__clkbuf_4
X_15914_ clknet_leaf_56_clk _01486_ VGND VGND VPWR VPWR cpuregs\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_160_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ clknet_leaf_35_clk _01417_ VGND VGND VPWR VPWR cpuregs\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_16 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15776_ clknet_leaf_50_clk _01351_ VGND VGND VPWR VPWR cpuregs\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12988_ _06629_ _06630_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14727_ clknet_leaf_136_clk _00385_ VGND VGND VPWR VPWR cpuregs\[15\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_11939_ _03581_ _05743_ _03547_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14658_ clknet_leaf_137_clk _00316_ VGND VGND VPWR VPWR cpuregs\[14\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13609_ cpuregs\[31\]\[26\] _06979_ _06967_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14589_ clknet_leaf_3_clk _00247_ VGND VGND VPWR VPWR cpuregs\[28\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_15_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_51_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput202 net202 VGND VGND VPWR VPWR pcpi_rs1[9] sky130_fd_sc_hd__buf_2
Xoutput213 net213 VGND VGND VPWR VPWR pcpi_rs2[19] sky130_fd_sc_hd__buf_2
Xoutput224 net224 VGND VGND VPWR VPWR pcpi_rs2[29] sky130_fd_sc_hd__buf_2
Xoutput235 net235 VGND VGND VPWR VPWR trap sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07963_ _01846_ _02503_ _02561_ _02563_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_79_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_145_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09702_ _01958_ _04144_ _04146_ _03397_ _04156_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__a32o_1
XFILLER_0_156_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07894_ _01992_ net251 VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09633_ _01870_ _04086_ _04089_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__nor3_1
X_09564_ _03766_ _03897_ _04018_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08515_ _03034_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09495_ _02154_ _03956_ _03395_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08446_ reg_next_pc\[20\] reg_out\[20\] _02969_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_136_827 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08377_ net221 _02252_ _02930_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__a21o_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07328_ net193 VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_793 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07259_ _01895_ _01896_ cpu_state\[4\] VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_234 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10270_ _04609_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13960_ _01597_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__clkbuf_1
X_12911_ _06590_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__clkbuf_1
X_13891_ _01560_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__clkbuf_1
X_15630_ clknet_leaf_1_clk _01205_ VGND VGND VPWR VPWR cpuregs\[23\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_107_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ instr_lb _06554_ _06535_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _00822_
+ sky130_fd_sc_hd__a22o_1
X_15561_ clknet_leaf_12_clk _01136_ VGND VGND VPWR VPWR cpuregs\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12773_ _01891_ _01862_ cpu_state\[6\] VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14512_ clknet_leaf_33_clk _00170_ VGND VGND VPWR VPWR cpuregs\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11724_ _05589_ _05590_ _05593_ _05367_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__a22o_1
X_15492_ clknet_leaf_94_clk _01077_ VGND VGND VPWR VPWR mem_rdata_q\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11655_ _05481_ _05499_ _05510_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__and3_1
X_14443_ clknet_leaf_56_clk _00101_ VGND VGND VPWR VPWR cpuregs\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_791 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10606_ _04788_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11586_ _05273_ _05233_ _05467_ _01902_ _01872_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__a221o_1
X_14374_ clknet_leaf_52_clk _00037_ VGND VGND VPWR VPWR cpuregs\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10537_ net1302 _03215_ _04746_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__mux2_1
X_13325_ _06817_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__clkbuf_1
X_10468_ net1390 _03215_ _04709_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__mux2_1
X_13256_ net769 _04817_ _06780_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12207_ _03045_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__buf_4
X_13187_ decoded_imm\[30\] _06740_ _06737_ _06741_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__o22a_1
X_10399_ _04678_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__clkbuf_1
X_12138_ _03080_ _05880_ _05887_ _05902_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_127_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12069_ _01906_ _05838_ _01841_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_2
X_15828_ clknet_leaf_16_clk _01400_ VGND VGND VPWR VPWR cpuregs\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_140_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15759_ clknet_leaf_5_clk _01334_ VGND VGND VPWR VPWR cpuregs\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_08300_ _02458_ _02891_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09280_ _03746_ _03747_ _03603_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_630 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_51_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08231_ net185 _02828_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08162_ _02764_ _02756_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08093_ _02657_ _02700_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ _03434_ _03445_ _03453_ _03431_ _03469_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_71_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ _01931_ _02507_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07877_ net198 net249 VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__or2_1
X_09616_ _04067_ _04069_ _04071_ _04073_ _03760_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__a221o_2
X_09547_ _02165_ _03480_ _03906_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__o21ba_1
X_09478_ _03547_ _03935_ _03937_ _03939_ _03489_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_613 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08429_ _02165_ _02977_ _02971_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11440_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11371_ decoded_imm_j\[2\] _05191_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13110_ net137 net99 _06696_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__mux2_1
X_10322_ _04637_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__clkbuf_1
X_14090_ _01666_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13041_ _06635_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__buf_4
X_10253_ net580 _03179_ _04600_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__mux2_1
X_10184_ _04563_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14992_ clknet_leaf_84_clk _00650_ VGND VGND VPWR VPWR reg_next_pc\[7\] sky130_fd_sc_hd__dfxtp_1
X_13943_ net990 _06966_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13874_ net739 _06966_ _01551_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15613_ clknet_leaf_24_clk _01188_ VGND VGND VPWR VPWR cpuregs\[31\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12825_ _06531_ _06544_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_747 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15544_ clknet_leaf_81_clk _00017_ VGND VGND VPWR VPWR cpu_state\[0\] sky130_fd_sc_hd__dfxtp_1
X_12756_ cpuregs\[28\]\[31\] cpuregs\[29\]\[31\] cpuregs\[30\]\[31\] cpuregs\[31\]\[31\]
+ _06191_ _05914_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_155_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11707_ _05418_ net497 _05358_ _05578_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15475_ clknet_leaf_95_clk _00035_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__dfxtp_1
X_12687_ cpuregs\[16\]\[28\] cpuregs\[17\]\[28\] cpuregs\[18\]\[28\] cpuregs\[19\]\[28\]
+ _05984_ _05985_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_931 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14426_ clknet_leaf_58_clk _00084_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11638_ _05273_ _05242_ _05515_ _01903_ _05184_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14357_ net920 _03347_ _01800_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_690 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11569_ decoded_imm_j\[18\] _05230_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_40_625 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold707 cpuregs\[2\]\[7\] VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13308_ net1340 _04871_ _06802_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__mux2_1
Xhold718 cpuregs\[13\]\[26\] VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold729 cpuregs\[18\]\[23\] VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ _01769_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13239_ decoded_imm\[6\] _06626_ _06769_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07800_ net179 _02416_ _02419_ net178 VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__o22a_1
XFILLER_0_137_21 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08780_ _03271_ _03272_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07731_ reg_pc\[28\] decoded_imm\[28\] VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07662_ net16 _02202_ _02179_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__a21o_1
X_09401_ _03863_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__nand2_1
X_07593_ count_instr\[50\] _02013_ _02017_ _02226_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09332_ _03796_ _03797_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_793 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09263_ reg_pc\[6\] _03527_ _03731_ _03626_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__a211o_1
XFILLER_0_157_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_35_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08214_ net215 net213 _02791_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__nor3_2
XFILLER_0_56_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09194_ _03394_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08145_ net176 _02729_ _02743_ _02177_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08076_ _02682_ _02685_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_56_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08978_ _03448_ _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__or2_1
Xhold56 mem_rdata[25] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 mem_rdata[27] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 decoded_rd\[0\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ net252 net227 VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__and2b_1
Xhold89 is_compare VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10940_ _04980_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ net1385 _04858_ _04934_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__mux2_1
X_12610_ _06177_ _06350_ _06352_ _06354_ _06164_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ _06924_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_84_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12541_ _06285_ _06287_ _06288_ _03128_ _03035_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__o221a_1
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15260_ clknet_leaf_112_clk _00853_ VGND VGND VPWR VPWR instr_rdinstrh sky130_fd_sc_hd__dfxtp_4
XFILLER_0_81_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12472_ _06132_ _06210_ _06223_ _06153_ decoded_imm\[18\] VGND VGND VPWR VPWR _06224_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_152_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14211_ _01730_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__clkbuf_1
X_11423_ _05312_ _05317_ _05288_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15191_ clknet_leaf_74_clk alu_out\[4\] VGND VGND VPWR VPWR alu_out_q\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_9 _01932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ cpuregs\[7\]\[18\] _06962_ _01685_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__mux2_1
X_11354_ _01884_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10305_ net698 _03348_ _04622_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__mux2_1
X_14073_ _01657_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__clkbuf_1
X_11285_ reg_next_pc\[9\] _03237_ _02946_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__mux2_4
X_13024_ _06649_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__clkbuf_1
X_10236_ _04591_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__clkbuf_1
X_10167_ net1035 _03348_ _04548_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__mux2_1
X_14975_ clknet_leaf_112_clk _00633_ VGND VGND VPWR VPWR reg_pc\[21\] sky130_fd_sc_hd__dfxtp_2
X_10098_ net752 _03355_ _04509_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13926_ net579 _06950_ _01577_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__mux2_1
X_13857_ net1311 _06950_ _07111_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12808_ _06528_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13788_ _07077_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_18_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_128_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15527_ clknet_leaf_152_clk _01112_ VGND VGND VPWR VPWR cpuregs\[24\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12739_ _06475_ _06477_ _06478_ _03149_ _05815_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__o221a_1
XFILLER_0_139_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15458_ clknet_leaf_157_clk _01048_ VGND VGND VPWR VPWR cpuregs\[19\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_26_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14409_ clknet_leaf_56_clk _00030_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_135_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15389_ clknet_leaf_94_clk _00979_ VGND VGND VPWR VPWR decoded_imm\[19\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_152_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold504 cpuregs\[26\]\[14\] VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold515 cpuregs\[25\]\[0\] VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold526 cpuregs\[1\]\[22\] VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 cpuregs\[10\]\[17\] VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 cpuregs\[19\]\[13\] VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 cpuregs\[12\]\[18\] VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ _04305_ _04338_ _04395_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__and3_1
X_08901_ reg_out\[30\] alu_out_q\[30\] _03176_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__mux2_1
X_09881_ _03657_ _04209_ _04328_ _04330_ _01942_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__o311a_1
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ reg_pc\[21\] _03311_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08763_ reg_pc\[11\] _03245_ reg_pc\[12\] VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07714_ _02337_ _02338_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08694_ latched_branch latched_store VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__or2b_1
X_07645_ _02260_ _02273_ _02271_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ _02194_ _02198_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09315_ _03776_ _03778_ _03781_ _03434_ _03490_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_630 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09246_ _03713_ _03714_ _03401_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09177_ _03645_ _03646_ _03647_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08128_ _02733_ _02721_ _02718_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08059_ net202 _02669_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput35 net35 VGND VGND VPWR VPWR mem_addr[10] sky130_fd_sc_hd__clkbuf_4
Xoutput46 net46 VGND VGND VPWR VPWR mem_addr[21] sky130_fd_sc_hd__buf_2
XFILLER_0_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpicorv32_290 VGND VGND VPWR VPWR picorv32_290/HI pcpi_insn[0] sky130_fd_sc_hd__conb_1
X_11070_ count_instr\[8\] _05055_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__or2_1
Xoutput57 net57 VGND VGND VPWR VPWR mem_addr[31] sky130_fd_sc_hd__buf_2
Xoutput68 net68 VGND VGND VPWR VPWR mem_la_addr[12] sky130_fd_sc_hd__clkbuf_4
Xoutput79 net79 VGND VGND VPWR VPWR mem_la_addr[23] sky130_fd_sc_hd__buf_2
X_10021_ _03500_ _04465_ _03468_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_86_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ clknet_leaf_23_clk _00418_ VGND VGND VPWR VPWR cpuregs\[26\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11972_ net569 net92 _05767_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__mux2_1
X_13711_ _07036_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__clkbuf_1
X_10923_ cpuregs\[20\]\[11\] _04842_ _04970_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14691_ clknet_leaf_127_clk _00349_ VGND VGND VPWR VPWR cpuregs\[27\]\[25\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13642_ net1145 _06939_ _06992_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__mux2_1
X_10854_ _04935_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__clkbuf_1
X_13573_ _06955_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10785_ cpuregs\[16\]\[10\] _04839_ _04898_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__mux2_1
X_15312_ clknet_leaf_6_clk _00902_ VGND VGND VPWR VPWR cpuregs\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12524_ _06142_ _06272_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15243_ clknet_leaf_78_clk _00836_ VGND VGND VPWR VPWR instr_slli sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12455_ cpuregs\[8\]\[18\] cpuregs\[9\]\[18\] cpuregs\[10\]\[18\] cpuregs\[11\]\[18\]
+ _05907_ _03039_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_117_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11406_ decoded_imm_j\[5\] _05199_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15174_ clknet_leaf_97_clk _00799_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_22_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12386_ _05879_ _06135_ _06137_ _06140_ _03104_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14125_ _01673_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11337_ _05031_ _05244_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14056_ _01648_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11268_ _05194_ reg_pc\[3\] _01843_ _05196_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13007_ _06640_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__clkbuf_1
X_10219_ _04582_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__clkbuf_1
X_11199_ _05146_ _05147_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_45 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14958_ clknet_leaf_83_clk _00616_ VGND VGND VPWR VPWR reg_pc\[4\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13909_ net1011 _06933_ _01566_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__mux2_1
X_14889_ clknet_leaf_18_clk _00547_ VGND VGND VPWR VPWR cpuregs\[17\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07430_ reg_pc\[8\] decoded_imm\[8\] VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07361_ net4 net21 _01845_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09100_ _01978_ _03572_ _03395_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__mux2_1
X_07292_ _01943_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09031_ cpuregs\[30\]\[1\] cpuregs\[31\]\[1\] _03405_ VGND VGND VPWR VPWR _03505_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold301 cpuregs\[2\]\[28\] VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_230 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold312 cpuregs\[25\]\[31\] VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 reg_next_pc\[17\] VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 cpuregs\[10\]\[20\] VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 cpuregs\[29\]\[2\] VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_641 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold356 cpuregs\[3\]\[24\] VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 cpuregs\[6\]\[30\] VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 cpuregs\[23\]\[19\] VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 cpuregs\[14\]\[30\] VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _02331_ _03617_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09864_ cpuregs\[12\]\[25\] cpuregs\[13\]\[25\] cpuregs\[14\]\[25\] cpuregs\[15\]\[25\]
+ _03808_ _03801_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__mux4_1
Xhold1001 cpuregs\[1\]\[21\] VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 cpuregs\[21\]\[8\] VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ _03303_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__clkbuf_1
Xhold1023 cpuregs\[9\]\[3\] VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 cpuregs\[22\]\[16\] VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _04245_ _04246_ _03402_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__mux2_1
Xhold1045 count_cycle\[34\] VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08746_ reg_out\[10\] alu_out_q\[10\] _03174_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__mux2_2
XFILLER_0_96_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_207 net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_218 _04846_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_229 _03547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08677_ _03180_ _03183_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_37_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ net1411 _02054_ count_cycle\[21\] _02020_ _02258_ VGND VGND VPWR VPWR _02259_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07559_ _02193_ _02194_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10570_ _04769_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09229_ _03695_ _03698_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12240_ _03143_ _06000_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12171_ _05924_ _05928_ _05931_ _05934_ _03080_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11122_ count_instr\[23\] count_instr\[22\] count_instr\[21\] _05087_ VGND VGND VPWR
+ VPWR _05094_ sky130_fd_sc_hd__and4_1
Xhold890 cpuregs\[16\]\[11\] VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__dlygate4sd3_1
X_15930_ clknet_leaf_134_clk _01502_ VGND VGND VPWR VPWR cpuregs\[0\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11053_ net608 _05039_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10004_ _03616_ _04448_ _04449_ _01942_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__o211a_1
X_15861_ clknet_leaf_3_clk _01433_ VGND VGND VPWR VPWR cpuregs\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14812_ clknet_leaf_152_clk _00470_ VGND VGND VPWR VPWR cpuregs\[25\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15792_ clknet_leaf_7_clk _01367_ VGND VGND VPWR VPWR cpuregs\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14743_ clknet_leaf_152_clk _00401_ VGND VGND VPWR VPWR cpuregs\[26\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11955_ _02007_ _05759_ _03485_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10906_ net1233 _04825_ _04959_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14674_ clknet_leaf_54_clk _00332_ VGND VGND VPWR VPWR cpuregs\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11886_ _05703_ _05704_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13625_ _06990_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10837_ _04926_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13556_ net855 _06943_ _06925_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10768_ net664 _04823_ _04887_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12507_ cpuregs\[28\]\[20\] cpuregs\[29\]\[20\] cpuregs\[30\]\[20\] cpuregs\[31\]\[20\]
+ _06191_ _05914_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13487_ net859 _04846_ _06899_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__mux2_1
X_10699_ _04843_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15226_ clknet_leaf_76_clk _00819_ VGND VGND VPWR VPWR instr_bltu sky130_fd_sc_hd__dfxtp_1
X_12438_ _03062_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_625 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15157_ clknet_leaf_50_clk _00782_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dfxtp_2
X_12369_ cpuregs\[22\]\[14\] cpuregs\[23\]\[14\] _05816_ VGND VGND VPWR VPWR _06125_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14108_ _01676_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__clkbuf_1
X_15088_ clknet_leaf_81_clk _07142_ VGND VGND VPWR VPWR reg_out\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14039_ net887 _06927_ _01638_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08600_ _03080_ _03103_ _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__a21o_2
XFILLER_0_145_21 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09580_ _03448_ _04038_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__or2_1
X_08531_ _03038_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08462_ reg_out\[24\] _02949_ _03000_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_34_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07413_ cpu_state\[3\] VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__clkbuf_4
X_08393_ reg_next_pc\[3\] reg_out\[3\] _02949_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_45_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_620 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07344_ net3 net20 _01845_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07275_ _01928_ _01887_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09014_ _03475_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold120 count_cycle\[48\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold131 count_cycle\[59\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold142 count_cycle\[34\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 net45 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 reg_next_pc\[8\] VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 count_instr\[27\] VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 count_cycle\[46\] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 instr_lbu VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09916_ _04362_ _04363_ _03401_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__mux2_1
X_09847_ cpuregs\[28\]\[24\] cpuregs\[29\]\[24\] cpuregs\[30\]\[24\] cpuregs\[31\]\[24\]
+ _03641_ _03642_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__mux4_1
X_09778_ cpuregs\[4\]\[22\] cpuregs\[5\]\[22\] cpuregs\[6\]\[22\] cpuregs\[7\]\[22\]
+ _03457_ _03595_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__mux4_1
X_08729_ net731 _03228_ _03185_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ count_cycle\[4\] count_cycle\[5\] _05601_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__and3_1
X_11671_ _05541_ _05542_ _05545_ _05289_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13410_ net1179 _04837_ _06852_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10622_ cpuregs\[15\]\[13\] _03268_ _04793_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__mux2_1
X_14390_ clknet_leaf_12_clk _00053_ VGND VGND VPWR VPWR cpuregs\[11\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13341_ _06825_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__clkbuf_1
X_10553_ _04760_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_399 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_107_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_358 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13272_ net639 _04835_ _06780_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10484_ _04723_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_20_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15011_ clknet_leaf_109_clk _00669_ VGND VGND VPWR VPWR reg_next_pc\[26\] sky130_fd_sc_hd__dfxtp_1
X_12223_ _03052_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_94_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12154_ cpuregs\[8\]\[6\] cpuregs\[9\]\[6\] cpuregs\[10\]\[6\] cpuregs\[11\]\[6\]
+ _03150_ _05917_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__mux4_1
X_11105_ _05080_ _05078_ _05082_ _05052_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_9_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12085_ _03082_ _05853_ _03034_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__o21ai_1
X_11036_ _01891_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__clkbuf_4
X_15913_ clknet_leaf_34_clk _01485_ VGND VGND VPWR VPWR cpuregs\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15844_ clknet_leaf_26_clk _01416_ VGND VGND VPWR VPWR cpuregs\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_160_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ clknet_leaf_50_clk _01350_ VGND VGND VPWR VPWR cpuregs\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12987_ _01066_ _01068_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__nor2_1
X_14726_ clknet_leaf_137_clk _00384_ VGND VGND VPWR VPWR cpuregs\[15\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11938_ cpuregs\[16\]\[31\] cpuregs\[17\]\[31\] cpuregs\[18\]\[31\] cpuregs\[19\]\[31\]
+ _03598_ _03460_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14657_ clknet_leaf_137_clk _00315_ VGND VGND VPWR VPWR cpuregs\[14\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11869_ _05036_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_642 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13608_ _03354_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14588_ clknet_leaf_154_clk _00246_ VGND VGND VPWR VPWR cpuregs\[28\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13539_ _06932_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15209_ clknet_leaf_101_clk alu_out\[22\] VGND VGND VPWR VPWR alu_out_q\[22\] sky130_fd_sc_hd__dfxtp_1
Xoutput203 net203 VGND VGND VPWR VPWR pcpi_rs2[0] sky130_fd_sc_hd__buf_2
XFILLER_0_101_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput214 net214 VGND VGND VPWR VPWR pcpi_rs2[1] sky130_fd_sc_hd__buf_2
Xoutput225 net225 VGND VGND VPWR VPWR pcpi_rs2[2] sky130_fd_sc_hd__buf_2
XFILLER_0_2_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07962_ _02568_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_145_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ _04152_ _04155_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__xor2_1
XFILLER_0_156_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07893_ _01930_ _02503_ _02510_ _02512_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__a31o_1
X_09632_ _04026_ _04087_ _04088_ _04053_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_78_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09563_ _03900_ _04018_ _04019_ _04021_ _04011_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__o2111a_1
X_08514_ _00010_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__clkinv_4
X_09494_ _03651_ _03931_ _03932_ _03951_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__a311o_1
XFILLER_0_77_255 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_78_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08445_ _02988_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_1
XFILLER_0_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08376_ net220 _02927_ _02929_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__a21o_1
XFILLER_0_73_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07327_ _01958_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07258_ net652 _01874_ _01876_ _01913_ _01914_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07189_ _01853_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__buf_4
XFILLER_0_112_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12910_ mem_rdata_q\[25\] net18 _06589_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__mux2_1
X_13890_ net828 _06983_ _01551_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_509 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_159_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12841_ _06553_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15560_ clknet_leaf_11_clk _01135_ VGND VGND VPWR VPWR cpuregs\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12772_ _03032_ _06507_ _01885_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14511_ clknet_leaf_39_clk _00169_ VGND VGND VPWR VPWR cpuregs\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11723_ _05591_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15491_ clknet_leaf_86_clk _01076_ VGND VGND VPWR VPWR mem_rdata_q\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ clknet_leaf_52_clk _00100_ VGND VGND VPWR VPWR cpuregs\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11654_ _05494_ _05529_ _05508_ _05507_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10605_ cpuregs\[15\]\[5\] _03215_ _04782_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14373_ _05358_ net1397 _01813_ _01814_ _05767_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__a41o_1
XFILLER_0_51_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11585_ _05233_ _05457_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13324_ net982 _04817_ _06816_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__mux2_1
X_10536_ _04751_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__clkbuf_1
X_13255_ _06779_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_566 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10467_ _04714_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12206_ _03142_ _05963_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__or3_1
X_13186_ mem_rdata_q\[30\] _06738_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__and2_1
X_10398_ cpuregs\[21\]\[4\] _03209_ _04673_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__mux2_1
X_12137_ _03104_ _05893_ _05899_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__o31a_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12068_ _03104_ _05826_ _05837_ _03058_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__o211ai_4
X_11019_ _05022_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__clkbuf_1
X_15827_ clknet_leaf_7_clk _01399_ VGND VGND VPWR VPWR cpuregs\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_140_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_907 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15758_ clknet_leaf_8_clk _01333_ VGND VGND VPWR VPWR cpuregs\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_564 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14709_ clknet_leaf_10_clk _00367_ VGND VGND VPWR VPWR cpuregs\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15689_ clknet_leaf_8_clk _01264_ VGND VGND VPWR VPWR cpuregs\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08230_ net217 _02827_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08161_ _02756_ _02764_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__or2b_1
XFILLER_0_71_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08092_ net205 net248 net234 net233 VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_892 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08994_ _03455_ _03462_ _03466_ _03468_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_54_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07945_ _01847_ _02507_ _02561_ _02564_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_3_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07876_ net198 net249 VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__nand2_1
X_09615_ _03414_ _04072_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__or2_1
X_09546_ _03473_ _03996_ _04005_ _03526_ reg_pc\[15\] VGND VGND VPWR VPWR _04006_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_918 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09477_ _03807_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_940 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08428_ reg_next_pc\[14\] reg_out\[14\] _02969_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08359_ _02507_ net247 _02251_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_883 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11370_ _05264_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10321_ cpuregs\[28\]\[0\] _03179_ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13040_ _06657_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__clkbuf_1
X_10252_ _04599_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__buf_6
X_10183_ _04481_ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_109_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14991_ clknet_leaf_84_clk _00649_ VGND VGND VPWR VPWR reg_next_pc\[6\] sky130_fd_sc_hd__dfxtp_1
X_13942_ _01565_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13873_ _07099_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_122_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15612_ clknet_leaf_132_clk _01187_ VGND VGND VPWR VPWR cpuregs\[31\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12824_ _06532_ _06536_ _06533_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15543_ clknet_leaf_64_clk _00006_ VGND VGND VPWR VPWR reg_sh\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _03132_ _06493_ _05840_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11706_ _05193_ _05577_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15474_ clknet_leaf_97_clk _00034_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__dfxtp_2
X_12686_ _06142_ _06427_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_127_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14425_ clknet_leaf_60_clk _00083_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_127_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11637_ _05242_ _05503_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14356_ _01805_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__clkbuf_1
X_11568_ _05263_ net682 _05358_ _05450_ _05451_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_80_784 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13307_ _06807_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__clkbuf_1
Xhold708 cpuregs\[10\]\[24\] VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold719 cpuregs\[26\]\[27\] VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ _04741_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__clkbuf_1
X_14287_ net530 VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11499_ _05367_ _05387_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__nor2_1
X_13238_ _06763_ decoded_imm_j\[6\] _06733_ mem_rdata_q\[26\] _06541_ VGND VGND VPWR
+ VPWR _06769_ sky130_fd_sc_hd__a221o_1
X_13169_ is_slli_srli_srai _05838_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_33 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07730_ reg_pc\[28\] decoded_imm\[28\] VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__or2_1
X_07661_ net186 VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__clkbuf_8
X_09400_ decoded_imm\[11\] net173 VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07592_ count_instr\[18\] _01949_ count_cycle\[50\] _01947_ VGND VGND VPWR VPWR _02226_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_203 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09331_ decoded_imm\[8\] _02082_ _03767_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09262_ _03473_ _03722_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__and3_2
XFILLER_0_157_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08213_ _02584_ _02809_ _02810_ _02812_ _02405_ VGND VGND VPWR VPWR alu_out\[20\]
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09193_ _03651_ _03655_ _03656_ _03663_ _03488_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__a311o_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08144_ _02469_ _02741_ _02748_ _02585_ VGND VGND VPWR VPWR alu_out\[15\] sky130_fd_sc_hd__a22o_1
XFILLER_0_160_436 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08075_ _02671_ _02683_ _02684_ _02666_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08977_ cpuregs\[20\]\[0\] cpuregs\[21\]\[0\] cpuregs\[22\]\[0\] cpuregs\[23\]\[0\]
+ _03440_ _03451_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__mux4_1
Xhold57 mem_rdata[18] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _02488_ _02501_ _02541_ _02547_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__nor4b_1
Xhold68 decoded_rd\[2\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 instr_auipc VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ _02112_ net248 VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10870_ _04943_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_715 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09529_ cpuregs\[4\]\[15\] cpuregs\[5\]\[15\] cpuregs\[6\]\[15\] cpuregs\[7\]\[15\]
+ _03439_ _03576_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12540_ cpuregs\[0\]\[22\] cpuregs\[1\]\[22\] cpuregs\[2\]\[22\] cpuregs\[3\]\[22\]
+ _05819_ _03125_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_271 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_770 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12471_ _05886_ _06212_ _06216_ _05978_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__a311o_2
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14210_ cpuregs\[8\]\[18\] _06962_ _01721_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11422_ _05315_ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__xor2_1
X_15190_ clknet_leaf_73_clk alu_out\[3\] VGND VGND VPWR VPWR alu_out_q\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14141_ _01693_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__clkbuf_1
X_11353_ _05231_ reg_pc\[29\] VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_89_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10304_ _04627_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__clkbuf_1
X_14072_ net1368 _06960_ _01649_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__mux2_1
X_11284_ _05194_ reg_pc\[8\] _01843_ _05207_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__o211a_1
X_13023_ cpuregs\[1\]\[11\] _04842_ _06647_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__mux2_1
X_10235_ net1055 _03341_ _04586_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_889 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_100_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10166_ _04553_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__clkbuf_1
X_14974_ clknet_leaf_106_clk _00632_ VGND VGND VPWR VPWR reg_pc\[20\] sky130_fd_sc_hd__dfxtp_2
X_10097_ _04515_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__clkbuf_1
X_13925_ _01579_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_98_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13856_ _07113_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12807_ _06529_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13787_ net1025 _06948_ _07075_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__mux2_1
X_10999_ cpuregs\[17\]\[15\] _04850_ _05006_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15526_ clknet_leaf_159_clk _01111_ VGND VGND VPWR VPWR cpuregs\[24\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12738_ cpuregs\[16\]\[30\] cpuregs\[17\]\[30\] cpuregs\[18\]\[30\] cpuregs\[19\]\[30\]
+ _05921_ _05922_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_26_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15457_ clknet_leaf_159_clk _01047_ VGND VGND VPWR VPWR cpuregs\[19\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12669_ cpuregs\[22\]\[27\] cpuregs\[23\]\[27\] _05979_ VGND VGND VPWR VPWR _06412_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_155_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14408_ clknet_leaf_57_clk _00029_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15388_ clknet_leaf_94_clk _00978_ VGND VGND VPWR VPWR decoded_imm\[20\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_924 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14339_ _01796_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold505 cpuregs\[10\]\[1\] VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 cpuregs\[25\]\[18\] VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold527 cpuregs\[28\]\[6\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 cpuregs\[4\]\[0\] VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 cpuregs\[21\]\[18\] VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__dlygate4sd3_1
X_08900_ reg_pc\[30\] _03371_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09880_ _04211_ _04329_ _03657_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_51_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ reg_out\[21\] alu_out_q\[21\] _03175_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08762_ reg_out\[12\] alu_out_q\[12\] _03174_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__mux2_1
X_07713_ _02327_ _02329_ _02326_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__a21o_1
X_08693_ reg_pc\[3\] _01971_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07644_ _02260_ _02271_ _02273_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07575_ _02208_ _02209_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09314_ _03779_ _03780_ _03455_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_91_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09245_ cpuregs\[16\]\[6\] cpuregs\[17\]\[6\] cpuregs\[18\]\[6\] cpuregs\[19\]\[6\]
+ _03404_ _03408_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09176_ _03579_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__buf_6
XFILLER_0_160_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08127_ net175 _02717_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_98_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08058_ _02482_ _02668_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput36 net36 VGND VGND VPWR VPWR mem_addr[11] sky130_fd_sc_hd__clkbuf_4
Xoutput47 net47 VGND VGND VPWR VPWR mem_addr[22] sky130_fd_sc_hd__buf_2
XFILLER_0_12_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput58 net58 VGND VGND VPWR VPWR mem_addr[3] sky130_fd_sc_hd__clkbuf_4
Xpicorv32_280 VGND VGND VPWR VPWR picorv32_280/HI eoi[26] sky130_fd_sc_hd__conb_1
Xpicorv32_291 VGND VGND VPWR VPWR picorv32_291/HI pcpi_insn[1] sky130_fd_sc_hd__conb_1
Xoutput69 net69 VGND VGND VPWR VPWR mem_la_addr[13] sky130_fd_sc_hd__clkbuf_4
X_10020_ cpuregs\[24\]\[30\] cpuregs\[25\]\[30\] cpuregs\[26\]\[30\] cpuregs\[27\]\[30\]
+ _03458_ _03637_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _05771_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__clkbuf_1
X_13710_ net627 _06939_ _07028_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__mux2_1
X_10922_ _04971_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__clkbuf_1
X_14690_ clknet_leaf_127_clk _00348_ VGND VGND VPWR VPWR cpuregs\[27\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13641_ _06999_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__clkbuf_1
X_10853_ cpuregs\[25\]\[10\] _04839_ _04934_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_539 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13572_ net640 _06954_ _06946_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__mux2_1
X_10784_ _04886_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__buf_4
XFILLER_0_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15311_ clknet_leaf_8_clk _00901_ VGND VGND VPWR VPWR cpuregs\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12523_ cpuregs\[20\]\[21\] cpuregs\[21\]\[21\] cpuregs\[22\]\[21\] cpuregs\[23\]\[21\]
+ _06065_ _03144_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_125_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15242_ clknet_leaf_77_clk _00835_ VGND VGND VPWR VPWR instr_sw sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12454_ cpuregs\[12\]\[18\] cpuregs\[13\]\[18\] cpuregs\[14\]\[18\] cpuregs\[15\]\[18\]
+ _05834_ _03129_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_117_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11405_ _05258_ net1027 _05239_ _05301_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__o211a_1
X_15173_ clknet_leaf_96_clk _00798_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dfxtp_1
X_12385_ _06138_ _06139_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14124_ _01684_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_97_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_607 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11336_ _02947_ _03336_ _03000_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_104_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14055_ cpuregs\[6\]\[9\] _06943_ _01638_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__mux2_1
X_11267_ _01872_ _05195_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__or2_1
X_13006_ net792 _04825_ _06636_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__mux2_1
X_10218_ cpuregs\[13\]\[16\] _03287_ _04575_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__mux2_1
X_11198_ net554 _05143_ _05133_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10149_ _04544_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14957_ clknet_leaf_83_clk _00615_ VGND VGND VPWR VPWR reg_pc\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13908_ _01570_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__clkbuf_1
X_14888_ clknet_leaf_23_clk _00546_ VGND VGND VPWR VPWR cpuregs\[17\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13839_ _07104_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07360_ net197 VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15509_ clknet_leaf_54_clk _01094_ VGND VGND VPWR VPWR cpuregs\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_07291_ _01942_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09030_ cpuregs\[28\]\[1\] cpuregs\[29\]\[1\] _03406_ VGND VGND VPWR VPWR _03504_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_795 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_130_406 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold302 cpuregs\[15\]\[12\] VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold313 instr_sw VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 cpuregs\[15\]\[17\] VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold335 cpuregs\[27\]\[30\] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 cpuregs\[11\]\[26\] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 cpuregs\[24\]\[1\] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 cpuregs\[27\]\[21\] VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net252 _03617_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold379 cpuregs\[22\]\[19\] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09863_ _03557_ _04312_ _03417_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__o21a_1
X_08814_ net984 _03302_ _03249_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__mux2_1
Xhold1002 reg_next_pc\[28\] VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 cpuregs\[19\]\[23\] VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ cpuregs\[0\]\[23\] cpuregs\[1\]\[23\] cpuregs\[2\]\[23\] cpuregs\[3\]\[23\]
+ _03405_ _03496_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__mux4_1
Xhold1024 cpuregs\[14\]\[0\] VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 cpuregs\[21\]\[3\] VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 reg_sh\[2\] VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _03242_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_208 net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_219 _04846_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08676_ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ count_instr\[53\] _02052_ _02014_ count_cycle\[53\] VGND VGND VPWR VPWR _02258_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ reg_pc\[16\] decoded_imm\[16\] VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07489_ count_instr\[11\] _01965_ count_cycle\[11\] _01951_ _02129_ VGND VGND VPWR
+ VPWR _02130_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09228_ _03696_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09159_ _03437_ _03629_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12170_ _03149_ _05933_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11121_ _05092_ _05093_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold880 cpuregs\[5\]\[8\] VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 cpuregs\[31\]\[31\] VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ _05040_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_196 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10003_ _04335_ _04392_ _03482_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__o21ai_1
X_15860_ clknet_leaf_16_clk _01432_ VGND VGND VPWR VPWR cpuregs\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14811_ clknet_leaf_160_clk _00469_ VGND VGND VPWR VPWR cpuregs\[25\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15791_ clknet_leaf_5_clk _01366_ VGND VGND VPWR VPWR cpuregs\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14742_ clknet_leaf_156_clk _00400_ VGND VGND VPWR VPWR cpuregs\[26\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11954_ _03483_ _05758_ _03390_ _01897_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10905_ _04962_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__clkbuf_1
X_14673_ clknet_leaf_36_clk _00331_ VGND VGND VPWR VPWR cpuregs\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11885_ count_cycle\[50\] _05700_ _05647_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_15_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13624_ net1250 _06989_ _06924_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__mux2_1
X_10836_ cpuregs\[25\]\[2\] _04823_ _04923_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_82_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13555_ _03240_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_17_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_857 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10767_ _04889_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12506_ _06023_ _06255_ _05840_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__o21a_1
X_13486_ _06902_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10698_ cpuregs\[26\]\[11\] _04842_ _04840_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15225_ clknet_leaf_80_clk _00818_ VGND VGND VPWR VPWR instr_bge sky130_fd_sc_hd__dfxtp_1
X_12437_ _06023_ _06189_ _05927_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15156_ clknet_leaf_49_clk _00781_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_1
X_12368_ _05872_ _06123_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__and2_1
X_14107_ cpuregs\[7\]\[1\] _06927_ _01674_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11319_ _05227_ _05230_ _05232_ _05224_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__o211a_1
X_15087_ clknet_leaf_81_clk _07141_ VGND VGND VPWR VPWR reg_out\[5\] sky130_fd_sc_hd__dfxtp_1
X_12299_ _06054_ _06056_ _06014_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14038_ _01639_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_26_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_33 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08530_ _03036_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08461_ reg_next_pc\[24\] _02999_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07412_ count_cycle\[7\] _02051_ _02053_ _02056_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__a211o_2
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08392_ _02952_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_1
XFILLER_0_18_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07343_ net196 VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07274_ _01927_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_531 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09013_ _01847_ _03396_ _03478_ _03487_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_732 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_85_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold110 instr_bgeu VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 count_instr\[25\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 instr_slti VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 count_cycle\[31\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 count_instr\[44\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 cpuregs\[0\]\[0\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 count_instr\[40\] VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 count_instr\[62\] VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold198 instr_sltiu VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ cpuregs\[0\]\[27\] cpuregs\[1\]\[27\] cpuregs\[2\]\[27\] cpuregs\[3\]\[27\]
+ _03439_ _03576_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__mux4_1
X_09846_ _03415_ _04296_ _03420_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__o21a_1
X_09777_ _03746_ _04229_ _03467_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08728_ _03227_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08659_ mem_rdata_q\[24\] net17 _03017_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__mux2_1
X_11670_ _05543_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10621_ _04796_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_37_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13340_ net1303 _04835_ _06816_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__mux2_1
X_10552_ net667 _03263_ _04757_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13271_ _06788_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10483_ net603 _03263_ _04720_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15010_ clknet_leaf_109_clk _00668_ VGND VGND VPWR VPWR reg_next_pc\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12222_ _03051_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__buf_6
XFILLER_0_121_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12153_ _03052_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11104_ count_instr\[15\] count_instr\[14\] _05072_ _05081_ VGND VGND VPWR VPWR _05082_
+ sky130_fd_sc_hd__and4_4
X_12084_ cpuregs\[20\]\[1\] cpuregs\[21\]\[1\] cpuregs\[22\]\[1\] cpuregs\[23\]\[1\]
+ _05816_ _03086_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_9_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15912_ clknet_leaf_32_clk _01484_ VGND VGND VPWR VPWR cpuregs\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11035_ _05030_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__clkbuf_1
X_15843_ clknet_leaf_50_clk _01415_ VGND VGND VPWR VPWR cpuregs\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ clknet_leaf_22_clk _01349_ VGND VGND VPWR VPWR cpuregs\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12986_ _01065_ _01064_ _06518_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__nor3b_2
XTAP_TAPCELL_ROW_125_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ clknet_leaf_21_clk _00383_ VGND VGND VPWR VPWR cpuregs\[15\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11937_ _03593_ _05741_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11868_ count_cycle\[43\] net473 count_cycle\[45\] _05686_ VGND VGND VPWR VPWR _05692_
+ sky130_fd_sc_hd__and4_4
X_14656_ clknet_leaf_138_clk _00314_ VGND VGND VPWR VPWR cpuregs\[14\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13607_ _06978_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__clkbuf_1
X_10819_ _04916_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14587_ clknet_leaf_2_clk _00245_ VGND VGND VPWR VPWR cpuregs\[28\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_11799_ _05645_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13538_ cpuregs\[31\]\[3\] _06931_ _06925_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13469_ _06893_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_401 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15208_ clknet_leaf_102_clk alu_out\[21\] VGND VGND VPWR VPWR alu_out_q\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_445 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput204 net204 VGND VGND VPWR VPWR pcpi_rs2[10] sky130_fd_sc_hd__buf_2
Xoutput215 net215 VGND VGND VPWR VPWR pcpi_rs2[20] sky130_fd_sc_hd__buf_2
Xoutput226 net226 VGND VGND VPWR VPWR pcpi_rs2[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15139_ clknet_leaf_110_clk _00765_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfxtp_1
X_07961_ _02566_ _02578_ net1416 VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__o21a_1
X_09700_ _04153_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07892_ _01978_ _02509_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09631_ _04085_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__inv_2
X_09562_ _03963_ _04012_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08513_ _00011_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__inv_4
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09493_ _03657_ _03839_ _03952_ _03954_ _01942_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_156_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_156_clk sky130_fd_sc_hd__clkbuf_2
X_08444_ _02237_ _02987_ _02971_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_46_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ net246 _02927_ _02928_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__a21o_1
XFILLER_0_46_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07326_ _01972_ _01975_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_564 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07257_ net529 instr_lh _01866_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_52_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07188_ cpu_state\[6\] cpu_state\[5\] VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_76_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ _04149_ _04276_ _04279_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__o21ai_1
X_12840_ _06540_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_61_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _01893_ _05193_ _05269_ _06506_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_147_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_147_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_139_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11722_ _05495_ _05261_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__xnor2_1
X_14510_ clknet_leaf_44_clk _00168_ VGND VGND VPWR VPWR cpuregs\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15490_ clknet_leaf_86_clk _01075_ VGND VGND VPWR VPWR mem_rdata_q\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _05244_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14441_ clknet_leaf_65_clk _00099_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_139_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10604_ _04787_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14372_ net420 net235 VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__nand2_1
X_11584_ _05463_ _05465_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13323_ _06815_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_122_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10535_ net1140 _03209_ _04746_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_70_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13254_ _04524_ _04885_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__nor2_4
X_10466_ net1100 _03209_ _04709_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12205_ _05845_ _05964_ _05966_ _03139_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13185_ _06531_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__buf_2
X_10397_ _04677_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__clkbuf_1
X_12136_ _05900_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__buf_4
X_12067_ _05828_ _05831_ _05833_ _05836_ _03033_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_127_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11018_ cpuregs\[17\]\[24\] _04869_ _05017_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__mux2_1
X_15826_ clknet_leaf_6_clk _01398_ VGND VGND VPWR VPWR cpuregs\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15757_ clknet_leaf_142_clk _01332_ VGND VGND VPWR VPWR cpuregs\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_138_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_138_clk sky130_fd_sc_hd__clkbuf_2
X_12969_ _06619_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14708_ clknet_leaf_10_clk _00366_ VGND VGND VPWR VPWR cpuregs\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15688_ clknet_leaf_32_clk _01263_ VGND VGND VPWR VPWR cpuregs\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14639_ clknet_leaf_39_clk _00297_ VGND VGND VPWR VPWR cpuregs\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08160_ _02762_ _02763_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_659 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08091_ _02485_ _02691_ _02698_ _02699_ VGND VGND VPWR VPWR alu_out\[11\] sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08993_ _03467_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_118_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07944_ _01847_ _02507_ _02563_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_71_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07875_ _02493_ _02494_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__and2_1
X_09614_ cpuregs\[24\]\[17\] cpuregs\[25\]\[17\] cpuregs\[26\]\[17\] cpuregs\[27\]\[17\]
+ _03516_ _03409_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09545_ _03998_ _04000_ _04002_ _04004_ _03430_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__a221o_2
Xclkbuf_leaf_129_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_129_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_149_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09476_ cpuregs\[12\]\[13\] cpuregs\[13\]\[13\] cpuregs\[14\]\[13\] cpuregs\[15\]\[13\]
+ _03808_ _03801_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08427_ _02976_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_102_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08358_ net209 _02927_ _02935_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__a21o_1
XFILLER_0_74_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07309_ net9 _01937_ _01959_ _01935_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_292 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08289_ _02757_ _02881_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10320_ _04635_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10251_ _04483_ _04524_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__nor2_2
X_10182_ _04561_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout250 net123 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__buf_2
X_14990_ clknet_leaf_84_clk _00648_ VGND VGND VPWR VPWR reg_next_pc\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13941_ _01587_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13872_ _01550_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15611_ clknet_leaf_129_clk _01186_ VGND VGND VPWR VPWR cpuregs\[31\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12823_ _05358_ _06542_ _06543_ _06530_ net474 VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_159_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ clknet_leaf_72_clk _00005_ VGND VGND VPWR VPWR reg_sh\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12754_ cpuregs\[16\]\[31\] cpuregs\[17\]\[31\] cpuregs\[18\]\[31\] cpuregs\[19\]\[31\]
+ _05984_ _05985_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11705_ _01903_ _05569_ _05575_ _05264_ _05576_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_401 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12685_ cpuregs\[20\]\[28\] cpuregs\[21\]\[28\] cpuregs\[22\]\[28\] cpuregs\[23\]\[28\]
+ _03095_ _03144_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__mux4_1
X_15473_ clknet_leaf_99_clk _00033_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11636_ _05269_ _05511_ _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__and3_1
X_14424_ clknet_leaf_57_clk _00082_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14355_ net1067 _03340_ _01800_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__mux2_1
X_11567_ _05300_ _05431_ _05228_ _05184_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13306_ net964 _04869_ _06802_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__mux2_1
X_10518_ net821 _03374_ _04731_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__mux2_1
Xhold709 cpuregs\[30\]\[23\] VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__dlygate4sd3_1
X_14286_ _01768_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11498_ _05215_ _05380_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13237_ decoded_imm\[7\] _06626_ _06768_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__o21a_1
X_10449_ _04704_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_150_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13168_ net434 _03670_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__or2_1
X_12119_ cpuregs\[28\]\[5\] cpuregs\[29\]\[5\] _03096_ VGND VGND VPWR VPWR _05884_
+ sky130_fd_sc_hd__mux2_1
X_13099_ net163 _02492_ _06685_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07660_ _02287_ _02288_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__xor2_1
X_15809_ clknet_leaf_73_clk _00026_ VGND VGND VPWR VPWR mem_wordsize\[2\] sky130_fd_sc_hd__dfxtp_2
X_07591_ _01970_ _02221_ _02224_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09330_ _03794_ _03795_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09261_ _03724_ _03726_ _03729_ _03426_ _03489_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08212_ _02595_ _02811_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09192_ _03657_ _03658_ _03661_ _03662_ _01953_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__o221a_1
XFILLER_0_161_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08143_ _02746_ _02747_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_454 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_448 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_487 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_125_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08074_ _02662_ _02670_ _02671_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08976_ _03450_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__clkbuf_8
Xhold58 mem_rdata[11] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _02546_ _02510_ _02508_ _02506_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__and4b_1
Xhold69 mem_rdata[8] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
X_07858_ _02082_ _02476_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_27_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07789_ net213 VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09528_ _02165_ _03624_ _03988_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09459_ cpuregs\[0\]\[12\] cpuregs\[1\]\[12\] cpuregs\[2\]\[12\] cpuregs\[3\]\[12\]
+ _03457_ _03595_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_283 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_207 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12470_ _06218_ _06220_ _06221_ _03132_ _05815_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11421_ _05304_ _05305_ _05303_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14140_ net1116 _06960_ _01685_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11352_ reg_next_pc\[29\] _03369_ _02948_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__mux2_2
X_10303_ net1347 _03341_ _04622_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14071_ _01656_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__clkbuf_1
X_11283_ _01872_ _05206_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_115_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13022_ _06648_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__clkbuf_1
X_10234_ _04590_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__clkbuf_1
X_10165_ net838 _03341_ _04548_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__mux2_1
X_14973_ clknet_leaf_106_clk _00631_ VGND VGND VPWR VPWR reg_pc\[19\] sky130_fd_sc_hd__dfxtp_2
X_10096_ net1214 _03348_ _04509_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__mux2_1
X_13924_ cpuregs\[4\]\[11\] _06948_ _01577_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__mux2_1
X_13855_ cpuregs\[22\]\[11\] _06948_ _07111_ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__mux2_1
X_12806_ _01820_ _06528_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__nor2_2
X_10998_ _05011_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__clkbuf_1
X_13786_ _07076_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15525_ clknet_leaf_156_clk _01110_ VGND VGND VPWR VPWR cpuregs\[24\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_710 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_84_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12737_ _05896_ _06476_ _03153_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_139_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_760 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15456_ clknet_leaf_159_clk _01046_ VGND VGND VPWR VPWR cpuregs\[19\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12668_ _05872_ _06410_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ clknet_leaf_57_clk _00028_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__dfxtp_2
X_11619_ decoded_imm_j\[20\] _05240_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15387_ clknet_leaf_94_clk _00977_ VGND VGND VPWR VPWR decoded_imm\[21\] sky130_fd_sc_hd__dfxtp_2
X_12599_ _06338_ _06340_ _06342_ _06344_ _06151_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_41_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_104 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_41_936 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14338_ net924 _03286_ _01789_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold506 cpuregs\[9\]\[27\] VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 cpuregs\[28\]\[1\] VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap236 _02844_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
Xhold528 cpuregs\[6\]\[1\] VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 cpuregs\[22\]\[23\] VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ net486 VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _03316_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08761_ _03256_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__clkbuf_1
X_07712_ _02335_ _02336_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__nand2_1
X_08692_ reg_out\[3\] alu_out_q\[3\] latched_stalu VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__mux2_1
X_07643_ _02247_ _02272_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07574_ reg_pc\[17\] decoded_imm\[17\] VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_822 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09313_ cpuregs\[0\]\[8\] cpuregs\[1\]\[8\] cpuregs\[2\]\[8\] cpuregs\[3\]\[8\] _03641_
+ _03642_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_60_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_2
X_09244_ cpuregs\[20\]\[6\] cpuregs\[21\]\[6\] cpuregs\[22\]\[6\] cpuregs\[23\]\[6\]
+ _03404_ _03576_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_63_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09175_ cpuregs\[16\]\[4\] cpuregs\[17\]\[4\] cpuregs\[18\]\[4\] cpuregs\[19\]\[4\]
+ _03458_ _03461_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08126_ _02730_ _02731_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08057_ _02476_ _02657_ _02656_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput37 net37 VGND VGND VPWR VPWR mem_addr[12] sky130_fd_sc_hd__clkbuf_4
Xpicorv32_270 VGND VGND VPWR VPWR picorv32_270/HI eoi[16] sky130_fd_sc_hd__conb_1
Xoutput48 net48 VGND VGND VPWR VPWR mem_addr[23] sky130_fd_sc_hd__clkbuf_4
Xpicorv32_281 VGND VGND VPWR VPWR picorv32_281/HI eoi[27] sky130_fd_sc_hd__conb_1
Xoutput59 net59 VGND VGND VPWR VPWR mem_addr[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpicorv32_292 VGND VGND VPWR VPWR picorv32_292/HI pcpi_insn[2] sky130_fd_sc_hd__conb_1
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08959_ _03433_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_86_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11970_ net60 net91 _05767_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10921_ cpuregs\[20\]\[10\] _04839_ _04970_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10852_ _04922_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__buf_4
X_13640_ net1049 _06937_ _06992_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _03274_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__buf_2
XFILLER_0_67_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10783_ _04897_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_51_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_2
X_15310_ clknet_leaf_142_clk _00900_ VGND VGND VPWR VPWR cpuregs\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12522_ _06177_ _06266_ _06268_ _06270_ _06164_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15241_ clknet_leaf_76_clk _00834_ VGND VGND VPWR VPWR instr_andi sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12453_ _06201_ _06203_ _06204_ _03128_ _03035_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_10_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11404_ _05285_ _05198_ _05299_ _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__a22o_1
X_12384_ cpuregs\[8\]\[15\] cpuregs\[9\]\[15\] cpuregs\[10\]\[15\] cpuregs\[11\]\[15\]
+ _06061_ _05917_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__mux4_1
X_15172_ clknet_leaf_61_clk _00797_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11335_ _05227_ _05242_ _05243_ _05224_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__o211a_1
X_14123_ net1274 _06943_ _01674_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_619 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14054_ _01647_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__clkbuf_1
X_11266_ reg_next_pc\[3\] _03196_ _02945_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__mux2_2
X_10217_ _04581_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__clkbuf_1
X_13005_ _06639_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__clkbuf_1
X_11197_ count_instr\[46\] count_instr\[45\] net513 _05139_ VGND VGND VPWR VPWR _05146_
+ sky130_fd_sc_hd__and4_1
X_10148_ net1193 _03287_ _04537_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__mux2_1
X_10079_ cpuregs\[12\]\[17\] _03295_ _04498_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__mux2_1
X_14956_ clknet_leaf_92_clk _00614_ VGND VGND VPWR VPWR reg_pc\[2\] sky130_fd_sc_hd__dfxtp_1
X_13907_ net566 _06931_ _01566_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__mux2_1
X_14887_ clknet_leaf_125_clk _00545_ VGND VGND VPWR VPWR cpuregs\[17\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13838_ cpuregs\[22\]\[3\] _06931_ _07100_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13769_ _07067_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_2
X_15508_ clknet_leaf_88_clk _01093_ VGND VGND VPWR VPWR mem_rdata_q\[31\] sky130_fd_sc_hd__dfxtp_2
X_07290_ cpu_state\[4\] VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15439_ clknet_leaf_18_clk _01029_ VGND VGND VPWR VPWR cpuregs\[18\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_41_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold303 cpuregs\[16\]\[1\] VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold314 instr_sb VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__buf_1
XFILLER_0_142_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold325 cpuregs\[15\]\[22\] VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold336 cpuregs\[31\]\[27\] VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 cpuregs\[23\]\[24\] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold358 cpuregs\[26\]\[12\] VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 cpuregs\[9\]\[29\] VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _03473_ _04369_ _04378_ _03526_ reg_pc\[27\] VGND VGND VPWR VPWR _04379_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09862_ cpuregs\[8\]\[25\] cpuregs\[9\]\[25\] cpuregs\[10\]\[25\] cpuregs\[11\]\[25\]
+ _03586_ _03449_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold1003 cpuregs\[7\]\[19\] VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ _03301_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__clkbuf_4
X_09793_ cpuregs\[4\]\[23\] cpuregs\[5\]\[23\] cpuregs\[6\]\[23\] cpuregs\[7\]\[23\]
+ _03405_ _03496_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__mux4_1
Xhold1014 mem_rdata[3] VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1025 cpuregs\[11\]\[14\] VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 cpuregs\[2\]\[10\] VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 is_sb_sh_sw VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ net825 _03241_ _03185_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _03181_ _01877_ latched_rd\[0\] latched_rd\[1\] VGND VGND VPWR VPWR _03182_
+ sky130_fd_sc_hd__or4bb_1
*XANTENNA_209 net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07626_ _02249_ _02254_ _02257_ _02018_ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_37_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07557_ reg_pc\[16\] decoded_imm\[16\] VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_81_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_49_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07488_ count_instr\[43\] instr_rdinstrh instr_rdcycleh count_cycle\[43\] VGND VGND
+ VPWR VPWR _02129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09227_ decoded_imm\[5\] net198 VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_437 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_134_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09158_ cpuregs\[0\]\[4\] cpuregs\[1\]\[4\] cpuregs\[2\]\[4\] cpuregs\[3\]\[4\] _03458_
+ _03461_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08109_ _02463_ _02701_ _02656_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_79_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09089_ _03446_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11120_ net575 _05089_ _05090_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold870 net155 VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 cpuregs\[1\]\[1\] VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ count_instr\[3\] count_instr\[2\] _05037_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__and3_1
Xhold892 cpuregs\[2\]\[8\] VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__dlygate4sd3_1
X_10002_ net191 _02380_ _03617_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__mux2_1
X_14810_ clknet_leaf_156_clk _00468_ VGND VGND VPWR VPWR cpuregs\[25\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15790_ clknet_leaf_8_clk _01365_ VGND VGND VPWR VPWR cpuregs\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_14741_ clknet_leaf_159_clk _00399_ VGND VGND VPWR VPWR cpuregs\[26\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11953_ instr_srl instr_sll instr_slli instr_srli VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__nor4_2
X_10904_ net1083 _04823_ _04959_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__mux2_1
X_14672_ clknet_leaf_30_clk _00330_ VGND VGND VPWR VPWR cpuregs\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11884_ count_cycle\[50\] net379 VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_15_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ _03385_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__buf_2
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10835_ _04925_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_2
X_13554_ _06942_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10766_ net662 _04821_ _04887_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_81_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12505_ cpuregs\[16\]\[20\] cpuregs\[17\]\[20\] cpuregs\[18\]\[20\] cpuregs\[19\]\[20\]
+ _05948_ _06068_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__mux4_1
X_13485_ net714 _04844_ _06899_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__mux2_1
X_10697_ _03254_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__clkbuf_4
X_15224_ clknet_leaf_76_clk _00817_ VGND VGND VPWR VPWR instr_blt sky130_fd_sc_hd__dfxtp_1
X_12436_ cpuregs\[16\]\[17\] cpuregs\[17\]\[17\] cpuregs\[18\]\[17\] cpuregs\[19\]\[17\]
+ _05948_ _06068_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__mux4_1
X_15155_ clknet_leaf_49_clk _00780_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_1
X_12367_ cpuregs\[20\]\[14\] cpuregs\[21\]\[14\] _05979_ VGND VGND VPWR VPWR _06123_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14106_ _01675_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__clkbuf_1
X_11318_ _05231_ reg_pc\[18\] VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12298_ cpuregs\[0\]\[12\] cpuregs\[1\]\[12\] cpuregs\[2\]\[12\] cpuregs\[3\]\[12\]
+ _06055_ _05909_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__mux4_1
X_15086_ clknet_leaf_81_clk _07140_ VGND VGND VPWR VPWR reg_out\[4\] sky130_fd_sc_hd__dfxtp_1
X_11249_ net546 _05178_ _05169_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__o21ai_1
X_14037_ cpuregs\[6\]\[0\] _06923_ _01638_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14939_ clknet_leaf_120_clk _00597_ VGND VGND VPWR VPWR count_instr\[48\] sky130_fd_sc_hd__dfxtp_1
X_08460_ latched_branch latched_store VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__nand2_4
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07411_ count_instr\[7\] _02054_ count_cycle\[39\] _02055_ VGND VGND VPWR VPWR _02056_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08391_ _01978_ _02950_ _02951_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_663 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_2
X_07342_ _01986_ _01987_ _01989_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_195 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_644 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_724 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07273_ cpu_state\[6\] VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09012_ _01944_ _03481_ _03484_ _03486_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold100 count_cycle\[63\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold111 instr_beq VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 instr_or VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 mem_rdata[13] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold144 count_cycle\[42\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold155 net65 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 count_instr\[50\] VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 count_instr\[39\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold188 instr_srai VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 count_cycle\[12\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ cpuregs\[4\]\[27\] cpuregs\[5\]\[27\] cpuregs\[6\]\[27\] cpuregs\[7\]\[27\]
+ _03439_ _03576_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09845_ cpuregs\[24\]\[24\] cpuregs\[25\]\[24\] cpuregs\[26\]\[24\] cpuregs\[27\]\[24\]
+ _03494_ _03497_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__mux4_2
X_09776_ cpuregs\[8\]\[22\] cpuregs\[9\]\[22\] cpuregs\[10\]\[22\] cpuregs\[11\]\[22\]
+ _03601_ _03583_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__mux4_1
X_08727_ _03223_ _03225_ _03173_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_1_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08658_ _03167_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07609_ _02219_ _02234_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08589_ _03047_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__buf_8
XFILLER_0_138_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10620_ net661 _03263_ _04793_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10551_ _04759_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_510 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10482_ _04722_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__clkbuf_1
X_13270_ net1198 _04833_ _06780_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12221_ _03087_ _05982_ _03153_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12152_ _05912_ _05915_ _03123_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__o21a_1
X_11103_ count_instr\[17\] count_instr\[16\] VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12083_ _03061_ _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11034_ _01905_ net690 VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__and2_1
X_15911_ clknet_leaf_38_clk _01483_ VGND VGND VPWR VPWR cpuregs\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15842_ clknet_leaf_50_clk _01414_ VGND VGND VPWR VPWR cpuregs\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15773_ clknet_leaf_58_clk _01348_ VGND VGND VPWR VPWR cpuregs\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_714 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12985_ decoded_imm\[0\] _06626_ _06628_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_125_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ clknet_leaf_138_clk _00382_ VGND VGND VPWR VPWR cpuregs\[15\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_142_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ cpuregs\[20\]\[31\] cpuregs\[21\]\[31\] cpuregs\[22\]\[31\] cpuregs\[23\]\[31\]
+ _03594_ _03442_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__mux4_1
X_14655_ clknet_leaf_97_clk _00313_ VGND VGND VPWR VPWR cpuregs\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_11867_ _05691_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13606_ cpuregs\[31\]\[25\] _06977_ _06967_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__mux2_1
X_10818_ net1375 _04873_ _04909_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__mux2_1
X_14586_ clknet_leaf_3_clk _00244_ VGND VGND VPWR VPWR cpuregs\[28\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11798_ _05643_ _05625_ _05644_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__and3b_1
XFILLER_0_83_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13537_ _03201_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_41_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10749_ _03366_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xload_slew1 _06576_ VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__buf_1
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13468_ cpuregs\[9\]\[4\] _04827_ _06888_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15207_ clknet_leaf_98_clk alu_out\[20\] VGND VGND VPWR VPWR alu_out_q\[20\] sky130_fd_sc_hd__dfxtp_1
X_12419_ _06073_ _06172_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__or2_1
X_13399_ _06856_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__clkbuf_1
Xoutput205 net205 VGND VGND VPWR VPWR pcpi_rs2[11] sky130_fd_sc_hd__buf_2
XFILLER_0_2_457 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput216 net216 VGND VGND VPWR VPWR pcpi_rs2[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput227 net227 VGND VGND VPWR VPWR pcpi_rs2[31] sky130_fd_sc_hd__buf_2
X_15138_ clknet_leaf_102_clk _00764_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15069_ clknet_leaf_122_clk _00727_ VGND VGND VPWR VPWR count_cycle\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07960_ _02566_ _02578_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_2
X_07891_ _02506_ _02508_ _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09630_ decoded_imm\[16\] net178 net179 decoded_imm\[17\] VGND VGND VPWR VPWR _04087_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09561_ _03894_ _03964_ _03928_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__o21a_1
X_08512_ _01870_ _03032_ _03022_ _00809_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__o2bb2a_1
X_09492_ _03837_ _03953_ _03657_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08443_ reg_next_pc\[19\] reg_out\[19\] _02969_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08374_ _02943_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07325_ _01971_ decoded_imm\[2\] decoded_imm\[1\] reg_pc\[1\] VGND VGND VPWR VPWR
+ _01975_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_129_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07256_ _01848_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__buf_4
XFILLER_0_116_576 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_144_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07187_ _01838_ _01841_ _01843_ _01852_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_76_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09828_ _04275_ _04277_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09759_ _04139_ _04211_ _03483_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_107_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ instr_jalr _01894_ _06503_ latched_branch VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11721_ _05579_ _05581_ _05580_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_739 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ clknet_leaf_64_clk _00098_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_25_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _05246_ _05523_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10603_ net1101 _03209_ _04782_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__mux2_1
X_14371_ net235 _01855_ _06678_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__or3_1
X_11583_ _05452_ _05455_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13322_ _03183_ _04885_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__nor2_4
X_10534_ _04750_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13253_ decoded_imm\[1\] _06531_ _06777_ _06778_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__o22a_1
X_10465_ _04713_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12204_ _03042_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13184_ net781 _06626_ _06737_ _06739_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__o22a_1
X_10396_ net1394 _03202_ _04673_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12135_ _01917_ net245 VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__nor2_4
X_12066_ _03124_ _05835_ _03054_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_127_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11017_ _05021_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__clkbuf_1
X_15825_ clknet_leaf_7_clk _01397_ VGND VGND VPWR VPWR cpuregs\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15756_ clknet_leaf_17_clk _01331_ VGND VGND VPWR VPWR cpuregs\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12968_ decoded_imm_j\[16\] _01078_ _06587_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__mux2_1
X_14707_ clknet_leaf_31_clk _00365_ VGND VGND VPWR VPWR cpuregs\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11919_ _05726_ _05727_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15687_ clknet_leaf_55_clk _01262_ VGND VGND VPWR VPWR cpuregs\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12899_ mem_rdata_q\[20\] _06580_ mem_rdata_q\[21\] VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_118_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14638_ clknet_leaf_44_clk _00296_ VGND VGND VPWR VPWR cpuregs\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14569_ clknet_leaf_19_clk _00227_ VGND VGND VPWR VPWR cpuregs\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_08090_ _02696_ _02697_ _02584_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_155_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_488 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_100_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08992_ _03418_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_71_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07943_ _02562_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_71_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07874_ _02044_ _02492_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__nand2_1
X_09613_ _03448_ _04070_ _03468_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__o21a_1
X_09544_ _03436_ _04003_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_148_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09475_ _03557_ _03936_ _03417_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08426_ _02154_ _02975_ _02971_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_430 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08357_ _01880_ _02489_ net209 _01848_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07308_ net32 net18 _01844_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08288_ net221 net220 net246 _02850_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07239_ _01888_ _01892_ _01894_ _01898_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__or4b_1
XFILLER_0_131_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10250_ _04598_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10181_ latched_rd\[1\] _03181_ _01877_ latched_rd\[0\] VGND VGND VPWR VPWR _04561_
+ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_161_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout251 net122 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_4
X_13940_ net1374 _06964_ _01577_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13871_ net738 _06964_ _07111_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15610_ clknet_leaf_143_clk _01185_ VGND VGND VPWR VPWR cpuregs\[31\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12822_ _06533_ _06532_ _06536_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__and3b_1
X_15541_ clknet_leaf_64_clk _00004_ VGND VGND VPWR VPWR reg_sh\[2\] sky130_fd_sc_hd__dfxtp_1
X_12753_ _03113_ _06491_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11704_ _05032_ _05561_ _05255_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__a21oi_1
X_15472_ clknet_leaf_95_clk _00032_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__dfxtp_4
X_12684_ _06177_ _06421_ _06423_ _06425_ _06164_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14423_ clknet_leaf_60_clk _00081_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dfxtp_4
X_11635_ _05496_ _05498_ _05510_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__a211o_1
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14354_ _01804_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11566_ _05446_ _05447_ _05449_ _05193_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_107_362 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_123_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_123_822 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_764 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13305_ _06806_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10517_ _04740_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__clkbuf_1
X_14285_ net552 VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__clkbuf_1
X_11497_ _05215_ _05380_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_123_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13236_ _06763_ decoded_imm_j\[7\] _06733_ mem_rdata_q\[27\] _06541_ VGND VGND VPWR
+ VPWR _06768_ sky130_fd_sc_hd__a221o_1
X_10448_ net1039 _03367_ _04695_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13167_ latched_rd\[4\] _06724_ _06725_ net436 VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__a22o_1
X_10379_ net685 _03367_ _04658_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12118_ _03096_ cpuregs\[30\]\[5\] _03098_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__o21a_1
X_13098_ _06691_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12049_ _03038_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__buf_6
XFILLER_0_137_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07590_ _02007_ _02222_ _02201_ _02223_ _01955_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__a221o_1
X_15808_ clknet_leaf_73_clk _00025_ VGND VGND VPWR VPWR mem_wordsize\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15739_ clknet_leaf_146_clk _01314_ VGND VGND VPWR VPWR cpuregs\[22\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_886 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09260_ _03727_ _03728_ _03579_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08211_ _02560_ _02568_ _02406_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__mux2_1
X_09191_ _02030_ _03480_ _03482_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08142_ _02732_ _02734_ _02730_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_764 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08073_ _02660_ _02670_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_541 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_585 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08975_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__clkbuf_8
X_07926_ _01931_ _02507_ _02514_ _02515_ _02474_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__a221o_1
Xhold48 net7 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 mem_rdata[26] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ net201 _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07788_ _02395_ _02398_ _02407_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09527_ _03672_ _03969_ _03987_ _03665_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09458_ cpuregs\[4\]\[12\] cpuregs\[5\]\[12\] cpuregs\[6\]\[12\] cpuregs\[7\]\[12\]
+ _03463_ _03464_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08409_ _02082_ _02963_ _02951_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_923 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09389_ _03413_ _03853_ _03418_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11420_ _05313_ _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__or2b_1
XFILLER_0_151_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11351_ _05227_ _05253_ _05254_ _05224_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_120_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10302_ _04626_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14070_ net1256 _06958_ _01649_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11282_ reg_next_pc\[8\] _03230_ _02945_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_115_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13021_ net901 _04839_ _06647_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__mux2_1
X_10233_ net1265 _03334_ _04586_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10164_ _04552_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__clkbuf_1
X_10095_ _04514_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__clkbuf_1
X_14972_ clknet_leaf_106_clk _00630_ VGND VGND VPWR VPWR reg_pc\[18\] sky130_fd_sc_hd__dfxtp_2
X_13923_ _01578_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13854_ _07112_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_137_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12805_ _01901_ decoder_pseudo_trigger VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__nor2_2
X_13785_ cpuregs\[3\]\[10\] _06945_ _07075_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10997_ net1105 _04848_ _05006_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15524_ clknet_leaf_160_clk _01109_ VGND VGND VPWR VPWR cpuregs\[24\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12736_ cpuregs\[22\]\[30\] cpuregs\[23\]\[30\] _05979_ VGND VGND VPWR VPWR _06476_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15455_ clknet_leaf_158_clk _01045_ VGND VGND VPWR VPWR cpuregs\[19\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12667_ cpuregs\[20\]\[27\] cpuregs\[21\]\[27\] _05979_ VGND VGND VPWR VPWR _06410_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ clknet_leaf_59_clk _00027_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_13_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ decoded_imm_j\[20\] _05240_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15386_ clknet_leaf_94_clk _00976_ VGND VGND VPWR VPWR decoded_imm\[22\] sky130_fd_sc_hd__dfxtp_2
X_12598_ _06073_ _06343_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14337_ _01795_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__clkbuf_1
X_11549_ _05432_ _05433_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold507 cpuregs\[1\]\[13\] VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 cpuregs\[19\]\[27\] VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 cpuregs\[21\]\[7\] VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14268_ _01759_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13219_ decoded_imm\[15\] _06752_ _06735_ _06758_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14199_ _01724_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ cpuregs\[11\]\[11\] _03255_ _03249_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07711_ reg_pc\[27\] decoded_imm\[27\] VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__nand2_1
X_08691_ _03195_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__clkbuf_1
X_07642_ reg_pc\[20\] decoded_imm\[20\] decoded_imm\[21\] reg_pc\[21\] VGND VGND VPWR
+ VPWR _02272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07573_ reg_pc\[17\] decoded_imm\[17\] VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09312_ cpuregs\[4\]\[8\] cpuregs\[5\]\[8\] cpuregs\[6\]\[8\] cpuregs\[7\]\[8\] _03641_
+ _03642_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09243_ _03651_ _03707_ _03711_ _03476_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09174_ cpuregs\[20\]\[4\] cpuregs\[21\]\[4\] cpuregs\[22\]\[4\] cpuregs\[23\]\[4\]
+ _03458_ _03461_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_133_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08125_ net176 _02729_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08056_ _02477_ _02655_ _02667_ _02585_ VGND VGND VPWR VPWR alu_out\[8\] sky130_fd_sc_hd__a22o_1
XFILLER_0_141_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput38 net38 VGND VGND VPWR VPWR mem_addr[13] sky130_fd_sc_hd__clkbuf_4
Xpicorv32_260 VGND VGND VPWR VPWR picorv32_260/HI eoi[6] sky130_fd_sc_hd__conb_1
Xpicorv32_271 VGND VGND VPWR VPWR picorv32_271/HI eoi[17] sky130_fd_sc_hd__conb_1
Xoutput49 net49 VGND VGND VPWR VPWR mem_addr[24] sky130_fd_sc_hd__buf_2
Xpicorv32_282 VGND VGND VPWR VPWR picorv32_282/HI eoi[28] sky130_fd_sc_hd__conb_1
Xpicorv32_293 VGND VGND VPWR VPWR picorv32_293/HI pcpi_insn[3] sky130_fd_sc_hd__conb_1
X_08958_ _03426_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__buf_4
X_07909_ _02481_ _02527_ _02528_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__o21ai_1
X_08889_ net889 _03367_ _03315_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ _04958_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10851_ _04933_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__clkbuf_1
X_13570_ _06953_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__clkbuf_1
X_10782_ net1199 _04837_ _04887_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12521_ _06138_ _06269_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15240_ clknet_leaf_76_clk _00833_ VGND VGND VPWR VPWR instr_ori sky130_fd_sc_hd__dfxtp_1
X_12452_ cpuregs\[0\]\[18\] cpuregs\[1\]\[18\] cpuregs\[2\]\[18\] cpuregs\[3\]\[18\]
+ _05819_ _03125_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_10_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11403_ decoder_trigger VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__clkbuf_4
X_15171_ clknet_leaf_56_clk _00796_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dfxtp_4
X_12383_ _03045_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14122_ _01683_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11334_ _05231_ reg_pc\[23\] VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__or2_1
X_14053_ net1320 _06941_ _01638_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11265_ _05193_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__clkbuf_4
X_13004_ net1317 _04823_ _06636_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__mux2_1
X_10216_ net1010 _03282_ _04575_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__mux2_1
X_11196_ _05145_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__clkbuf_1
X_10147_ _04543_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14955_ clknet_leaf_82_clk _00613_ VGND VGND VPWR VPWR reg_pc\[1\] sky130_fd_sc_hd__dfxtp_4
XPHY_EDGE_ROW_145_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10078_ _04505_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13906_ _01569_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__clkbuf_1
X_14886_ clknet_leaf_126_clk _00544_ VGND VGND VPWR VPWR cpuregs\[17\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13837_ _07103_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_18_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_480 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13768_ cpuregs\[3\]\[2\] _06929_ _07064_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15507_ clknet_leaf_87_clk _01092_ VGND VGND VPWR VPWR mem_rdata_q\[30\] sky130_fd_sc_hd__dfxtp_1
X_12719_ cpuregs\[6\]\[30\] cpuregs\[7\]\[30\] _03084_ VGND VGND VPWR VPWR _06459_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_906 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13699_ _07030_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_859 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15438_ clknet_leaf_23_clk _01028_ VGND VGND VPWR VPWR cpuregs\[18\]\[30\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_154_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15369_ clknet_leaf_73_clk _00959_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold304 cpuregs\[0\]\[3\] VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 cpuregs\[0\]\[17\] VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 cpuregs\[28\]\[28\] VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 cpuregs\[4\]\[6\] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 instr_jalr VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09930_ _04371_ _04373_ _04375_ _04377_ _03430_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__a221o_2
XFILLER_0_1_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold359 cpuregs\[13\]\[11\] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09861_ _04309_ _04310_ _03552_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__mux2_1
X_08812_ _03297_ _03300_ _03293_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__mux2_4
X_09792_ _04242_ _04243_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__nor2_1
Xhold1004 cpuregs\[24\]\[8\] VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 cpuregs\[4\]\[19\] VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold1026 cpuregs\[25\]\[19\] VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 count_cycle\[45\] VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ _03240_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__buf_2
Xhold1048 count_cycle\[40\] VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ latched_branch latched_store VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__nor2_2
X_07625_ count_cycle\[20\] _02020_ _02255_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07556_ count_instr\[48\] _02013_ count_cycle\[16\] _02020_ _02191_ VGND VGND VPWR
+ VPWR _02192_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07487_ _01944_ _02125_ _02127_ _01928_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09226_ decoded_imm\[5\] _02030_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09157_ _03448_ _03627_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08108_ _02584_ _02712_ _02713_ _02715_ _02464_ VGND VGND VPWR VPWR alu_out\[12\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_79_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09088_ cpuregs\[20\]\[2\] cpuregs\[21\]\[2\] cpuregs\[22\]\[2\] cpuregs\[23\]\[2\]
+ _03554_ _03459_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08039_ _02066_ _02489_ _02561_ _02595_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_112_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold860 cpuregs\[24\]\[15\] VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 cpuregs\[8\]\[17\] VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 count_instr\[47\] VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _05039_ net995 VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__nor2_1
Xhold893 cpuregs\[11\]\[5\] VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__dlygate4sd3_1
X_10001_ _03475_ _04446_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__and2_1
X_14740_ clknet_leaf_159_clk _00398_ VGND VGND VPWR VPWR cpuregs\[26\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11952_ _03476_ _05750_ _05752_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10903_ _04961_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__clkbuf_1
X_14671_ clknet_leaf_38_clk _00329_ VGND VGND VPWR VPWR cpuregs\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11883_ _05702_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_631 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13622_ _06988_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10834_ net819 _04821_ _04923_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_67_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13553_ net1343 _06941_ _06925_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10765_ _04888_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12504_ _06142_ _06253_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__or2_1
X_13484_ _06901_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__clkbuf_1
X_10696_ _04841_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15223_ clknet_leaf_77_clk _00816_ VGND VGND VPWR VPWR instr_bne sky130_fd_sc_hd__dfxtp_1
X_12435_ _06142_ _06187_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15154_ clknet_leaf_67_clk _00779_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_1
X_12366_ _06119_ _06120_ _06121_ _05873_ _03113_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14105_ cpuregs\[7\]\[0\] _06923_ _01674_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11317_ _01891_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__clkbuf_2
X_15085_ clknet_leaf_81_clk _07139_ VGND VGND VPWR VPWR reg_out\[3\] sky130_fd_sc_hd__dfxtp_1
X_12297_ _05907_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__buf_6
X_14036_ _01637_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__buf_6
X_11248_ count_instr\[62\] count_instr\[61\] net475 _05175_ VGND VGND VPWR VPWR _05181_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_129_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11179_ net535 _05130_ _05133_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_147_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14938_ clknet_leaf_121_clk _00596_ VGND VGND VPWR VPWR count_instr\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_54_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14869_ clknet_leaf_159_clk _00527_ VGND VGND VPWR VPWR cpuregs\[17\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_817 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07410_ _01947_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_46_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08390_ _01816_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07341_ _01986_ _01987_ _01989_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_656 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07272_ _01840_ is_lb_lh_lw_lbu_lhu _01838_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09011_ _03485_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_155_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold101 mem_rdata[14] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 count_instr\[33\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold123 mem_rdata[12] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold134 reg_next_pc\[21\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold145 count_cycle\[25\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold156 count_cycle\[39\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 count_instr\[56\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_463 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold178 cpuregs\[0\]\[18\] VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _02331_ _03624_ _04361_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__a21o_1
Xhold189 instr_srli VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09844_ _04293_ _04294_ _03437_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__mux2_1
X_09775_ _03454_ _04227_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__or2_1
X_08726_ reg_out\[7\] alu_out_q\[7\] latched_stalu VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_428 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08657_ decoded_imm_j\[3\] _01085_ _03022_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07608_ _02019_ _02231_ _02240_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__o21a_1
X_08588_ _03046_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__clkbuf_8
X_07539_ _02172_ _02173_ _02174_ _01893_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_48_174 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_325 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_91_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10550_ net967 _03255_ _04757_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09209_ _03500_ _03678_ _03468_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10481_ cpuregs\[14\]\[11\] _03255_ _04720_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__mux2_1
X_12220_ cpuregs\[22\]\[8\] cpuregs\[23\]\[8\] _05816_ VGND VGND VPWR VPWR _05982_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12151_ cpuregs\[12\]\[6\] cpuregs\[13\]\[6\] cpuregs\[14\]\[6\] cpuregs\[15\]\[6\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11102_ net465 VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12082_ cpuregs\[16\]\[1\] cpuregs\[17\]\[1\] cpuregs\[18\]\[1\] cpuregs\[19\]\[1\]
+ _03091_ _03125_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__mux4_1
Xhold690 cpuregs\[23\]\[6\] VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11033_ _05029_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__clkbuf_1
X_15910_ clknet_leaf_43_clk _01482_ VGND VGND VPWR VPWR cpuregs\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_129_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ clknet_leaf_22_clk _01413_ VGND VGND VPWR VPWR cpuregs\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15772_ clknet_leaf_102_clk _01347_ VGND VGND VPWR VPWR cpuregs\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12984_ net1406 net445 _06627_ mem_rdata_q\[20\] _06553_ VGND VGND VPWR VPWR _06628_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_125_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14723_ clknet_leaf_97_clk _00381_ VGND VGND VPWR VPWR cpuregs\[15\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11935_ _03575_ _05735_ _05737_ _05739_ _03489_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_142_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14654_ clknet_leaf_21_clk _00312_ VGND VGND VPWR VPWR cpuregs\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_11866_ _05689_ _01842_ _05690_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__and3b_1
XFILLER_0_86_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13605_ _03347_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__clkbuf_4
X_10817_ _04915_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14585_ clknet_leaf_3_clk _00243_ VGND VGND VPWR VPWR cpuregs\[28\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11797_ count_cycle\[22\] _05640_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13536_ _06930_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__clkbuf_1
X_10748_ _04876_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_41_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_706 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13467_ _06892_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__clkbuf_1
X_10679_ net1142 _04829_ _04819_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15206_ clknet_leaf_98_clk alu_out\[19\] VGND VGND VPWR VPWR alu_out_q\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12418_ cpuregs\[24\]\[16\] cpuregs\[25\]\[16\] cpuregs\[26\]\[16\] cpuregs\[27\]\[16\]
+ _06074_ _05932_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__mux4_1
X_13398_ cpuregs\[24\]\[3\] _04825_ _06852_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__mux2_1
Xoutput206 net206 VGND VGND VPWR VPWR pcpi_rs2[12] sky130_fd_sc_hd__clkbuf_4
Xoutput217 net217 VGND VGND VPWR VPWR pcpi_rs2[22] sky130_fd_sc_hd__buf_2
X_15137_ clknet_leaf_102_clk _00763_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12349_ _06105_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__clkbuf_1
Xoutput228 net228 VGND VGND VPWR VPWR pcpi_rs2[3] sky130_fd_sc_hd__buf_2
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15068_ clknet_leaf_123_clk _00726_ VGND VGND VPWR VPWR count_cycle\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14019_ net1339 _06975_ _01624_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__mux2_1
X_07890_ net193 _02509_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09560_ _03962_ _04010_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__or2b_1
X_08511_ _01945_ is_beq_bne_blt_bge_bltu_bgeu _02558_ VGND VGND VPWR VPWR _03032_
+ sky130_fd_sc_hd__and3_1
X_09491_ _02139_ _03617_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__nor2_1
X_08442_ _02986_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08373_ _02489_ net218 _01932_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07324_ reg_pc\[1\] decoded_imm\[1\] _01972_ _01973_ VGND VGND VPWR VPWR _01974_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_61_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07255_ _01912_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__clkbuf_1
X_07186_ cpu_state\[0\] _01851_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ _04213_ _04239_ _04276_ _04151_ _04240_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__o221a_1
X_09758_ _02331_ _03660_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_107_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08709_ reg_pc\[5\] _03206_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__and2_1
X_09689_ _02306_ _03619_ _04077_ _03075_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__a211o_1
X_11720_ _05261_ _05584_ _05367_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11651_ _05418_ net452 _05343_ _05527_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10602_ _04786_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14370_ _01812_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__clkbuf_1
X_11582_ _05453_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13321_ _06814_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10533_ cpuregs\[27\]\[3\] _03202_ _04746_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_823 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13252_ _06763_ decoded_imm_j\[1\] _06732_ net852 _06540_ VGND VGND VPWR VPWR _06778_
+ sky130_fd_sc_hd__a221o_1
X_10464_ net1305 _03202_ _04709_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__mux2_1
X_12203_ cpuregs\[8\]\[8\] cpuregs\[9\]\[8\] cpuregs\[10\]\[8\] cpuregs\[11\]\[8\]
+ _05907_ _03047_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__mux4_1
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13183_ mem_rdata_q\[31\] _06738_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__and2_1
X_10395_ _04676_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12134_ _03083_ _05894_ _05898_ _05886_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12065_ cpuregs\[28\]\[0\] cpuregs\[29\]\[0\] cpuregs\[30\]\[0\] cpuregs\[31\]\[0\]
+ _05834_ _03097_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_127_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ cpuregs\[17\]\[23\] _04867_ _05017_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15824_ clknet_leaf_142_clk _01396_ VGND VGND VPWR VPWR cpuregs\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_512 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15755_ clknet_leaf_4_clk _01330_ VGND VGND VPWR VPWR cpuregs\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12967_ _06618_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11918_ net824 _05724_ _05141_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__o21ai_1
X_14706_ clknet_leaf_56_clk _00364_ VGND VGND VPWR VPWR cpuregs\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12898_ _02055_ _06554_ _06581_ _06582_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__a22o_1
X_15686_ clknet_leaf_34_clk _01261_ VGND VGND VPWR VPWR cpuregs\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11849_ _05678_ _05679_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14637_ clknet_leaf_39_clk _00295_ VGND VGND VPWR VPWR cpuregs\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_431 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_16_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14568_ clknet_leaf_58_clk _00226_ VGND VGND VPWR VPWR cpuregs\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_16_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13519_ _06919_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__clkbuf_1
X_14499_ clknet_leaf_130_clk _00157_ VGND VGND VPWR VPWR cpuregs\[30\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_569 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08991_ _03436_ _03465_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__or2_1
X_07942_ instr_or instr_ori VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_71_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07873_ net199 _02492_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__or2_1
X_09612_ cpuregs\[28\]\[17\] cpuregs\[29\]\[17\] cpuregs\[30\]\[17\] cpuregs\[31\]\[17\]
+ _03680_ _03443_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__mux4_1
X_09543_ cpuregs\[24\]\[15\] cpuregs\[25\]\[15\] cpuregs\[26\]\[15\] cpuregs\[27\]\[15\]
+ _03594_ _03442_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__mux4_2
X_09474_ cpuregs\[8\]\[13\] cpuregs\[9\]\[13\] cpuregs\[10\]\[13\] cpuregs\[11\]\[13\]
+ _03586_ _03449_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08425_ reg_next_pc\[13\] reg_out\[13\] _02969_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__mux2_2
XFILLER_0_65_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08356_ _02466_ _02927_ _02934_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__a21o_2
XFILLER_0_117_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07307_ _01953_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08287_ _02432_ _02581_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07238_ cpu_state\[4\] _01897_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07169_ instr_fence instr_and instr_lbu instr_lb VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10180_ _04560_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_161_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout252 net195 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_4
X_13870_ _01549_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12821_ _05803_ _06541_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_122_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ clknet_leaf_19_clk _01125_ VGND VGND VPWR VPWR cpuregs\[24\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12752_ cpuregs\[20\]\[31\] cpuregs\[21\]\[31\] cpuregs\[22\]\[31\] cpuregs\[23\]\[31\]
+ _03095_ _03144_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_159_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _05571_ _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__xnor2_1
X_15471_ clknet_leaf_18_clk _01061_ VGND VGND VPWR VPWR cpuregs\[19\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12683_ _06138_ _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14422_ clknet_leaf_61_clk _00080_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dfxtp_2
X_11634_ _05497_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14353_ net628 _03333_ _01800_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__mux2_1
X_11565_ _05367_ _05448_ net361 VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13304_ net1088 _04867_ _06802_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10516_ net1189 _03367_ _04731_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14284_ _01767_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11496_ _05372_ _05375_ _05383_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__o21ai_1
X_13235_ decoded_imm\[8\] _06626_ _06767_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10447_ _04703_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13166_ latched_rd\[3\] _06724_ _06725_ net439 VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10378_ _04666_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_591 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12117_ cpuregs\[31\]\[5\] _03096_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__or2b_1
X_13097_ net162 net249 _06685_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12048_ _03124_ _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15807_ clknet_leaf_73_clk _00024_ VGND VGND VPWR VPWR mem_wordsize\[0\] sky130_fd_sc_hd__dfxtp_1
X_13999_ _01618_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15738_ clknet_leaf_144_clk _01313_ VGND VGND VPWR VPWR cpuregs\[22\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_526 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_932 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15669_ clknet_leaf_144_clk _01244_ VGND VGND VPWR VPWR cpuregs\[29\]\[22\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_190 _06191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08210_ _02801_ _02808_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09190_ _01992_ _03660_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08141_ _02744_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08072_ _02680_ _02681_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_597 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08974_ _00013_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07925_ _02394_ _02544_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__nor2_1
Xhold49 mem_rdata[1] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07856_ net233 VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_27_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07787_ _02405_ _02406_ _02400_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__a21bo_1
X_09526_ reg_pc\[14\] _03528_ _03986_ _03626_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ _03746_ _03919_ _03603_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08408_ reg_next_pc\[8\] reg_out\[8\] _02949_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09388_ cpuregs\[8\]\[10\] cpuregs\[9\]\[10\] cpuregs\[10\]\[10\] cpuregs\[11\]\[10\]
+ _03404_ _03408_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_935 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08339_ _02925_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_151_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11350_ _05231_ reg_pc\[28\] VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10301_ net1248 _03334_ _04622_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11281_ _05186_ _05204_ _05205_ _01885_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__o211a_1
X_13020_ _06635_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_115_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10232_ _04589_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10163_ net1068 _03334_ _04548_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_58_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10094_ net747 _03341_ _04509_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__mux2_1
X_14971_ clknet_leaf_105_clk _00629_ VGND VGND VPWR VPWR reg_pc\[17\] sky130_fd_sc_hd__dfxtp_2
X_13922_ cpuregs\[4\]\[10\] _06945_ _01577_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_89_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13853_ net1273 _06945_ _07111_ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__mux2_1
X_12804_ _06525_ _06513_ _06518_ _06527_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__a22o_1
X_10996_ _05010_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__clkbuf_1
X_13784_ _07063_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_684 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15523_ clknet_leaf_153_clk _01108_ VGND VGND VPWR VPWR cpuregs\[24\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12735_ _05872_ _06474_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_139_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _06406_ _06407_ _06408_ _05873_ _05845_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__a221o_1
X_15454_ clknet_leaf_152_clk _01044_ VGND VGND VPWR VPWR cpuregs\[19\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11617_ _05495_ _05237_ _05488_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__a21o_1
X_14405_ clknet_leaf_21_clk _00068_ VGND VGND VPWR VPWR cpuregs\[11\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ cpuregs\[24\]\[24\] cpuregs\[25\]\[24\] cpuregs\[26\]\[24\] cpuregs\[27\]\[24\]
+ _06074_ _03151_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_13_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15385_ clknet_leaf_94_clk _00975_ VGND VGND VPWR VPWR decoded_imm\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_142_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14336_ net589 _03281_ _01789_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__mux2_1
X_11548_ decoded_imm_j\[16\] _05225_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_123_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold508 cpuregs\[27\]\[31\] VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ net611 VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__clkbuf_1
Xhold519 cpuregs\[10\]\[28\] VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11479_ _05184_ _05210_ _05269_ _05344_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__or4_1
XFILLER_0_111_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13218_ _06525_ decoded_imm_j\[15\] _06738_ mem_rdata_q\[15\] VGND VGND VPWR VPWR
+ _06758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14198_ net1129 _06950_ _01721_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__mux2_1
X_13149_ net1141 net120 _06684_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07710_ reg_pc\[27\] decoded_imm\[27\] VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__or2_1
X_08690_ cpuregs\[11\]\[2\] _03194_ _03185_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07641_ _02269_ _02270_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__and2_1
X_07572_ count_instr\[17\] _02054_ count_cycle\[17\] _02020_ _02206_ VGND VGND VPWR
+ VPWR _02207_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09311_ _03415_ _03777_ _03420_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_66_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09242_ _03657_ _03708_ _03710_ _01953_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_378 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09173_ _03455_ _03643_ _03468_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_32_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08124_ net176 _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_631 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_32_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08055_ _02662_ _02666_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_261 VGND VGND VPWR VPWR picorv32_261/HI eoi[7] sky130_fd_sc_hd__conb_1
Xoutput39 net39 VGND VGND VPWR VPWR mem_addr[14] sky130_fd_sc_hd__clkbuf_4
Xpicorv32_272 VGND VGND VPWR VPWR picorv32_272/HI eoi[18] sky130_fd_sc_hd__conb_1
Xpicorv32_283 VGND VGND VPWR VPWR picorv32_283/HI eoi[29] sky130_fd_sc_hd__conb_1
Xpicorv32_294 VGND VGND VPWR VPWR picorv32_294/HI pcpi_insn[4] sky130_fd_sc_hd__conb_1
X_08957_ _03412_ _03421_ _03423_ _03428_ _03431_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__o221a_1
X_07908_ _02112_ net248 VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__or2b_1
X_08888_ _03366_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_86_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07839_ _02458_ net223 _02442_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__and3_1
X_10850_ cpuregs\[25\]\[9\] _04837_ _04923_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09509_ cpuregs\[20\]\[14\] cpuregs\[21\]\[14\] cpuregs\[22\]\[14\] cpuregs\[23\]\[14\]
+ _03587_ _03588_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__mux4_1
X_10781_ _04896_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__clkbuf_1
X_12520_ cpuregs\[8\]\[21\] cpuregs\[9\]\[21\] cpuregs\[10\]\[21\] cpuregs\[11\]\[21\]
+ _06061_ _03137_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_594 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_136_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12451_ _05925_ _06202_ _03050_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_10_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11402_ _05289_ _05293_ _05295_ _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_117_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15170_ clknet_leaf_62_clk _00795_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_151_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12382_ _06058_ _06136_ _03123_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_491 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_90 _04958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14121_ net1054 _06941_ _01674_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__mux2_1
X_11333_ reg_next_pc\[23\] _03331_ _02947_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__mux2_2
XFILLER_0_132_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14052_ _01646_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__clkbuf_1
X_11264_ _01891_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13003_ _06638_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__clkbuf_1
X_10215_ _04580_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__clkbuf_1
X_11195_ _05143_ _05113_ _05144_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__and3b_1
X_10146_ cpuregs\[30\]\[15\] _03282_ _04537_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__mux2_1
X_14954_ clknet_leaf_115_clk _00612_ VGND VGND VPWR VPWR count_instr\[63\] sky130_fd_sc_hd__dfxtp_1
X_10077_ net787 _03287_ _04498_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__mux2_1
X_13905_ cpuregs\[4\]\[2\] _06929_ _01566_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__mux2_1
X_14885_ clknet_leaf_151_clk _00543_ VGND VGND VPWR VPWR cpuregs\[17\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13836_ net688 _06929_ _07100_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13767_ _07066_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__clkbuf_1
X_10979_ _05001_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__clkbuf_1
X_15506_ clknet_leaf_87_clk _01091_ VGND VGND VPWR VPWR mem_rdata_q\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_127_211 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12718_ _05871_ _06457_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13698_ net1018 _06927_ _07028_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15437_ clknet_leaf_125_clk _01027_ VGND VGND VPWR VPWR cpuregs\[18\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12649_ _06392_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_882 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15368_ clknet_leaf_75_clk _00958_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold305 cpuregs\[16\]\[2\] VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ net1194 _03227_ _01778_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__mux2_1
Xhold316 cpuregs\[25\]\[12\] VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ clknet_leaf_35_clk _00889_ VGND VGND VPWR VPWR cpuregs\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold327 count_cycle\[51\] VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold338 cpuregs\[4\]\[27\] VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 cpuregs\[19\]\[5\] VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09860_ cpuregs\[0\]\[25\] cpuregs\[1\]\[25\] cpuregs\[2\]\[25\] cpuregs\[3\]\[25\]
+ _03800_ _03407_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__mux4_1
X_08811_ _03298_ _03299_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__nor2_1
X_09791_ _04213_ _04238_ _04241_ _01870_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__a31o_1
Xhold1005 cpuregs\[15\]\[23\] VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 cpuregs\[16\]\[26\] VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 cpuregs\[1\]\[20\] VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _03173_ _03237_ _03238_ _03239_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__a22o_2
Xhold1038 net134 VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 count_cycle\[25\] VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08673_ latched_rd\[4\] latched_rd\[2\] latched_rd\[3\] VGND VGND VPWR VPWR _03180_
+ sky130_fd_sc_hd__or3b_4
X_07624_ count_instr\[20\] _01965_ count_cycle\[52\] _02014_ VGND VGND VPWR VPWR _02256_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_95_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07555_ count_instr\[16\] _01965_ count_cycle\[48\] _02014_ VGND VGND VPWR VPWR _02191_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_119_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07486_ _02083_ _02126_ _02085_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09225_ _03652_ _03655_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09156_ cpuregs\[4\]\[4\] cpuregs\[5\]\[4\] cpuregs\[6\]\[4\] cpuregs\[7\]\[4\] _03458_
+ _03461_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08107_ _02465_ _02569_ _02714_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09087_ _03547_ _03553_ _03556_ _03559_ _03489_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_110_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_110_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_79_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08038_ _02066_ _02489_ _02593_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_112_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold850 cpuregs\[27\]\[8\] VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 cpuregs\[8\]\[20\] VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_678 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold872 cpuregs\[7\]\[24\] VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold883 cpuregs\[13\]\[1\] VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 cpuregs\[26\]\[23\] VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _03472_ _04436_ _04445_ _03525_ reg_pc\[29\] VGND VGND VPWR VPWR _04446_
+ sky130_fd_sc_hd__a32o_1
X_09989_ _03552_ _04434_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__or2_1
X_11951_ _05754_ _05755_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__nor2_1
X_10902_ net891 _04821_ _04959_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__mux2_1
X_11882_ _05700_ _01842_ _05701_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14670_ clknet_leaf_44_clk _00328_ VGND VGND VPWR VPWR cpuregs\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13621_ net736 _06987_ _06924_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__mux2_1
X_10833_ _04924_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13552_ _03234_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__buf_2
X_10764_ net1056 _04817_ _04887_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12503_ cpuregs\[20\]\[20\] cpuregs\[21\]\[20\] cpuregs\[22\]\[20\] cpuregs\[23\]\[20\]
+ _06065_ _03144_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__mux4_1
X_13483_ net1040 _04842_ _06899_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_501 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10695_ cpuregs\[26\]\[10\] _04839_ _04840_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12434_ cpuregs\[20\]\[17\] cpuregs\[21\]\[17\] cpuregs\[22\]\[17\] cpuregs\[23\]\[17\]
+ _06065_ _05922_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__mux4_1
X_15222_ clknet_leaf_77_clk _00815_ VGND VGND VPWR VPWR instr_beq sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12365_ cpuregs\[28\]\[14\] cpuregs\[29\]\[14\] _03085_ VGND VGND VPWR VPWR _06121_
+ sky130_fd_sc_hd__mux2_1
X_15153_ clknet_leaf_69_clk _00778_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_101_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_101_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_105_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11316_ reg_next_pc\[18\] _03297_ _02947_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__mux2_2
X_14104_ _01673_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__buf_6
X_15084_ clknet_leaf_72_clk _07136_ VGND VGND VPWR VPWR reg_out\[2\] sky130_fd_sc_hd__dfxtp_1
X_12296_ cpuregs\[4\]\[12\] cpuregs\[5\]\[12\] cpuregs\[6\]\[12\] cpuregs\[7\]\[12\]
+ _06011_ _03097_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__mux4_1
X_14035_ _04524_ _01564_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__nor2_2
XFILLER_0_129_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11247_ _05180_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11178_ _05040_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_147_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10129_ net699 _03228_ _04526_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14937_ clknet_leaf_121_clk _00595_ VGND VGND VPWR VPWR count_instr\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14868_ clknet_leaf_158_clk _00526_ VGND VGND VPWR VPWR cpuregs\[17\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_148_829 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13819_ _07093_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14799_ clknet_leaf_43_clk _00457_ VGND VGND VPWR VPWR cpuregs\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07340_ _01988_ _01975_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07271_ _01922_ _01925_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_203 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_92_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09010_ _03388_ _01864_ _03393_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__or3b_4
XFILLER_0_14_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold102 decoded_imm_j\[16\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 instr_ori VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 reg_next_pc\[27\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 count_instr\[1\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 count_instr\[54\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_598 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold157 count_instr\[20\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 reg_next_pc\[15\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09912_ _03672_ _04342_ _04360_ _03665_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__o211a_1
Xhold179 instr_blt VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09843_ cpuregs\[20\]\[24\] cpuregs\[21\]\[24\] cpuregs\[22\]\[24\] cpuregs\[23\]\[24\]
+ _03636_ _03637_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_13_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09774_ cpuregs\[12\]\[22\] cpuregs\[13\]\[22\] cpuregs\[14\]\[22\] cpuregs\[15\]\[22\]
+ _03598_ _03716_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__mux4_1
X_08725_ _03199_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_159_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_159_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08656_ _03166_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _02058_ _02236_ _02239_ _02071_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08587_ _03045_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07538_ _02172_ _02173_ _02174_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_862 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_48_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07469_ _02074_ _02079_ _02108_ _02107_ _02094_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09208_ cpuregs\[8\]\[5\] cpuregs\[9\]\[5\] cpuregs\[10\]\[5\] cpuregs\[11\]\[5\]
+ _03636_ _03637_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10480_ _04721_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09139_ decoded_imm\[3\] net196 VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12150_ _03063_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_94_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11101_ _05079_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__clkbuf_1
X_12081_ _05840_ _05842_ _05844_ _05847_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__o32a_1
Xhold680 cpuregs\[21\]\[28\] VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold691 cpuregs\[30\]\[4\] VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ net759 _04883_ _04994_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ clknet_leaf_25_clk _01412_ VGND VGND VPWR VPWR cpuregs\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15771_ clknet_leaf_129_clk _01346_ VGND VGND VPWR VPWR cpuregs\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12983_ instr_jalr is_lb_lh_lw_lbu_lhu is_alu_reg_imm VGND VGND VPWR VPWR _06627_
+ sky130_fd_sc_hd__or3_4
X_14722_ clknet_leaf_136_clk _00380_ VGND VGND VPWR VPWR cpuregs\[15\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11934_ _03447_ _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_142_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14653_ clknet_leaf_14_clk _00311_ VGND VGND VPWR VPWR cpuregs\[14\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11865_ count_cycle\[43\] _05686_ count_cycle\[44\] VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13604_ _06976_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10816_ net1298 _04871_ _04909_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14584_ clknet_leaf_143_clk _00242_ VGND VGND VPWR VPWR cpuregs\[28\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11796_ count_cycle\[22\] _05640_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_851 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13535_ net766 _06929_ _06925_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__mux2_1
X_10747_ net1078 _04875_ _04861_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_605 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_82_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13466_ net1382 _04825_ _06888_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__mux2_1
X_10678_ _03214_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__buf_2
XFILLER_0_153_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_23_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15205_ clknet_leaf_99_clk alu_out\[18\] VGND VGND VPWR VPWR alu_out_q\[18\] sky130_fd_sc_hd__dfxtp_1
X_12417_ _06026_ _06170_ _03081_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__o21a_1
X_13397_ _06855_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__clkbuf_1
Xoutput207 net207 VGND VGND VPWR VPWR pcpi_rs2[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput218 net218 VGND VGND VPWR VPWR pcpi_rs2[23] sky130_fd_sc_hd__buf_2
X_15136_ clknet_leaf_112_clk _00762_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12348_ _02471_ _06104_ _06052_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__mux2_1
Xoutput229 net229 VGND VGND VPWR VPWR pcpi_rs2[4] sky130_fd_sc_hd__buf_2
X_15067_ clknet_leaf_122_clk _00725_ VGND VGND VPWR VPWR count_cycle\[50\] sky130_fd_sc_hd__dfxtp_1
X_12279_ _05912_ _06037_ _03123_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__o21a_1
X_14018_ _01628_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__clkbuf_1
X_15969_ clknet_leaf_21_clk _01541_ VGND VGND VPWR VPWR cpuregs\[10\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_08510_ _03031_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__clkbuf_1
X_09490_ _02213_ _03617_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__and2_1
X_08441_ _02222_ _02985_ _02971_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_604 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08372_ _02942_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_98_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07323_ _01971_ decoded_imm\[2\] VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07254_ _01905_ _01851_ _01911_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_882 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07185_ mem_do_rinst reg_pc\[1\] _01850_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_76_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_793 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ _04153_ _04178_ _04177_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__o21a_1
X_09757_ _02290_ _03619_ _04209_ _03616_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_107_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _03210_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__clkbuf_1
X_09688_ _04143_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08639_ _03142_ _03148_ _03156_ net244 VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__a31o_1
X_11650_ _05285_ _05245_ _05526_ _05300_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10601_ cpuregs\[15\]\[3\] _03202_ _04782_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__mux2_1
X_11581_ _05461_ _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13320_ net1295 _04883_ _06779_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10532_ _04749_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10463_ _04712_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__clkbuf_1
X_13251_ mem_rdata_q\[21\] _06627_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12202_ cpuregs\[12\]\[8\] cpuregs\[13\]\[8\] cpuregs\[14\]\[8\] cpuregs\[15\]\[8\]
+ _03107_ _03129_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__mux4_1
X_13182_ _01823_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__clkbuf_4
X_10394_ net590 _03194_ _04673_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_384 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12133_ _03090_ _05897_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12064_ _03046_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__buf_8
X_11015_ _05020_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_144_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ clknet_leaf_16_clk _01395_ VGND VGND VPWR VPWR cpuregs\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15754_ clknet_leaf_8_clk _01329_ VGND VGND VPWR VPWR cpuregs\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12966_ decoded_imm_j\[15\] _01077_ _06587_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14705_ clknet_leaf_34_clk _00363_ VGND VGND VPWR VPWR cpuregs\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11917_ count_cycle\[60\] _05724_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__and2_1
X_15685_ clknet_leaf_32_clk _01260_ VGND VGND VPWR VPWR cpuregs\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12897_ net564 _06575_ net443 VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_142_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14636_ clknet_leaf_28_clk _00294_ VGND VGND VPWR VPWR cpuregs\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11848_ net630 _05675_ _05647_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14567_ clknet_leaf_133_clk _00225_ VGND VGND VPWR VPWR cpuregs\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11779_ count_cycle\[16\] count_cycle\[17\] _05628_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13518_ net1234 _04877_ _06910_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__mux2_1
X_14498_ clknet_leaf_129_clk _00156_ VGND VGND VPWR VPWR cpuregs\[30\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13449_ _06882_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15119_ clknet_leaf_74_clk _00745_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08990_ cpuregs\[24\]\[0\] cpuregs\[25\]\[0\] cpuregs\[26\]\[0\] cpuregs\[27\]\[0\]
+ _03463_ _03464_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__mux4_1
X_07941_ _02560_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_71_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07872_ net125 VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__clkbuf_4
X_09611_ _03437_ _04068_ _03426_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__o21a_1
X_09542_ _03402_ _04001_ _03603_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__o21a_1
X_09473_ _03933_ _03934_ _03552_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_90_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_2
X_08424_ _02974_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_456 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08355_ _01880_ _02492_ _02466_ _01913_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07306_ _01928_ _01941_ _01957_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08286_ _02340_ net222 _02561_ _02563_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07237_ _01895_ _01896_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07168_ instr_sltu instr_slt instr_sw instr_sh VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_161_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout253 net191 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__buf_4
X_09809_ _04254_ _04256_ _04258_ _04260_ _03760_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_89_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12820_ _06540_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12751_ _06177_ _06485_ _06487_ _06489_ _03142_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_2
X_11702_ _05572_ _05573_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__nand2_1
X_15470_ clknet_leaf_23_clk _01060_ VGND VGND VPWR VPWR cpuregs\[19\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12682_ cpuregs\[8\]\[28\] cpuregs\[9\]\[28\] cpuregs\[10\]\[28\] cpuregs\[11\]\[28\]
+ _05970_ _03137_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14421_ clknet_leaf_57_clk _00079_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dfxtp_2
X_11633_ _05488_ _05507_ _05510_ _05498_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_108_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_92_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14352_ _01803_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__clkbuf_1
X_11564_ _05414_ _05228_ _05225_ _05222_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__and4b_1
XFILLER_0_135_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _06805_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__clkbuf_1
X_10515_ _04739_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_137_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14283_ net581 VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__clkbuf_1
X_11495_ _05372_ _05375_ _05383_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__or3_1
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10446_ cpuregs\[21\]\[27\] _03360_ _04695_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__mux2_1
X_13234_ _06763_ decoded_imm_j\[8\] _06733_ mem_rdata_q\[28\] _06541_ VGND VGND VPWR
+ VPWR _06767_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10377_ net1104 _03360_ _04658_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__mux2_1
X_13165_ latched_rd\[2\] _06724_ _06725_ net427 VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12116_ cpuregs\[24\]\[5\] cpuregs\[25\]\[5\] cpuregs\[26\]\[5\] cpuregs\[27\]\[5\]
+ _03096_ _03098_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__mux4_1
X_13096_ _06690_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12047_ cpuregs\[4\]\[0\] cpuregs\[5\]\[0\] cpuregs\[6\]\[0\] cpuregs\[7\]\[0\] _05816_
+ _03086_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__mux4_1
X_15806_ clknet_leaf_22_clk _01381_ VGND VGND VPWR VPWR cpuregs\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13998_ net1243 _06954_ _01613_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__mux2_1
X_15737_ clknet_leaf_153_clk _01312_ VGND VGND VPWR VPWR cpuregs\[22\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_12949_ _06609_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_72_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_87_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15668_ clknet_leaf_121_clk _01243_ VGND VGND VPWR VPWR cpuregs\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
*XANTENNA_180 _04877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_191 _06759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14619_ clknet_leaf_0_clk _00277_ VGND VGND VPWR VPWR cpuregs\[21\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15599_ clknet_leaf_6_clk _01174_ VGND VGND VPWR VPWR cpuregs\[31\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08140_ net177 _02743_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08071_ net172 _02679_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08973_ _03447_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__buf_6
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07924_ _02461_ _02542_ _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__or3b_2
X_07855_ net205 VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07786_ _02250_ net215 VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__nand2_1
X_09525_ _03574_ _03977_ _03985_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_63_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_2
X_09456_ cpuregs\[8\]\[12\] cpuregs\[9\]\[12\] cpuregs\[10\]\[12\] cpuregs\[11\]\[12\]
+ _03601_ _03583_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_84_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08407_ _02962_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_1
X_09387_ _03401_ _03851_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08338_ _02251_ _01937_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08269_ _02316_ _02863_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__xnor2_1
X_10300_ _04625_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11280_ _05188_ reg_pc\[7\] VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10231_ cpuregs\[13\]\[22\] _03329_ _04586_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10162_ _04551_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_5_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10093_ _04513_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__clkbuf_1
X_14970_ clknet_leaf_106_clk _00628_ VGND VGND VPWR VPWR reg_pc\[16\] sky130_fd_sc_hd__dfxtp_2
X_13921_ _01565_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__buf_4
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13852_ _07099_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__buf_4
X_12803_ _01065_ _01064_ _06526_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13783_ _07074_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__clkbuf_1
X_10995_ cpuregs\[17\]\[13\] _04846_ _05006_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_54_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_2
X_15522_ clknet_leaf_153_clk _01107_ VGND VGND VPWR VPWR cpuregs\[24\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12734_ cpuregs\[20\]\[30\] cpuregs\[21\]\[30\] _03084_ VGND VGND VPWR VPWR _06474_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_696 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ clknet_leaf_151_clk _01043_ VGND VGND VPWR VPWR cpuregs\[19\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12665_ cpuregs\[28\]\[27\] cpuregs\[29\]\[27\] _03085_ VGND VGND VPWR VPWR _06408_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_155_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14404_ clknet_leaf_22_clk _00067_ VGND VGND VPWR VPWR cpuregs\[11\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11616_ _05494_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15384_ clknet_leaf_94_clk _00974_ VGND VGND VPWR VPWR decoded_imm\[24\] sky130_fd_sc_hd__dfxtp_2
X_12596_ _05912_ _06341_ _06193_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14335_ _01794_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__clkbuf_1
X_11547_ decoded_imm_j\[16\] _05225_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_152_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_788 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_122_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold509 cpuregs\[16\]\[5\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ _01758_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__clkbuf_1
X_11478_ _05289_ _05364_ _05366_ _05368_ _05184_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13217_ decoded_imm\[16\] _06752_ _06735_ _06757_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__o22a_1
X_10429_ net629 _03307_ _04684_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14197_ _01723_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13148_ _06717_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_78 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13079_ _01839_ _06679_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__nand2_1
X_07640_ reg_pc\[22\] decoded_imm\[22\] VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07571_ count_instr\[49\] _02052_ _02014_ count_cycle\[49\] VGND VGND VPWR VPWR _02206_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_45_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09310_ cpuregs\[8\]\[8\] cpuregs\[9\]\[8\] cpuregs\[10\]\[8\] cpuregs\[11\]\[8\]
+ _03494_ _03497_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_66_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09241_ _02066_ _03480_ _03709_ _03482_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09172_ cpuregs\[28\]\[4\] cpuregs\[29\]\[4\] cpuregs\[30\]\[4\] cpuregs\[31\]\[4\]
+ _03641_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08123_ _02466_ _02728_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_585 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08054_ _02625_ _02663_ _02637_ _02648_ _02665_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__a41o_1
XFILLER_0_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_262 VGND VGND VPWR VPWR picorv32_262/HI eoi[8] sky130_fd_sc_hd__conb_1
Xpicorv32_273 VGND VGND VPWR VPWR picorv32_273/HI eoi[19] sky130_fd_sc_hd__conb_1
Xpicorv32_284 VGND VGND VPWR VPWR picorv32_284/HI eoi[30] sky130_fd_sc_hd__conb_1
Xpicorv32_295 VGND VGND VPWR VPWR picorv32_295/HI pcpi_insn[5] sky130_fd_sc_hd__conb_1
XFILLER_0_110_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08956_ _03430_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__buf_6
X_07907_ _02099_ _02525_ _02526_ _02082_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__o22a_1
X_08887_ _03362_ _03365_ _03199_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_86_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07838_ net253 VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__inv_2
X_07769_ reg_pc\[31\] decoded_imm\[31\] VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_36_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09508_ _01958_ _03958_ _03960_ _03397_ _03968_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_156_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10780_ net1334 _04835_ _04887_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09439_ _03898_ _03900_ _03895_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_251 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_82_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12450_ cpuregs\[6\]\[18\] cpuregs\[7\]\[18\] _03084_ VGND VGND VPWR VPWR _06202_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11401_ _05197_ _05283_ _05297_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_117_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_917 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12381_ cpuregs\[12\]\[15\] cpuregs\[13\]\[15\] cpuregs\[14\]\[15\] cpuregs\[15\]\[15\]
+ _05913_ _05994_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_134_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_80 _04839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_91 _05815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14120_ _01682_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__clkbuf_1
X_11332_ _05194_ net709 _05239_ _05241_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_793 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_132_484 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14051_ cpuregs\[6\]\[7\] _06939_ _01638_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11263_ _05186_ _05191_ _05192_ _01885_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13002_ net1240 _04821_ _06636_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__mux2_1
X_10214_ net1300 _03275_ _04575_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__mux2_1
X_11194_ count_instr\[44\] net381 count_instr\[45\] VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__a21o_1
X_10145_ _04542_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__clkbuf_1
X_14953_ clknet_leaf_117_clk _00611_ VGND VGND VPWR VPWR count_instr\[62\] sky130_fd_sc_hd__dfxtp_1
X_10076_ _04504_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
X_13904_ _01568_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__clkbuf_1
X_14884_ clknet_leaf_149_clk _00542_ VGND VGND VPWR VPWR cpuregs\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_13835_ _07102_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_18_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13766_ net763 _06927_ _07064_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10978_ net831 _04829_ _04995_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15505_ clknet_leaf_88_clk _01090_ VGND VGND VPWR VPWR mem_rdata_q\[28\] sky130_fd_sc_hd__dfxtp_1
X_12717_ cpuregs\[4\]\[30\] cpuregs\[5\]\[30\] _03051_ VGND VGND VPWR VPWR _06457_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13697_ _07029_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15436_ clknet_leaf_148_clk _01026_ VGND VGND VPWR VPWR cpuregs\[18\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12648_ net221 _06391_ _06282_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15367_ clknet_leaf_73_clk _00957_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dfxtp_1
X_12579_ _06319_ _06321_ _06323_ _06325_ _06151_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14318_ _01785_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold306 cpuregs\[13\]\[30\] VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ clknet_leaf_26_clk _00888_ VGND VGND VPWR VPWR cpuregs\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold317 cpuregs\[22\]\[31\] VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 cpuregs\[15\]\[2\] VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold339 cpuregs\[2\]\[25\] VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ net613 VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_68_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08810_ reg_pc\[18\] _03291_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__and2_1
X_09790_ _04213_ _04238_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__a21oi_1
Xhold1006 cpuregs\[27\]\[7\] VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 cpuregs\[20\]\[0\] VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ reg_pc\[9\] _03232_ _03199_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__o21a_1
Xhold1028 cpuregs\[27\]\[0\] VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 count_instr\[16\] VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08672_ _03178_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_77_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07623_ count_instr\[52\] _01946_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_18_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07554_ _02187_ _02190_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XFILLER_0_9_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_76_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07485_ _01846_ _01848_ net20 net3 _01933_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09224_ _01977_ _03668_ _03671_ _03672_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09155_ _03625_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08106_ _02139_ _02463_ _02618_ _02641_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__a31o_1
X_09086_ _03557_ _03558_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08037_ _02648_ _02649_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold840 cpuregs\[16\]\[9\] VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold851 mem_rdata_q\[28\] VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold862 reg_pc\[12\] VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold873 cpuregs\[12\]\[21\] VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 cpuregs\[5\]\[14\] VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 cpuregs\[27\]\[27\] VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__dlygate4sd3_1
X_09988_ cpuregs\[12\]\[29\] cpuregs\[13\]\[29\] cpuregs\[14\]\[29\] cpuregs\[15\]\[29\]
+ _03808_ _03801_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__mux4_1
X_08939_ _03413_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_95_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11950_ _04453_ _04457_ _05753_ _01869_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__a31o_1
X_10901_ _04960_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__clkbuf_1
X_11881_ count_cycle\[48\] _05695_ count_cycle\[49\] VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__a21o_1
X_13620_ _03380_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__clkbuf_4
X_10832_ net874 _04817_ _04923_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_201 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13551_ _06940_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10763_ _04886_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_463 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12502_ _06177_ _06247_ _06249_ _06251_ _06164_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__a221o_1
X_13482_ _06900_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__clkbuf_1
X_10694_ _04818_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15221_ clknet_leaf_78_clk _00814_ VGND VGND VPWR VPWR instr_jal sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_43_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12433_ _06177_ _06180_ _06183_ _06185_ _06164_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15152_ clknet_leaf_71_clk _00777_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_1
X_12364_ _05974_ cpuregs\[30\]\[14\] _05896_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14103_ _03183_ _01564_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__nor2_2
X_11315_ _05227_ _05228_ _05229_ _05224_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__o211a_1
X_15083_ clknet_leaf_91_clk _07125_ VGND VGND VPWR VPWR reg_out\[1\] sky130_fd_sc_hd__dfxtp_1
X_12295_ _06053_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__clkbuf_1
X_14034_ _01636_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__clkbuf_1
X_11246_ _05178_ _05113_ _05179_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__and3b_1
XFILLER_0_129_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11177_ count_instr\[40\] count_instr\[39\] count_instr\[38\] _05127_ VGND VGND VPWR
+ VPWR _05132_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_147_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10128_ _04533_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14936_ clknet_leaf_121_clk _00594_ VGND VGND VPWR VPWR count_instr\[45\] sky130_fd_sc_hd__dfxtp_1
X_10059_ _04495_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14867_ clknet_leaf_29_clk _00525_ VGND VGND VPWR VPWR cpuregs\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13818_ net1125 _06979_ _07086_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14798_ clknet_leaf_45_clk _00456_ VGND VGND VPWR VPWR cpuregs\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13749_ _07056_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07270_ cpu_state\[5\] _01887_ _01924_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15419_ clknet_leaf_159_clk _01009_ VGND VGND VPWR VPWR cpuregs\[18\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_14_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold103 count_instr\[5\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold114 count_cycle\[44\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold125 mem_rdata_q\[23\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold136 _00550_ VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold147 count_cycle\[40\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold158 reg_next_pc\[19\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ reg_pc\[26\] _03528_ _04359_ _03626_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__a211o_1
Xhold169 count_cycle\[3\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09842_ cpuregs\[16\]\[24\] cpuregs\[17\]\[24\] cpuregs\[18\]\[24\] cpuregs\[19\]\[24\]
+ _03636_ _03637_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09773_ _03433_ _04221_ _04223_ _04225_ _03760_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__a221o_1
X_08724_ reg_pc\[6\] reg_pc\[5\] _03206_ reg_pc\[7\] VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__a31o_1
X_08655_ mem_rdata_q\[23\] net16 _03017_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07606_ _02065_ _02237_ _02201_ _02238_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__a22o_1
X_08586_ cpuregs\[20\]\[3\] cpuregs\[21\]\[3\] cpuregs\[22\]\[3\] cpuregs\[23\]\[3\]
+ _03092_ _03098_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__mux4_1
XFILLER_0_135_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_817 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07537_ _02161_ _02163_ _02160_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_688 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07468_ _02107_ _02109_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_716 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_107_738 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09207_ _03675_ _03676_ _03402_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__mux2_1
X_07399_ net6 net24 _01845_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09138_ _03539_ _03540_ _03541_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_20_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09069_ _03539_ _03540_ _03541_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11100_ _01884_ _05077_ _05078_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12080_ _03128_ _05848_ _03035_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__o21ai_1
Xhold670 cpuregs\[4\]\[16\] VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold681 cpuregs\[9\]\[11\] VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 cpuregs\[5\]\[20\] VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _05028_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_129_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15770_ clknet_leaf_138_clk _01345_ VGND VGND VPWR VPWR cpuregs\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12982_ _06531_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__clkbuf_4
X_14721_ clknet_leaf_137_clk _00379_ VGND VGND VPWR VPWR cpuregs\[15\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_11933_ cpuregs\[12\]\[31\] cpuregs\[13\]\[31\] cpuregs\[14\]\[31\] cpuregs\[15\]\[31\]
+ _03719_ _03588_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_142_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14652_ clknet_leaf_14_clk _00310_ VGND VGND VPWR VPWR cpuregs\[14\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11864_ count_cycle\[43\] net473 _05686_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13603_ net800 _06975_ _06967_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _04914_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__clkbuf_1
X_14583_ clknet_leaf_154_clk _00241_ VGND VGND VPWR VPWR cpuregs\[28\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11795_ _05642_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13534_ _03193_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_198 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10746_ _03359_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13465_ _06891_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10677_ _04828_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__clkbuf_1
X_15204_ clknet_leaf_98_clk alu_out\[17\] VGND VGND VPWR VPWR alu_out_q\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12416_ cpuregs\[28\]\[16\] cpuregs\[29\]\[16\] cpuregs\[30\]\[16\] cpuregs\[31\]\[16\]
+ _05895_ _05929_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13396_ net1291 _04823_ _06852_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15135_ clknet_leaf_102_clk _00761_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dfxtp_1
Xoutput208 net208 VGND VGND VPWR VPWR pcpi_rs2[14] sky130_fd_sc_hd__clkbuf_4
X_12347_ _05901_ _06090_ _06103_ _05904_ decoded_imm\[13\] VGND VGND VPWR VPWR _06104_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_590 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput219 net246 VGND VGND VPWR VPWR pcpi_rs2[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15066_ clknet_leaf_121_clk _00724_ VGND VGND VPWR VPWR count_cycle\[49\] sky130_fd_sc_hd__dfxtp_1
X_12278_ cpuregs\[12\]\[11\] cpuregs\[13\]\[11\] cpuregs\[14\]\[11\] cpuregs\[15\]\[11\]
+ _05913_ _05994_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14017_ net957 _06973_ _01624_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__mux2_1
X_11229_ count_instr\[56\] count_instr\[55\] count_instr\[54\] _05162_ VGND VGND VPWR
+ VPWR _05168_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ clknet_leaf_22_clk _01540_ VGND VGND VPWR VPWR cpuregs\[10\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_14919_ clknet_leaf_117_clk _00577_ VGND VGND VPWR VPWR count_instr\[28\] sky130_fd_sc_hd__dfxtp_1
X_15899_ clknet_leaf_101_clk _01471_ VGND VGND VPWR VPWR cpuregs\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08440_ reg_next_pc\[18\] reg_out\[18\] _02969_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08371_ _02492_ net217 _01932_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_129_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07322_ _01971_ decoded_imm\[2\] VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_98_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07253_ cpu_state\[3\] is_beq_bne_blt_bge_bltu_bgeu _01886_ _01910_ _01840_ VGND
+ VGND VPWR VPWR _01911_ sky130_fd_sc_hd__a32o_1
XFILLER_0_155_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_144_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07184_ mem_do_wdata mem_do_rdata _01846_ _01847_ _01849_ VGND VGND VPWR VPWR _01850_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09825_ _04155_ _04180_ _04275_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__or3_1
X_09756_ _02265_ net243 VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__and2_1
X_08707_ net1332 _03209_ _03185_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _02237_ _04142_ _03395_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08638_ _03149_ _03152_ _03155_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08569_ cpuregs\[4\]\[3\] cpuregs\[5\]\[3\] cpuregs\[6\]\[3\] cpuregs\[7\]\[3\] _03085_
+ _03087_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ _04785_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11580_ decoded_imm_j\[19\] _05233_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_582 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_107_524 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10531_ net1070 _03194_ _04746_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13250_ decoded_imm\[2\] _06531_ _06775_ _06776_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10462_ net653 _03194_ _04709_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12201_ _05959_ _05961_ _05962_ _03128_ _03035_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_847 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13181_ _06736_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__buf_2
XFILLER_0_150_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10393_ _04675_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_396 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12132_ cpuregs\[8\]\[5\] cpuregs\[9\]\[5\] cpuregs\[10\]\[5\] cpuregs\[11\]\[5\]
+ _05895_ _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12063_ _03061_ _05832_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__or2_1
X_11014_ net829 _04865_ _05017_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ clknet_leaf_5_clk _01394_ VGND VGND VPWR VPWR cpuregs\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15753_ clknet_leaf_8_clk _01328_ VGND VGND VPWR VPWR cpuregs\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_12965_ _06617_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__clkbuf_1
X_11916_ _05724_ _05725_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__nor2_1
X_14704_ clknet_leaf_32_clk _00362_ VGND VGND VPWR VPWR cpuregs\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15684_ clknet_leaf_41_clk _01259_ VGND VGND VPWR VPWR cpuregs\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12896_ instr_rdcycle _06554_ _06576_ _06581_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14635_ clknet_leaf_56_clk _00293_ VGND VGND VPWR VPWR cpuregs\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11847_ count_cycle\[37\] count_cycle\[38\] _05673_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_260 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14566_ clknet_leaf_134_clk _00224_ VGND VGND VPWR VPWR cpuregs\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11778_ net561 _05628_ _05630_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13517_ _06918_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__clkbuf_1
X_10729_ cpuregs\[26\]\[21\] _04863_ _04861_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__mux2_1
X_14497_ clknet_leaf_145_clk _00155_ VGND VGND VPWR VPWR cpuregs\[30\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13448_ net837 _04875_ _06874_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13379_ _06845_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15118_ clknet_leaf_75_clk _00744_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_1
X_15049_ clknet_leaf_115_clk _00707_ VGND VGND VPWR VPWR count_cycle\[32\] sky130_fd_sc_hd__dfxtp_1
X_07940_ _02559_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07871_ net200 _02489_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_3_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ cpuregs\[16\]\[17\] cpuregs\[17\]\[17\] cpuregs\[18\]\[17\] cpuregs\[19\]\[17\]
+ _03673_ _03674_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__mux4_1
X_09541_ cpuregs\[28\]\[15\] cpuregs\[29\]\[15\] cpuregs\[30\]\[15\] cpuregs\[31\]\[15\]
+ _03601_ _03492_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09472_ cpuregs\[0\]\[13\] cpuregs\[1\]\[13\] cpuregs\[2\]\[13\] cpuregs\[3\]\[13\]
+ _03800_ _03407_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_402 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08423_ _02139_ _02973_ _02971_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ _02471_ _02927_ _02933_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_22_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07305_ _01847_ _01944_ decoded_imm\[0\] _01945_ _01956_ VGND VGND VPWR VPWR _01957_
+ sky130_fd_sc_hd__a221o_1
X_08285_ _02584_ _02875_ _02876_ _02878_ _02426_ VGND VGND VPWR VPWR alu_out\[26\]
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_117_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07236_ reg_sh\[1\] reg_sh\[0\] VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__or2_2
XFILLER_0_15_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07167_ instr_or instr_sra instr_srl instr_xor VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__or4_1
XFILLER_0_112_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09808_ _03414_ _04259_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__or2_1
X_09739_ _03807_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_122_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12750_ _05969_ _06488_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _05495_ _05255_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12681_ _03143_ _06422_ _06182_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14420_ clknet_leaf_61_clk _00078_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dfxtp_4
X_11632_ _05508_ _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14351_ cpuregs\[10\]\[22\] _03328_ _01800_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11563_ _05445_ _05442_ _05444_ _01889_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13302_ net1211 _04865_ _06802_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__mux2_1
X_10514_ cpuregs\[14\]\[27\] _03360_ _04731_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _01766_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_137_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11494_ decoded_imm_j\[12\] _05215_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13233_ decoded_imm\[9\] _06626_ _06766_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__o21a_1
X_10445_ _04702_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13164_ latched_rd\[1\] _06724_ _06725_ net433 VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__a22o_1
X_10376_ _04665_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_150_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12115_ _05875_ _05877_ _05878_ _03090_ _05879_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__o221a_1
X_13095_ net161 net250 _06685_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12046_ _03038_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__clkbuf_8
X_15805_ clknet_leaf_22_clk _01380_ VGND VGND VPWR VPWR cpuregs\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_13997_ _01617_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15736_ clknet_leaf_128_clk _01311_ VGND VGND VPWR VPWR cpuregs\[22\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12948_ net437 _01069_ _06587_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15667_ clknet_leaf_146_clk _01242_ VGND VGND VPWR VPWR cpuregs\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_170 _03548_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12879_ _05041_ net242 _06569_ _06529_ net669 VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__a32o_1
*XANTENNA_181 _05040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_192 decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14618_ clknet_leaf_0_clk _00276_ VGND VGND VPWR VPWR cpuregs\[21\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15598_ clknet_leaf_2_clk _01173_ VGND VGND VPWR VPWR cpuregs\[31\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14549_ clknet_leaf_7_clk _00207_ VGND VGND VPWR VPWR cpuregs\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08070_ net172 _02679_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08972_ _03446_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__clkbuf_8
X_07923_ net194 _02394_ net226 VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__or3b_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07854_ _02464_ _02465_ _02473_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__a21o_1
X_07785_ _02250_ net215 VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ _03979_ _03981_ _03984_ _03433_ _03591_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09455_ _03454_ _03917_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08406_ _02066_ _02961_ _02951_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09386_ cpuregs\[12\]\[10\] cpuregs\[13\]\[10\] cpuregs\[14\]\[10\] cpuregs\[15\]\[10\]
+ _03554_ _03459_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__mux4_1
X_08337_ _01930_ _01847_ _01933_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__a21o_1
XFILLER_0_145_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08268_ net220 _02862_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07219_ instr_slt net491 net538 VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__or3_1
X_08199_ _02250_ _02798_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__and2_1
X_10230_ _04588_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_198 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10161_ cpuregs\[30\]\[22\] _03329_ _04548_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__mux2_1
X_10092_ net764 _03334_ _04509_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__mux2_1
X_13920_ _01576_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__clkbuf_1
X_13851_ _07110_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__clkbuf_1
X_12802_ _01066_ _01068_ _01067_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13782_ net1076 _06943_ _07064_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__mux2_1
X_10994_ _05009_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15521_ clknet_leaf_157_clk _01106_ VGND VGND VPWR VPWR cpuregs\[24\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12733_ _06470_ _06471_ _06472_ _05872_ _05845_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15452_ clknet_leaf_158_clk _01042_ VGND VGND VPWR VPWR cpuregs\[19\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _05974_ cpuregs\[30\]\[27\] _05896_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_106_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14403_ clknet_leaf_136_clk _00066_ VGND VGND VPWR VPWR cpuregs\[11\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_11615_ decoded_imm_j\[20\] VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_26_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15383_ clknet_leaf_89_clk _00973_ VGND VGND VPWR VPWR decoded_imm\[25\] sky130_fd_sc_hd__dfxtp_2
X_12595_ cpuregs\[28\]\[24\] cpuregs\[29\]\[24\] cpuregs\[30\]\[24\] cpuregs\[31\]\[24\]
+ _06191_ _05914_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_13_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14334_ net1262 _03274_ _01789_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11546_ _05222_ _05225_ _05429_ _05288_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_482 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14265_ net594 VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11477_ _05367_ net361 VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__nand2_2
XFILLER_0_123_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13216_ _06525_ net461 _06738_ mem_rdata_q\[16\] VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__a22o_1
X_10428_ _04693_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14196_ cpuregs\[8\]\[11\] _06948_ _01721_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13147_ net156 net118 _06707_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__mux2_1
X_10359_ _04656_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__clkbuf_1
X_13078_ _03020_ _01855_ _06678_ net235 VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__a211o_1
X_12029_ _01891_ _01840_ cpu_state\[0\] VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__nor3_1
XFILLER_0_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07570_ _02019_ _02192_ _02205_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15719_ clknet_leaf_25_clk _01294_ VGND VGND VPWR VPWR cpuregs\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_124_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09240_ _02030_ net243 VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09171_ _03492_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08122_ _02656_ _02727_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_542 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_255 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08053_ _02633_ _02664_ _02647_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_597 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_133_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpicorv32_263 VGND VGND VPWR VPWR picorv32_263/HI eoi[9] sky130_fd_sc_hd__conb_1
Xpicorv32_274 VGND VGND VPWR VPWR picorv32_274/HI eoi[20] sky130_fd_sc_hd__conb_1
Xpicorv32_285 VGND VGND VPWR VPWR picorv32_285/HI eoi[31] sky130_fd_sc_hd__conb_1
Xpicorv32_296 VGND VGND VPWR VPWR picorv32_296/HI pcpi_insn[6] sky130_fd_sc_hd__conb_1
X_08955_ _03429_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__clkbuf_8
X_07906_ _02476_ _02483_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__nand2_1
X_08886_ _03363_ _03364_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_86_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07837_ _02450_ net222 _02456_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_86_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07768_ _02376_ _02378_ _02375_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09507_ _03966_ _03967_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_156_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07699_ reg_pc\[26\] decoded_imm\[26\] VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09438_ _03895_ _03898_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09369_ _03832_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11400_ _05288_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12380_ _06133_ _06134_ _06014_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__mux2_1
*XANTENNA_70 _03588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
*XANTENNA_81 _04842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_929 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_105_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_406 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_90_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_50_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11331_ _01872_ _05240_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__or2_1
*XANTENNA_92 _05827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14050_ _01645_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__clkbuf_1
X_11262_ _05188_ _01971_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13001_ _06637_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__clkbuf_1
X_10213_ _04579_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__clkbuf_1
X_11193_ count_instr\[45\] net513 _05139_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__and3_1
X_10144_ cpuregs\[30\]\[14\] _03275_ _04537_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14952_ clknet_leaf_117_clk _00610_ VGND VGND VPWR VPWR count_instr\[61\] sky130_fd_sc_hd__dfxtp_1
X_10075_ cpuregs\[12\]\[15\] _03282_ _04498_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13903_ cpuregs\[4\]\[1\] _06927_ _01566_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__mux2_1
X_14883_ clknet_leaf_125_clk _00541_ VGND VGND VPWR VPWR cpuregs\[17\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13834_ net588 _06927_ _07100_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13765_ _07065_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_174 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10977_ _05000_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15504_ clknet_leaf_88_clk _01089_ VGND VGND VPWR VPWR mem_rdata_q\[27\] sky130_fd_sc_hd__dfxtp_1
X_12716_ _06456_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__clkbuf_1
X_13696_ net945 _06923_ _07028_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15435_ clknet_leaf_151_clk _01025_ VGND VGND VPWR VPWR cpuregs\[18\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12647_ _05900_ _06377_ _06390_ _01918_ decoded_imm\[26\] VGND VGND VPWR VPWR _06391_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_155_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15366_ clknet_leaf_74_clk _00956_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dfxtp_1
X_12578_ _06073_ _06324_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11529_ _05368_ _05411_ _05412_ _05415_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__o31a_1
X_14317_ cpuregs\[10\]\[6\] _03220_ _01778_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__mux2_1
X_15297_ clknet_leaf_50_clk _00887_ VGND VGND VPWR VPWR cpuregs\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold307 cpuregs\[0\]\[12\] VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold318 reg_next_pc\[11\] VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold329 cpuregs\[22\]\[2\] VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ _01749_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14179_ net1389 _06931_ _01710_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold1007 cpuregs\[20\]\[29\] VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__dlygate4sd3_1
X_08740_ reg_pc\[9\] _03232_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__nand2_1
Xhold1018 cpuregs\[7\]\[30\] VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 cpuregs\[21\]\[30\] VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__dlygate4sd3_1
X_08671_ _03173_ _03177_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_68_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07622_ _02007_ _02250_ _02201_ _02253_ _01968_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__a221o_1
X_07553_ count_cycle\[15\] _02051_ _02189_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_37_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07484_ net173 VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09223_ _03474_ _03683_ _03692_ _03527_ reg_pc\[5\] VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_583 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_57_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09154_ cpu_state\[4\] _01854_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08105_ _02706_ _02711_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_141_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09085_ cpuregs\[8\]\[2\] cpuregs\[9\]\[2\] cpuregs\[10\]\[2\] cpuregs\[11\]\[2\]
+ _03456_ _03441_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08036_ _02635_ _02638_ _02633_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__o21ai_1
Xhold830 cpuregs\[14\]\[28\] VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold841 cpuregs\[14\]\[23\] VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold852 cpuregs\[18\]\[22\] VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold863 cpuregs\[12\]\[22\] VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 cpuregs\[20\]\[3\] VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 cpuregs\[23\]\[4\] VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 cpuregs\[9\]\[5\] VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__dlygate4sd3_1
X_09987_ _03557_ _04432_ _03417_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__o21a_1
X_08938_ _00014_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_150_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08869_ reg_out\[26\] alu_out_q\[26\] _03176_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10900_ net1376 _04817_ _04959_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__mux2_1
X_11880_ count_cycle\[46\] count_cycle\[47\] _05692_ _05699_ VGND VGND VPWR VPWR _05700_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_67_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10831_ _04922_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13550_ net701 _06939_ _06925_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__mux2_1
X_10762_ _04485_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__nor2_4
XFILLER_0_27_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12501_ _06138_ _06250_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13481_ net642 _04839_ _06899_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10693_ _03247_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__clkbuf_4
X_15220_ clknet_leaf_78_clk _00813_ VGND VGND VPWR VPWR instr_auipc sky130_fd_sc_hd__dfxtp_1
X_12432_ _06138_ _06184_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15151_ clknet_leaf_69_clk _00776_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_1
X_12363_ cpuregs\[31\]\[14\] _03092_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__or2b_1
XFILLER_0_90_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14102_ _01672_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__clkbuf_1
X_11314_ _05188_ reg_pc\[17\] VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__or2_1
X_15082_ clknet_leaf_72_clk _07114_ VGND VGND VPWR VPWR reg_out\[0\] sky130_fd_sc_hd__dfxtp_1
X_12294_ net205 _06051_ _06052_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14033_ net1060 _06989_ _01601_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11245_ count_instr\[60\] _05175_ count_instr\[61\] VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11176_ _05130_ _05131_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__nor2_1
X_10127_ net1166 _03221_ _04526_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14935_ clknet_leaf_113_clk _00593_ VGND VGND VPWR VPWR count_instr\[44\] sky130_fd_sc_hd__dfxtp_1
X_10058_ cpuregs\[12\]\[7\] _03228_ _04487_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14866_ clknet_leaf_25_clk _00524_ VGND VGND VPWR VPWR cpuregs\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13817_ _07092_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__clkbuf_1
X_14797_ clknet_leaf_37_clk _00455_ VGND VGND VPWR VPWR cpuregs\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13748_ net586 _06977_ _07050_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_57_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_380 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13679_ _07019_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15418_ clknet_leaf_159_clk _01008_ VGND VGND VPWR VPWR cpuregs\[18\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15349_ clknet_leaf_69_clk _00939_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold104 _00554_ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 instr_blt VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 mem_rdata[21] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold137 reg_next_pc\[1\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 count_cycle\[30\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 count_instr\[23\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09910_ _03574_ _04350_ _04358_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09841_ _04286_ _04288_ _04291_ _03434_ _03490_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__a221o_1
X_09772_ _03593_ _04224_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__or2_1
X_08723_ reg_pc\[7\] reg_pc\[6\] _03211_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08654_ _03165_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07605_ net11 _02202_ _02179_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08585_ _00011_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07536_ reg_pc\[15\] decoded_imm\[15\] VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07467_ _02108_ _02097_ _02094_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09206_ cpuregs\[0\]\[5\] cpuregs\[1\]\[5\] cpuregs\[2\]\[5\] cpuregs\[3\]\[5\] _03673_
+ _03674_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_151_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07398_ net199 VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__buf_4
X_09137_ decoded_imm\[3\] net196 VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09068_ decoded_imm\[2\] net193 VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__and2_1
X_08019_ net199 _02632_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__nand2_1
Xhold660 cpuregs\[27\]\[23\] VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 cpuregs\[26\]\[9\] VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold682 cpuregs\[13\]\[21\] VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net917 _04881_ _04994_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__mux2_1
Xhold693 cpuregs\[2\]\[11\] VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _06625_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__clkbuf_1
X_14720_ clknet_leaf_138_clk _00378_ VGND VGND VPWR VPWR cpuregs\[15\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11932_ _03581_ _05736_ _03467_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ net565 net360 _05688_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__a21oi_1
X_14651_ clknet_leaf_10_clk _00309_ VGND VGND VPWR VPWR cpuregs\[14\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10814_ cpuregs\[16\]\[24\] _04869_ _04909_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _03340_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_45_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ clknet_leaf_154_clk _00240_ VGND VGND VPWR VPWR cpuregs\[28\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11794_ _05640_ _05625_ _05641_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10745_ _04874_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__clkbuf_1
X_13533_ _06928_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_54_147 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13464_ net939 _04823_ _06888_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__mux2_1
X_10676_ net1266 _04827_ _04819_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12415_ _06023_ _06168_ _05927_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__o21a_1
X_15203_ clknet_leaf_97_clk alu_out\[16\] VGND VGND VPWR VPWR alu_out_q\[16\] sky130_fd_sc_hd__dfxtp_1
X_13395_ _06854_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12346_ _05886_ _06092_ _06096_ _05978_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__a311o_2
X_15134_ clknet_leaf_102_clk _00760_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput209 net209 VGND VGND VPWR VPWR pcpi_rs2[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15065_ clknet_leaf_121_clk _00723_ VGND VGND VPWR VPWR count_cycle\[48\] sky130_fd_sc_hd__dfxtp_1
X_12277_ _06034_ _06035_ _06014_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__mux2_1
X_14016_ _01627_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11228_ _05167_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_56_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11159_ count_instr\[35\] count_instr\[34\] _05116_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15967_ clknet_leaf_101_clk _01539_ VGND VGND VPWR VPWR cpuregs\[10\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14918_ clknet_leaf_117_clk _00576_ VGND VGND VPWR VPWR count_instr\[27\] sky130_fd_sc_hd__dfxtp_1
X_15898_ clknet_leaf_133_clk _01470_ VGND VGND VPWR VPWR cpuregs\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14849_ clknet_leaf_147_clk _00507_ VGND VGND VPWR VPWR cpuregs\[20\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08370_ _02941_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_1
XFILLER_0_81_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07321_ reg_pc\[2\] VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_98_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_129_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07252_ _01906_ _01909_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_350 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07183_ _01847_ _01848_ mem_wordsize\[0\] VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_111_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09824_ _04215_ _04241_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__or2_1
X_09755_ _04208_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08706_ _03208_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__buf_2
X_09686_ _03651_ _04118_ _04137_ _04141_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_107_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _03153_ _03154_ _03054_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08568_ _03086_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07519_ _02058_ _02153_ _02157_ _02071_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_25_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ mem_rdata_q\[17\] net9 _03018_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10530_ _04748_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_536 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_134_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10461_ _04711_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12200_ cpuregs\[0\]\[8\] cpuregs\[1\]\[8\] cpuregs\[2\]\[8\] cpuregs\[3\]\[8\] _03091_
+ _03125_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__mux4_1
X_13180_ _05289_ _05495_ _06735_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10392_ net601 _03189_ _04673_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__mux2_1
X_12131_ _03063_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__clkbuf_8
X_12062_ cpuregs\[24\]\[0\] cpuregs\[25\]\[0\] cpuregs\[26\]\[0\] cpuregs\[27\]\[0\]
+ _03091_ _03125_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__mux4_1
Xhold490 cpuregs\[9\]\[26\] VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ _05019_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_144_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ clknet_leaf_7_clk _01393_ VGND VGND VPWR VPWR cpuregs\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15752_ clknet_leaf_32_clk _01327_ VGND VGND VPWR VPWR cpuregs\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12964_ net436 _01073_ _06587_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14703_ clknet_leaf_39_clk _00361_ VGND VGND VPWR VPWR cpuregs\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11915_ net490 _05721_ _05647_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15683_ clknet_leaf_43_clk _01258_ VGND VGND VPWR VPWR cpuregs\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12895_ mem_rdata_q\[21\] _06580_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_68_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14634_ clknet_leaf_54_clk _00292_ VGND VGND VPWR VPWR cpuregs\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11846_ _05677_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11777_ count_cycle\[16\] _05628_ _05622_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14565_ clknet_leaf_20_clk _00223_ VGND VGND VPWR VPWR cpuregs\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10728_ _03321_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__clkbuf_4
X_13516_ net865 _04875_ _06910_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__mux2_1
X_14496_ clknet_leaf_144_clk _00154_ VGND VGND VPWR VPWR cpuregs\[30\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13447_ _06881_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__clkbuf_1
X_10659_ net1276 _03386_ _04781_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13378_ net755 _04873_ _06838_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15117_ clknet_leaf_74_clk _00743_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_1
X_12329_ cpuregs\[12\]\[13\] cpuregs\[13\]\[13\] cpuregs\[14\]\[13\] cpuregs\[15\]\[13\]
+ _03107_ _03129_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15048_ clknet_leaf_114_clk _00706_ VGND VGND VPWR VPWR count_cycle\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07870_ _02489_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ _03581_ _03999_ _03547_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__o21a_1
X_09471_ cpuregs\[4\]\[13\] cpuregs\[5\]\[13\] cpuregs\[6\]\[13\] cpuregs\[7\]\[13\]
+ _03800_ _03801_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_751 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08422_ reg_next_pc\[12\] reg_out\[12\] _02969_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__mux2_2
XFILLER_0_148_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_626 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_650 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08353_ _01880_ net249 _02471_ _01913_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07304_ _01948_ _01952_ _01955_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__o21a_2
XFILLER_0_116_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08284_ _02427_ _02569_ _02877_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07235_ reg_sh\[3\] reg_sh\[2\] reg_sh\[4\] VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__or3_2
XFILLER_0_6_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07166_ _01829_ _01830_ _01831_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_161_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09807_ cpuregs\[24\]\[23\] cpuregs\[25\]\[23\] cpuregs\[26\]\[23\] cpuregs\[27\]\[23\]
+ _03516_ _03409_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__mux4_1
X_07999_ _02604_ _02606_ _02603_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__a21o_1
X_09738_ cpuregs\[20\]\[21\] cpuregs\[21\]\[21\] cpuregs\[22\]\[21\] cpuregs\[23\]\[21\]
+ _03438_ _03812_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_19_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09669_ _03807_ _04124_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_879 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _05495_ _05255_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_159_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ cpuregs\[12\]\[28\] cpuregs\[13\]\[28\] cpuregs\[14\]\[28\] cpuregs\[15\]\[28\]
+ _03133_ _03134_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11631_ decoded_imm_j\[20\] _05242_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14350_ _01802_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11562_ _05442_ _05444_ _05445_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13301_ _06804_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__clkbuf_1
X_10513_ _04738_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__clkbuf_1
X_14281_ net592 VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11493_ _05258_ net677 _05343_ _05382_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_137_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13232_ _06763_ decoded_imm_j\[9\] _06733_ mem_rdata_q\[29\] _06541_ VGND VGND VPWR
+ VPWR _06766_ sky130_fd_sc_hd__a221o_1
X_10444_ net973 _03355_ _04695_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13163_ latched_rd\[0\] _06724_ _06725_ net437 VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__a22o_1
X_10375_ cpuregs\[28\]\[26\] _03355_ _04658_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12114_ _05815_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_150_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13094_ _06689_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12045_ _03034_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_53_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15804_ clknet_leaf_132_clk _01379_ VGND VGND VPWR VPWR cpuregs\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_13996_ cpuregs\[5\]\[13\] _06952_ _01613_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__mux2_1
X_15735_ clknet_leaf_128_clk _01310_ VGND VGND VPWR VPWR cpuregs\[22\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_87_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12947_ _06608_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__buf_1
X_15666_ clknet_leaf_3_clk _01241_ VGND VGND VPWR VPWR cpuregs\[29\]\[19\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_160 _03193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12878_ is_alu_reg_reg _06528_ _06544_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__and3_1
*XANTENNA_171 _03552_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_182 _05113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_890 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14617_ clknet_leaf_1_clk _00275_ VGND VGND VPWR VPWR cpuregs\[21\]\[15\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_193 reg_next_pc\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11829_ _05664_ _05625_ _05665_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__and3b_1
X_15597_ clknet_leaf_143_clk _01172_ VGND VGND VPWR VPWR cpuregs\[31\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_16_618 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14548_ clknet_leaf_8_clk _00206_ VGND VGND VPWR VPWR cpuregs\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_491 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14479_ clknet_leaf_43_clk _00137_ VGND VGND VPWR VPWR cpuregs\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08971_ _03400_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__clkbuf_8
X_07922_ _02537_ _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__nor2_1
X_07853_ _02467_ _02470_ _02472_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__or3_1
X_07784_ _02398_ _02402_ _02403_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_88_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09523_ _03982_ _03983_ _03447_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__mux2_1
X_09454_ cpuregs\[12\]\[12\] cpuregs\[13\]\[12\] cpuregs\[14\]\[12\] cpuregs\[15\]\[12\]
+ _03582_ _03716_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_84_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08405_ reg_next_pc\[7\] reg_out\[7\] _02949_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__mux2_1
X_09385_ _03426_ _03845_ _03847_ _03849_ _03430_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_19_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08336_ _02920_ _02922_ _02393_ _02924_ VGND VGND VPWR VPWR alu_out\[31\] sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_148_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_798 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_642 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08267_ net246 _02850_ _02757_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_140_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_140_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07218_ net673 _01874_ _01876_ _01880_ _01881_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08198_ net215 _02797_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_678 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07149_ mem_do_rdata _01816_ _01817_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ _04550_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__clkbuf_1
X_10091_ _04512_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13850_ cpuregs\[22\]\[9\] _06943_ _07100_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12801_ _05289_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__buf_4
X_10993_ cpuregs\[17\]\[12\] _04844_ _05006_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__mux2_1
X_13781_ _07073_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15520_ clknet_leaf_160_clk _01105_ VGND VGND VPWR VPWR cpuregs\[24\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12732_ cpuregs\[28\]\[30\] cpuregs\[29\]\[30\] _05895_ VGND VGND VPWR VPWR _06472_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15451_ clknet_leaf_159_clk _01041_ VGND VGND VPWR VPWR cpuregs\[19\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ cpuregs\[31\]\[27\] _05974_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__or2b_1
XFILLER_0_139_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14402_ clknet_leaf_135_clk _00065_ VGND VGND VPWR VPWR cpuregs\[11\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11614_ _05418_ net493 _05343_ _05493_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_871 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15382_ clknet_leaf_89_clk _00972_ VGND VGND VPWR VPWR decoded_imm\[26\] sky130_fd_sc_hd__dfxtp_4
X_12594_ _03132_ _06339_ _05840_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14333_ _01793_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__clkbuf_1
X_11545_ _05222_ _05429_ _05225_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_131_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_131_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_152_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14264_ _01757_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__clkbuf_1
X_11476_ _05288_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10427_ net908 _03302_ _04684_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__mux2_1
X_13215_ decoded_imm\[17\] _06752_ _06735_ _06756_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__o22a_1
X_14195_ _01722_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__clkbuf_1
X_13146_ _06716_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__clkbuf_1
X_10358_ cpuregs\[28\]\[18\] _03302_ _04647_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13077_ mem_do_rdata _01816_ _06674_ _06677_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__o31ai_1
X_10289_ _04619_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12028_ _05800_ _01877_ _01890_ _05801_ _01860_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__o311a_1
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13979_ cpuregs\[5\]\[5\] _06935_ _01602_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__mux2_1
X_15718_ clknet_leaf_36_clk _01293_ VGND VGND VPWR VPWR cpuregs\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_66_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15649_ clknet_leaf_25_clk _01224_ VGND VGND VPWR VPWR cpuregs\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_726 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_56_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09170_ _03640_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__buf_8
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_404 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_521 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_83_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08121_ _02471_ _02463_ _02701_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_32_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_122_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_122_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08052_ _02646_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpicorv32_264 VGND VGND VPWR VPWR picorv32_264/HI eoi[10] sky130_fd_sc_hd__conb_1
Xpicorv32_275 VGND VGND VPWR VPWR picorv32_275/HI eoi[21] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_114_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_286 VGND VGND VPWR VPWR picorv32_286/HI mem_addr[0] sky130_fd_sc_hd__conb_1
Xpicorv32_297 VGND VGND VPWR VPWR picorv32_297/HI pcpi_insn[7] sky130_fd_sc_hd__conb_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08954_ _00016_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__inv_4
X_07905_ _02482_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__inv_2
X_08885_ reg_pc\[28\] reg_pc\[27\] _03352_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07836_ _02451_ _02455_ _02435_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__a21oi_1
X_07767_ count_cycle\[31\] _02051_ _02387_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__a21o_1
X_09506_ _03963_ _03965_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__or2_1
X_07698_ count_cycle\[26\] _02051_ _02322_ _02323_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_698 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09437_ decoded_imm\[10\] net172 _03863_ _03899_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_149_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09368_ decoded_imm\[10\] net172 VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08319_ net226 _02908_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_10_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_113_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_113_clk sky130_fd_sc_hd__clkbuf_2
X_09299_ _03734_ _03738_ _03735_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_60 _03500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_71 _03637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_82 _04844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ reg_next_pc\[22\] _03324_ _02947_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_134_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_93 _05886_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11261_ _05190_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__buf_2
X_10212_ net857 _03268_ _04575_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__mux2_1
X_13000_ net583 _04817_ _06636_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__mux2_1
X_11192_ net513 net382 _05142_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__a21oi_1
X_10143_ _04541_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14951_ clknet_leaf_115_clk _00609_ VGND VGND VPWR VPWR count_instr\[60\] sky130_fd_sc_hd__dfxtp_1
X_10074_ _04503_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_1
X_13902_ _01567_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__clkbuf_1
X_14882_ clknet_leaf_125_clk _00540_ VGND VGND VPWR VPWR cpuregs\[17\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_13833_ _07101_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_134_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13764_ net609 _06923_ _07064_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__mux2_1
X_10976_ net941 _04827_ _04995_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15503_ clknet_leaf_85_clk _01088_ VGND VGND VPWR VPWR mem_rdata_q\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12715_ net224 _06455_ _06282_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__mux2_1
X_13695_ _07027_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15434_ clknet_leaf_150_clk _01024_ VGND VGND VPWR VPWR cpuregs\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_12646_ _05886_ _06379_ _06383_ _05978_ _06389_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__a311o_2
XFILLER_0_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_104_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_104_clk sky130_fd_sc_hd__clkbuf_2
X_15365_ clknet_leaf_69_clk _00955_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dfxtp_1
X_12577_ cpuregs\[24\]\[23\] cpuregs\[25\]\[23\] cpuregs\[26\]\[23\] cpuregs\[27\]\[23\]
+ _06074_ _03151_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14316_ _01784_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__clkbuf_1
X_11528_ _01890_ _05414_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15296_ clknet_leaf_48_clk _00886_ VGND VGND VPWR VPWR cpuregs\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold308 cpuregs\[27\]\[12\] VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold319 cpuregs\[11\]\[16\] VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ net605 VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__clkbuf_1
X_11459_ _05323_ _05335_ _05350_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__nand3_1
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14178_ _01713_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13129_ net147 net109 _06707_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1008 cpuregs\[15\]\[21\] VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 cpuregs\[16\]\[16\] VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08670_ reg_out\[0\] alu_out_q\[0\] _03176_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07621_ net13 _02252_ _02180_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07552_ count_instr\[47\] _02013_ _02017_ _02188_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07483_ _01945_ _02122_ _02123_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09222_ _03685_ _03687_ _03689_ _03691_ _03431_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__a221o_2
XFILLER_0_17_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09153_ _03486_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08104_ _02706_ _02711_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__nand2_1
X_09084_ _00014_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08035_ _02646_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold820 cpuregs\[24\]\[9\] VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_626 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold831 cpuregs\[21\]\[25\] VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold842 cpuregs\[24\]\[7\] VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 cpuregs\[29\]\[17\] VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 cpuregs\[14\]\[31\] VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold875 cpuregs\[9\]\[28\] VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 cpuregs\[14\]\[6\] VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold897 cpuregs\[6\]\[16\] VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09986_ cpuregs\[8\]\[29\] cpuregs\[9\]\[29\] cpuregs\[10\]\[29\] cpuregs\[11\]\[29\]
+ _03548_ _03449_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__mux4_1
X_08937_ _03403_ _03411_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08868_ _03349_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__clkbuf_1
X_07819_ net253 net223 VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__and2_1
X_08799_ reg_out\[17\] alu_out_q\[17\] _03175_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__mux2_1
X_10830_ _04562_ _04744_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__nor2_4
XFILLER_0_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10761_ latched_rd\[3\] latched_rd\[2\] latched_rd\[4\] VGND VGND VPWR VPWR _04885_
+ sky130_fd_sc_hd__or3b_4
X_12500_ cpuregs\[8\]\[20\] cpuregs\[9\]\[20\] cpuregs\[10\]\[20\] cpuregs\[11\]\[20\]
+ _06061_ _03137_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_167 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13480_ _06887_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__buf_4
X_10692_ _04838_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12431_ cpuregs\[8\]\[17\] cpuregs\[9\]\[17\] cpuregs\[10\]\[17\] cpuregs\[11\]\[17\]
+ _06061_ _05917_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15150_ clknet_leaf_69_clk _00775_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
X_12362_ _05969_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14101_ net1156 _06989_ _01637_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__mux2_1
X_11313_ reg_next_pc\[17\] _03289_ _02947_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__mux2_2
X_15081_ clknet_leaf_92_clk _00739_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dfxtp_1
X_12293_ _05862_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__clkbuf_4
X_11244_ count_instr\[61\] count_instr\[60\] _05175_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__and3_1
X_14032_ _01635_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11175_ net536 _05128_ _05090_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__o21ai_1
X_10126_ _04532_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14934_ clknet_leaf_121_clk _00592_ VGND VGND VPWR VPWR count_instr\[43\] sky130_fd_sc_hd__dfxtp_1
X_10057_ _04494_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_1
X_14865_ clknet_leaf_26_clk _00523_ VGND VGND VPWR VPWR cpuregs\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13816_ net1120 _06977_ _07086_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14796_ clknet_leaf_27_clk _00454_ VGND VGND VPWR VPWR cpuregs\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13747_ _07055_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_63_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10959_ _04990_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13678_ net706 _06975_ _07014_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15417_ clknet_leaf_29_clk _01007_ VGND VGND VPWR VPWR cpuregs\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_852 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12629_ cpuregs\[12\]\[26\] cpuregs\[13\]\[26\] cpuregs\[14\]\[26\] cpuregs\[15\]\[26\]
+ _05834_ _03129_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15348_ clknet_leaf_68_clk _00938_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold105 instr_and VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 count_instr\[60\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ clknet_leaf_99_clk _00872_ VGND VGND VPWR VPWR decoded_imm_j\[16\] sky130_fd_sc_hd__dfxtp_2
Xhold127 cpuregs\[0\]\[15\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 reg_next_pc\[29\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 count_cycle\[4\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_793 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09840_ _04289_ _04290_ _03455_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ cpuregs\[28\]\[22\] cpuregs\[29\]\[22\] cpuregs\[30\]\[22\] cpuregs\[31\]\[22\]
+ _03463_ _03460_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__mux4_1
X_08722_ _03222_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08653_ decoded_imm_j\[2\] _01084_ _03022_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07604_ net181 VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08584_ _03081_ _03089_ _03094_ _03100_ _03102_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__o32a_1
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07535_ reg_pc\[15\] decoded_imm\[15\] VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07466_ reg_pc\[9\] decoded_imm\[9\] VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_45_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09205_ cpuregs\[4\]\[5\] cpuregs\[5\]\[5\] cpuregs\[6\]\[5\] cpuregs\[7\]\[5\] _03673_
+ _03674_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07397_ _02040_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09136_ _03574_ _03592_ _03607_ _03526_ reg_pc\[3\] VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09067_ decoded_imm\[2\] net193 VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_710 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_570 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08018_ _02492_ _02631_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__xnor2_1
Xhold650 cpuregs\[9\]\[20\] VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 cpuregs\[13\]\[0\] VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 cpuregs\[9\]\[30\] VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 cpuregs\[4\]\[17\] VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 cpuregs\[1\]\[17\] VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__dlygate4sd3_1
X_09969_ _03500_ _04415_ _03427_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_129_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ decoded_imm_j\[3\] _01085_ _03021_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__mux2_1
X_11931_ cpuregs\[8\]\[31\] cpuregs\[9\]\[31\] cpuregs\[10\]\[31\] cpuregs\[11\]\[31\]
+ _03582_ _03716_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_142_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ clknet_leaf_10_clk _00308_ VGND VGND VPWR VPWR cpuregs\[14\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11862_ count_cycle\[43\] net360 _05622_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__o21ai_1
X_13601_ _06974_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__clkbuf_1
X_10813_ _04913_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_45_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ clknet_leaf_2_clk _00239_ VGND VGND VPWR VPWR cpuregs\[28\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11793_ count_cycle\[21\] _05637_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13532_ cpuregs\[31\]\[1\] _06927_ _06925_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__mux2_1
X_10744_ net913 _04873_ _04861_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13463_ _06890_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10675_ _03208_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__buf_2
XFILLER_0_125_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15202_ clknet_leaf_65_clk alu_out\[15\] VGND VGND VPWR VPWR alu_out_q\[15\] sky130_fd_sc_hd__dfxtp_1
X_12414_ cpuregs\[16\]\[16\] cpuregs\[17\]\[16\] cpuregs\[18\]\[16\] cpuregs\[19\]\[16\]
+ _05948_ _06068_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13394_ net716 _04821_ _06852_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15133_ clknet_leaf_111_clk _00759_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_389 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12345_ _06098_ _06100_ _06101_ _03132_ _05815_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15064_ clknet_leaf_121_clk _00722_ VGND VGND VPWR VPWR count_cycle\[47\] sky130_fd_sc_hd__dfxtp_1
X_12276_ cpuregs\[0\]\[11\] cpuregs\[1\]\[11\] cpuregs\[2\]\[11\] cpuregs\[3\]\[11\]
+ _05908_ _05909_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__mux4_1
X_14015_ net1163 _06971_ _01624_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__mux2_1
X_11227_ _05165_ _05113_ _05166_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_56_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11158_ net595 net375 _05118_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_8_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10109_ _04521_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__clkbuf_1
X_11089_ count_instr\[13\] count_instr\[12\] VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__and2_1
X_15966_ clknet_leaf_135_clk _01538_ VGND VGND VPWR VPWR cpuregs\[10\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_14917_ clknet_leaf_117_clk _00575_ VGND VGND VPWR VPWR count_instr\[26\] sky130_fd_sc_hd__dfxtp_1
X_15897_ clknet_leaf_140_clk _01469_ VGND VGND VPWR VPWR cpuregs\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14848_ clknet_leaf_146_clk _00506_ VGND VGND VPWR VPWR cpuregs\[20\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14779_ clknet_leaf_158_clk _00437_ VGND VGND VPWR VPWR cpuregs\[16\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_07320_ cpu_state\[3\] VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_424 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07251_ is_sll_srl_sra is_lb_lh_lw_lbu_lhu is_sb_sh_sw _01908_ VGND VGND VPWR VPWR
+ _01909_ sky130_fd_sc_hd__or4_1
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07182_ mem_wordsize\[2\] VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__buf_4
XFILLER_0_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09823_ decoded_imm\[24\] net187 VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__or2_1
X_09754_ _02265_ _04207_ _03395_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__mux2_1
X_08705_ _03173_ _03204_ _03205_ _03207_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__a22o_2
X_09685_ _01953_ _04138_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_93_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_124_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ cpuregs\[28\]\[4\] cpuregs\[29\]\[4\] cpuregs\[30\]\[4\] cpuregs\[31\]\[4\]
+ _03062_ _03063_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__mux4_1
X_08567_ _03039_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07518_ _02065_ _02154_ _02156_ _01927_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_540 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_49_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08498_ _03025_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07449_ count_instr\[41\] _02052_ _02055_ count_cycle\[41\] VGND VGND VPWR VPWR _02092_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_548 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_885 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10460_ net1097 _03189_ _04709_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09119_ _03489_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__buf_4
XFILLER_0_115_570 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10391_ _04674_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12130_ _03062_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__buf_6
XFILLER_0_130_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12061_ _03124_ _05830_ _03034_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold480 net195 VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 cpuregs\[19\]\[22\] VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ net762 _04863_ _05017_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__mux2_1
X_15820_ clknet_leaf_8_clk _01392_ VGND VGND VPWR VPWR cpuregs\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ clknet_leaf_57_clk _01326_ VGND VGND VPWR VPWR cpuregs\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12963_ _06616_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_84_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_2
X_14702_ clknet_leaf_44_clk _00360_ VGND VGND VPWR VPWR cpuregs\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11914_ count_cycle\[59\] _05706_ _05713_ _05720_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__and4_1
XFILLER_0_158_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15682_ clknet_leaf_39_clk _01257_ VGND VGND VPWR VPWR cpuregs\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12894_ _06555_ _06577_ _06578_ _06579_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14633_ clknet_leaf_19_clk _00291_ VGND VGND VPWR VPWR cpuregs\[21\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11845_ _05675_ _05625_ _05676_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__and3b_1
XFILLER_0_142_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14564_ clknet_leaf_17_clk _00222_ VGND VGND VPWR VPWR cpuregs\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11776_ _05628_ _05629_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13515_ _06917_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_906 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10727_ _04862_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__clkbuf_1
X_14495_ clknet_leaf_130_clk _00153_ VGND VGND VPWR VPWR cpuregs\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13446_ net979 _04873_ _06874_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10658_ _04815_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13377_ _06844_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10589_ net694 _03381_ _04745_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15116_ clknet_leaf_74_clk _00742_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_1
X_12328_ _06081_ _06083_ _06084_ _03128_ _03035_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15047_ clknet_leaf_114_clk _00705_ VGND VGND VPWR VPWR count_cycle\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12259_ _03106_ _06018_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15949_ clknet_leaf_8_clk _01521_ VGND VGND VPWR VPWR cpuregs\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_75_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_2
X_09470_ _03894_ _03902_ _03930_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08421_ _02972_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08352_ _02463_ _02927_ _02932_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__a21o_1
XFILLER_0_19_638 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07303_ _01954_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__buf_4
X_08283_ _02331_ net221 _02618_ _02562_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_427 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07234_ _01893_ is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07165_ instr_ori instr_xori instr_addi instr_bltu VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_793 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_560 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09806_ _03448_ _04257_ _03419_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07998_ _02612_ _02613_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__and2_1
X_09737_ _03547_ _04186_ _04188_ _04190_ _00016_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__a221o_1
X_09668_ cpuregs\[12\]\[19\] cpuregs\[13\]\[19\] cpuregs\[14\]\[19\] cpuregs\[15\]\[19\]
+ _03438_ _03549_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_159_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _03052_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_159_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _04054_ _04055_ _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_139_459 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11630_ decoded_imm_j\[20\] _05242_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11561_ decoded_imm_j\[17\] _05228_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13300_ cpuregs\[18\]\[21\] _04863_ _06802_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__mux2_1
X_10512_ net836 _03355_ _04731_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__mux2_1
X_14280_ _01765_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__clkbuf_1
X_11492_ _05375_ _05376_ _05381_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_137_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_613 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13231_ decoded_imm\[10\] _06626_ _06765_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__o21a_1
X_10443_ _04701_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_32_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13162_ _02058_ _06724_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10374_ _04664_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__clkbuf_1
X_12113_ cpuregs\[16\]\[5\] cpuregs\[17\]\[5\] cpuregs\[18\]\[5\] cpuregs\[19\]\[5\]
+ _03096_ _03098_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_150_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13093_ net160 net251 _06685_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__mux2_1
X_12044_ decoded_imm\[0\] _01906_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_53_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15803_ clknet_leaf_130_clk _01378_ VGND VGND VPWR VPWR cpuregs\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13995_ _01616_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_57_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_2
X_15734_ clknet_leaf_146_clk _01309_ VGND VGND VPWR VPWR cpuregs\[22\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ mem_rdata_q\[7\] net30 _06589_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_87_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15665_ clknet_leaf_154_clk _01240_ VGND VGND VPWR VPWR cpuregs\[29\]\[18\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_150 _01869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12877_ _05041_ _06543_ _06568_ _06562_ net615 VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__a32o_1
XFILLER_0_158_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_161 _03220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14616_ clknet_leaf_153_clk _00274_ VGND VGND VPWR VPWR cpuregs\[21\]\[14\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_172 _03557_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11828_ count_cycle\[31\] net364 count_cycle\[32\] VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__a21o_1
*XANTENNA_183 _05113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15596_ clknet_leaf_154_clk _01171_ VGND VGND VPWR VPWR cpuregs\[31\]\[13\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_194 reg_next_pc\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14547_ clknet_leaf_31_clk _00205_ VGND VGND VPWR VPWR cpuregs\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11759_ net531 count_cycle\[11\] _05613_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14478_ clknet_leaf_45_clk _00136_ VGND VGND VPWR VPWR cpuregs\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13429_ net915 _04856_ _06863_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08970_ _03437_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__or2_1
X_16079_ net119 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_2
X_07921_ _02538_ _02539_ _02540_ _02408_ _02448_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__a2111o_1
X_07852_ net175 _02471_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__xor2_1
Xinput1 net412 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_07783_ _02277_ net217 VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_88_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_48_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_88_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09522_ cpuregs\[0\]\[14\] cpuregs\[1\]\[14\] cpuregs\[2\]\[14\] cpuregs\[3\]\[14\]
+ _03457_ _03595_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_104_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_847 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09453_ _03433_ _03911_ _03913_ _03915_ _03760_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08404_ _02960_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_1
XFILLER_0_47_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09384_ _03401_ _03848_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08335_ _02392_ _02581_ _02923_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_930 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08266_ _02428_ _02569_ _02860_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_641 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07217_ instr_lbu instr_lb _01866_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__o21a_1
X_08197_ net213 _02791_ _02656_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07148_ mem_state\[1\] mem_state\[0\] VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ net1222 _03329_ _04509_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_2
X_12800_ net438 _06513_ _06519_ _06524_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__a22o_1
X_13780_ net962 _06941_ _07064_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__mux2_1
X_10992_ _05008_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__clkbuf_1
X_12731_ _05974_ cpuregs\[30\]\[30\] _05896_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__o21a_1
X_15450_ clknet_leaf_158_clk _01040_ VGND VGND VPWR VPWR cpuregs\[19\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_12662_ _05969_ _06404_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ clknet_leaf_20_clk _00064_ VGND VGND VPWR VPWR cpuregs\[11\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11613_ _05263_ _05492_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__nand2_1
X_15381_ clknet_leaf_89_clk _00971_ VGND VGND VPWR VPWR decoded_imm\[27\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_148_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12593_ cpuregs\[16\]\[24\] cpuregs\[17\]\[24\] cpuregs\[18\]\[24\] cpuregs\[19\]\[24\]
+ _05984_ _06068_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ net904 _03267_ _01789_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11544_ _05217_ _05219_ _05387_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14263_ net666 VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11475_ _05032_ _05365_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__nand2_1
X_13214_ _06525_ net510 _06738_ mem_rdata_q\[17\] VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__a22o_1
X_10426_ _04692_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14194_ net745 _06945_ _01721_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13145_ net1229 net117 _06707_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__mux2_1
X_10357_ _04655_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13076_ _01817_ _01855_ _01857_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__or3_1
X_10288_ net899 _03295_ _04611_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__mux2_1
X_12027_ _01878_ _01903_ mem_do_prefetch VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__a21o_1
X_13978_ _01607_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__clkbuf_1
X_12929_ _06599_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
X_15717_ clknet_leaf_30_clk _01292_ VGND VGND VPWR VPWR cpuregs\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_519 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15648_ clknet_leaf_52_clk _01223_ VGND VGND VPWR VPWR cpuregs\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15579_ clknet_leaf_135_clk _01154_ VGND VGND VPWR VPWR cpuregs\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_894 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08120_ _02608_ _02722_ _02723_ _02726_ VGND VGND VPWR VPWR alu_out\[13\] sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_32_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08051_ _02635_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_254 VGND VGND VPWR VPWR picorv32_254/HI eoi[0] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_114_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_265 VGND VGND VPWR VPWR picorv32_265/HI eoi[11] sky130_fd_sc_hd__conb_1
Xpicorv32_276 VGND VGND VPWR VPWR picorv32_276/HI eoi[22] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_114_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_287 VGND VGND VPWR VPWR picorv32_287/HI mem_addr[1] sky130_fd_sc_hd__conb_1
Xpicorv32_298 VGND VGND VPWR VPWR picorv32_298/HI pcpi_insn[8] sky130_fd_sc_hd__conb_1
X_08953_ _03415_ _03424_ _03427_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07904_ _02066_ _02490_ _02501_ _02517_ _02523_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__o221a_1
X_08884_ reg_pc\[27\] _03352_ reg_pc\[28\] VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07835_ _02426_ _02427_ _02452_ _02454_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__a22o_1
X_07766_ count_instr\[63\] _02013_ _02017_ _02386_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_655 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09505_ _03963_ _03965_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_817 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07697_ count_instr\[26\] _02054_ count_cycle\[58\] _02055_ VGND VGND VPWR VPWR _02323_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _03795_ _03830_ _03896_ net173 decoded_imm\[11\] VGND VGND VPWR VPWR _03899_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_137_705 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09367_ decoded_imm\[10\] net172 VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08318_ _02757_ net224 _02900_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_10_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09298_ decoded_imm\[8\] net201 VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__xnor2_1
*XANTENNA_50 _03402_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_61 _03516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_72 _03673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_83 _04846_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08249_ net186 _02837_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_134_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_94 _05921_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11260_ reg_next_pc\[2\] _03192_ _02945_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__mux2_1
X_10211_ _04578_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__clkbuf_1
X_11191_ net1400 net382 _05141_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__o21ai_1
X_10142_ cpuregs\[30\]\[13\] _03268_ _04537_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput190 net190 VGND VGND VPWR VPWR pcpi_rs1[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ clknet_leaf_115_clk _00608_ VGND VGND VPWR VPWR count_instr\[59\] sky130_fd_sc_hd__dfxtp_1
X_10073_ cpuregs\[12\]\[14\] _03275_ _04498_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__mux2_1
X_13901_ net897 _06923_ _01566_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__mux2_1
X_14881_ clknet_leaf_148_clk _00539_ VGND VGND VPWR VPWR cpuregs\[17\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_13832_ net1346 _06923_ _07100_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13763_ _07063_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__buf_6
X_10975_ _04999_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12714_ _05900_ _06445_ _06454_ _01918_ decoded_imm\[29\] VGND VGND VPWR VPWR _06455_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_84_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15502_ clknet_leaf_82_clk _01087_ VGND VGND VPWR VPWR mem_rdata_q\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_198 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13694_ _04522_ _04562_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__nor2_4
XFILLER_0_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15433_ clknet_leaf_125_clk _01023_ VGND VGND VPWR VPWR cpuregs\[18\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12645_ _06385_ _06387_ _06388_ _03149_ _05815_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_26_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_259 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15364_ clknet_leaf_69_clk _00954_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dfxtp_1
X_12576_ _06026_ _06322_ _06193_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_61_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14315_ net1026 _03214_ _01778_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11527_ _05215_ _05413_ _05380_ _05219_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__or4b_2
XFILLER_0_124_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15295_ clknet_leaf_78_clk _00885_ VGND VGND VPWR VPWR is_beq_bne_blt_bge_bltu_bgeu
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_151_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_22_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold309 cpuregs\[0\]\[27\] VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__dlygate4sd3_1
X_14246_ _01748_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11458_ decoded_imm_j\[5\] _05199_ _05314_ _05313_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10409_ _04683_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__clkbuf_1
X_14177_ cpuregs\[8\]\[2\] _06929_ _01710_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__mux2_1
X_11389_ _05269_ _05279_ _05281_ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__a31o_1
X_13128_ _06684_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__clkbuf_4
X_13059_ _06667_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__clkbuf_1
Xhold1009 cpuregs\[6\]\[17\] VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07620_ _02251_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07551_ count_instr\[15\] _01949_ count_cycle\[47\] _02014_ VGND VGND VPWR VPWR _02188_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07482_ _02105_ _02111_ _02121_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__or3_1
XFILLER_0_76_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09221_ _03437_ _03690_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09152_ _03623_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08103_ _02709_ _02710_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_116_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09083_ _03401_ _03555_ _03418_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08034_ net200 _02645_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold810 cpuregs\[5\]\[7\] VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold821 cpuregs\[21\]\[16\] VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 cpuregs\[29\]\[12\] VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold843 cpuregs\[19\]\[20\] VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 cpuregs\[28\]\[22\] VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold865 cpuregs\[19\]\[19\] VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 cpuregs\[9\]\[21\] VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 cpuregs\[4\]\[9\] VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_660 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold898 cpuregs\[6\]\[6\] VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _04429_ _04430_ _03552_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08936_ cpuregs\[12\]\[0\] cpuregs\[13\]\[0\] cpuregs\[14\]\[0\] cpuregs\[15\]\[0\]
+ _03406_ _03410_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__mux4_1
X_08867_ net783 _03348_ _03315_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07818_ net253 net223 VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08798_ _03288_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_64_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07749_ _01945_ _02368_ _02371_ _01968_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10760_ _04884_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09419_ cpuregs\[24\]\[11\] cpuregs\[25\]\[11\] cpuregs\[26\]\[11\] cpuregs\[27\]\[11\]
+ _03516_ _03409_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10691_ net1030 _04837_ _04819_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12430_ _06058_ _06181_ _06182_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12361_ cpuregs\[24\]\[14\] cpuregs\[25\]\[14\] cpuregs\[26\]\[14\] cpuregs\[27\]\[14\]
+ _05970_ _03108_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14100_ _01671_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11312_ _05184_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__buf_2
X_15080_ clknet_leaf_115_clk _00738_ VGND VGND VPWR VPWR count_cycle\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_914 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12292_ _05901_ _06041_ _06050_ _05904_ decoded_imm\[11\] VGND VGND VPWR VPWR _06051_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14031_ cpuregs\[5\]\[30\] _06987_ _01601_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__mux2_1
X_11243_ net475 _05175_ _05177_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__a21oi_1
X_11174_ count_instr\[39\] count_instr\[38\] net373 VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__and3_1
X_10125_ cpuregs\[30\]\[5\] _03215_ _04526_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14933_ clknet_leaf_121_clk _00591_ VGND VGND VPWR VPWR count_instr\[42\] sky130_fd_sc_hd__dfxtp_1
X_10056_ net1017 _03221_ _04487_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14864_ clknet_leaf_27_clk _00522_ VGND VGND VPWR VPWR cpuregs\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_901 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13815_ _07091_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14795_ clknet_leaf_46_clk _00453_ VGND VGND VPWR VPWR cpuregs\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13746_ net743 _06975_ _07050_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10958_ net803 _04877_ _04981_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_513 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13677_ _07018_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10889_ _04953_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12628_ _06368_ _06370_ _06371_ _03128_ _03035_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__o221a_1
X_15416_ clknet_leaf_25_clk _01006_ VGND VGND VPWR VPWR cpuregs\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15347_ clknet_leaf_69_clk _00937_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12559_ _05886_ _06296_ _06300_ _05978_ _06306_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__a311o_1
XFILLER_0_53_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_91_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold106 count_instr\[17\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15278_ clknet_leaf_95_clk _00871_ VGND VGND VPWR VPWR decoded_imm_j\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold117 count_cycle\[57\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_569 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_111_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold128 count_cycle\[27\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 count_instr\[59\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ cpuregs\[8\]\[27\] _06981_ _01732_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09770_ _03746_ _04222_ _03419_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_91_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ cpuregs\[11\]\[6\] _03221_ _03185_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08652_ _03164_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__buf_1
XFILLER_0_89_750 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ _02234_ _02235_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08583_ _03083_ _03101_ _03081_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_647 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07534_ _01970_ _02164_ _02171_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07465_ _02106_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09204_ _03576_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__buf_6
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07396_ _02038_ _02041_ _01945_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_161_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09135_ _03597_ _03600_ _03604_ _03606_ _03430_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09066_ _03398_ _03530_ _03538_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08017_ _02609_ _02630_ _02573_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_295 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold640 cpuregs\[6\]\[23\] VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 cpuregs\[13\]\[15\] VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 cpuregs\[30\]\[12\] VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 cpuregs\[6\]\[20\] VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 reg_next_pc\[10\] VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold695 cpuregs\[7\]\[8\] VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__dlygate4sd3_1
X_09968_ cpuregs\[16\]\[28\] cpuregs\[17\]\[28\] cpuregs\[18\]\[28\] cpuregs\[19\]\[28\]
+ _03641_ _03642_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_129_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _03388_ _01864_ _03393_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09899_ cpuregs\[28\]\[26\] cpuregs\[29\]\[26\] cpuregs\[30\]\[26\] cpuregs\[31\]\[26\]
+ _03463_ _03464_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__mux4_1
X_11930_ _05733_ _05734_ _03401_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _05686_ _05687_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_142_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ net952 _06973_ _06967_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10812_ cpuregs\[16\]\[23\] _04867_ _04909_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__mux2_1
X_14580_ clknet_leaf_2_clk _00238_ VGND VGND VPWR VPWR cpuregs\[28\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11792_ count_cycle\[19\] count_cycle\[20\] count_cycle\[21\] _05634_ VGND VGND VPWR
+ VPWR _05640_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_45_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _03188_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10743_ _03354_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13462_ net1045 _04821_ _06888_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__mux2_1
X_10674_ _04826_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__clkbuf_1
X_15201_ clknet_leaf_71_clk alu_out\[14\] VGND VGND VPWR VPWR alu_out_q\[14\] sky130_fd_sc_hd__dfxtp_1
X_12413_ _06142_ _06166_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_106_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13393_ _06853_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15132_ clknet_leaf_108_clk _00758_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12344_ cpuregs\[16\]\[13\] cpuregs\[17\]\[13\] cpuregs\[18\]\[13\] cpuregs\[19\]\[13\]
+ _05984_ _05985_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15063_ clknet_leaf_132_clk _00721_ VGND VGND VPWR VPWR count_cycle\[46\] sky130_fd_sc_hd__dfxtp_1
X_12275_ cpuregs\[4\]\[11\] cpuregs\[5\]\[11\] cpuregs\[6\]\[11\] cpuregs\[7\]\[11\]
+ _06011_ _03097_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__mux4_1
X_14014_ _01626_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__clkbuf_1
X_11226_ count_instr\[54\] _05162_ count_instr\[55\] VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_56_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11157_ count_instr\[34\] net386 _05036_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ net777 _03386_ _04486_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__mux2_1
X_11088_ net467 VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__inv_2
X_15965_ clknet_leaf_20_clk _01537_ VGND VGND VPWR VPWR cpuregs\[10\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_14916_ clknet_leaf_118_clk _00574_ VGND VGND VPWR VPWR count_instr\[25\] sky130_fd_sc_hd__dfxtp_1
X_10039_ latched_rd\[3\] latched_rd\[4\] latched_rd\[2\] VGND VGND VPWR VPWR _04483_
+ sky130_fd_sc_hd__or3_4
X_15896_ clknet_leaf_141_clk _01468_ VGND VGND VPWR VPWR cpuregs\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_14847_ clknet_leaf_124_clk _00505_ VGND VGND VPWR VPWR cpuregs\[20\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14778_ clknet_leaf_158_clk _00436_ VGND VGND VPWR VPWR cpuregs\[16\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_86_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13729_ net949 _06958_ _07039_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07250_ _01907_ _01838_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__or2b_1
XFILLER_0_156_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_54_661 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07181_ net171 VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09822_ decoded_imm\[24\] _02306_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__nand2_1
X_09753_ _03651_ _04182_ _04183_ _04202_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__a311o_1
X_08704_ _03172_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__nor2_1
X_09684_ _04029_ _04139_ _03657_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08635_ _03037_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_539 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08566_ _03084_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__buf_8
XFILLER_0_65_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07517_ _02083_ _02155_ _02085_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_138_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08497_ decoded_imm_j\[16\] _01078_ _03022_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07448_ _02091_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_650 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07379_ _02024_ _02025_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09118_ _03447_ _03589_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__or2_1
X_10390_ net976 _03179_ _04673_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09049_ _03490_ _03502_ _03508_ _03514_ _03522_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__a32o_1
X_12060_ cpuregs\[20\]\[0\] cpuregs\[21\]\[0\] cpuregs\[22\]\[0\] cpuregs\[23\]\[0\]
+ _03091_ _05829_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__mux4_1
Xhold470 cpuregs\[17\]\[22\] VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 cpuregs\[29\]\[11\] VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ _05018_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__clkbuf_1
Xhold492 cpuregs\[21\]\[6\] VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ mem_rdata_q\[11\] net3 _03018_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__mux2_1
X_15750_ clknet_leaf_34_clk _01325_ VGND VGND VPWR VPWR cpuregs\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11913_ _05723_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__clkbuf_1
X_14701_ clknet_leaf_39_clk _00359_ VGND VGND VPWR VPWR cpuregs\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12893_ mem_rdata_q\[17\] mem_rdata_q\[16\] mem_rdata_q\[15\] VGND VGND VPWR VPWR
+ _06579_ sky130_fd_sc_hd__or3_1
X_15681_ clknet_leaf_26_clk _01256_ VGND VGND VPWR VPWR cpuregs\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11844_ count_cycle\[37\] _05673_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__or2_1
X_14632_ clknet_leaf_22_clk _00290_ VGND VGND VPWR VPWR cpuregs\[21\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14563_ clknet_leaf_134_clk _00221_ VGND VGND VPWR VPWR cpuregs\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11775_ net637 _05624_ _05169_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10726_ net1013 _04860_ _04861_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__mux2_1
X_13514_ net849 _04873_ _06910_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__mux2_1
X_14494_ clknet_leaf_146_clk _00152_ VGND VGND VPWR VPWR cpuregs\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13445_ _06880_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10657_ net786 _03381_ _04781_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_677 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_152_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13376_ cpuregs\[19\]\[25\] _04871_ _06838_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__mux2_1
X_10588_ _04778_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12327_ cpuregs\[0\]\[13\] cpuregs\[1\]\[13\] cpuregs\[2\]\[13\] cpuregs\[3\]\[13\]
+ _05819_ _03125_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__mux4_1
X_15115_ clknet_leaf_74_clk _00741_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15046_ clknet_leaf_120_clk _00704_ VGND VGND VPWR VPWR count_cycle\[29\] sky130_fd_sc_hd__dfxtp_1
X_12258_ cpuregs\[8\]\[10\] cpuregs\[9\]\[10\] cpuregs\[10\]\[10\] cpuregs\[11\]\[10\]
+ _03150_ _05917_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11209_ count_instr\[47\] _05146_ _05154_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__and3_1
X_12189_ _03083_ _05951_ _03081_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_71_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15948_ clknet_leaf_11_clk _01520_ VGND VGND VPWR VPWR cpuregs\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15879_ clknet_leaf_38_clk _01451_ VGND VGND VPWR VPWR cpuregs\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_08420_ _02125_ _02970_ _02971_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08351_ _01880_ net250 _02463_ _01913_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07302_ cpu_state\[3\] cpu_state\[6\] _01953_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_22_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_129_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08282_ _02871_ _02874_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07233_ cpu_state\[3\] VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07164_ instr_blt instr_bne instr_beq instr_rdcycle VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xfanout246 net219 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_161_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09805_ cpuregs\[28\]\[23\] cpuregs\[29\]\[23\] cpuregs\[30\]\[23\] cpuregs\[31\]\[23\]
+ _03680_ _03443_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__mux4_1
X_07997_ net197 _02611_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09736_ _03807_ _04189_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__or2_1
X_09667_ _03413_ _04122_ _03418_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08618_ _03132_ _03135_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_159_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _04054_ _04055_ _01870_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_159_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_241 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08549_ _03045_ _03066_ _03068_ _03054_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_77_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11560_ _05394_ _05399_ _05443_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_53_907 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_107_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10511_ _04737_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11491_ _01903_ _05377_ _05380_ _05285_ _05213_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _06525_ decoded_imm_j\[10\] _06733_ mem_rdata_q\[30\] _06553_ VGND VGND VPWR
+ VPWR _06765_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10442_ net1190 _03348_ _04695_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_625 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_21_804 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13161_ _06723_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__clkbuf_2
X_10373_ net622 _03348_ _04658_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_859 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12112_ _03098_ _05876_ _03083_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_150_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13092_ _06688_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12043_ mem_do_wdata _01860_ _05813_ _01862_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15802_ clknet_leaf_20_clk _01377_ VGND VGND VPWR VPWR cpuregs\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_13994_ net621 _06950_ _01613_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__mux2_1
X_15733_ clknet_leaf_144_clk _01308_ VGND VGND VPWR VPWR cpuregs\[22\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _06607_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15664_ clknet_leaf_2_clk _01239_ VGND VGND VPWR VPWR cpuregs\[29\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
*XANTENNA_140 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ _05041_ _06561_ _06568_ _06562_ net597 VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__a32o_1
*XANTENNA_151 _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_162 _03431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14615_ clknet_leaf_154_clk _00273_ VGND VGND VPWR VPWR cpuregs\[21\]\[13\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_173 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11827_ count_cycle\[32\] count_cycle\[31\] _05661_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__and3_1
*XANTENNA_184 _05273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15595_ clknet_leaf_2_clk _01170_ VGND VGND VPWR VPWR cpuregs\[31\]\[12\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_195 reg_pc\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_419 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_126_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11758_ net531 _05613_ _05616_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__a21oi_1
X_14546_ clknet_leaf_55_clk _00204_ VGND VGND VPWR VPWR cpuregs\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10709_ _03281_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__buf_4
XFILLER_0_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11689_ _05551_ _05555_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__and2_1
X_14477_ clknet_leaf_37_clk _00135_ VGND VGND VPWR VPWR cpuregs\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13428_ _06871_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13359_ cpuregs\[19\]\[17\] _04854_ _06827_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__mux2_1
X_16078_ net108 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_1
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_8 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07920_ _02410_ _02411_ _02417_ _02418_ _02415_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__a221o_1
X_15029_ clknet_leaf_132_clk _00687_ VGND VGND VPWR VPWR count_cycle\[12\] sky130_fd_sc_hd__dfxtp_1
X_07851_ net207 VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__clkbuf_4
Xinput2 net422 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
X_07782_ _02265_ _02399_ _02401_ _02250_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09521_ cpuregs\[4\]\[14\] cpuregs\[5\]\[14\] cpuregs\[6\]\[14\] cpuregs\[7\]\[14\]
+ _03457_ _03464_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_88_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09452_ _03454_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08403_ _02044_ _02959_ _02951_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09383_ cpuregs\[28\]\[10\] cpuregs\[29\]\[10\] cpuregs\[30\]\[10\] cpuregs\[31\]\[10\]
+ _03554_ _03459_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__mux4_1
XFILLER_0_87_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_734 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08334_ net252 net227 _02561_ _02595_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08265_ _02316_ net220 _02598_ _02641_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_806 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_940 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07216_ mem_wordsize\[1\] VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08196_ _02411_ _02790_ _02796_ _02585_ VGND VGND VPWR VPWR alu_out\[19\] sky130_fd_sc_hd__a22o_2
XFILLER_0_131_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07147_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09719_ _03574_ _04165_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__and3_1
X_10991_ net1370 _04842_ _05006_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_623 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12730_ cpuregs\[31\]\[30\] _05974_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12661_ cpuregs\[24\]\[27\] cpuregs\[25\]\[27\] cpuregs\[26\]\[27\] cpuregs\[27\]\[27\]
+ _05970_ _03108_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14400_ clknet_leaf_138_clk _00063_ VGND VGND VPWR VPWR cpuregs\[11\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11612_ _05264_ _05489_ _05490_ _01903_ _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12592_ _06142_ _06337_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__or2_1
X_15380_ clknet_leaf_89_clk _00970_ VGND VGND VPWR VPWR decoded_imm\[28\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14331_ _01792_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__clkbuf_1
X_11543_ _05418_ net527 _05343_ _05428_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _01756_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_152_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11474_ _05208_ _05210_ _05338_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13213_ decoded_imm\[18\] _06752_ _06735_ _06755_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__o22a_1
X_10425_ net1344 _03295_ _04684_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__mux2_1
X_14193_ _01709_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_150_488 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13144_ _06715_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__clkbuf_1
X_10356_ net1165 _03295_ _04647_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13075_ _06674_ _06675_ _05763_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__a21oi_1
X_10287_ _04618_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__clkbuf_1
X_12026_ instr_jalr VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13977_ net633 _06933_ _01602_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15716_ clknet_leaf_38_clk _01291_ VGND VGND VPWR VPWR cpuregs\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12928_ decoded_imm_j\[9\] _01091_ _03169_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15647_ clknet_leaf_46_clk _01222_ VGND VGND VPWR VPWR cpuregs\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _06546_ _06559_ _06561_ _06562_ net557 VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__a32o_1
XFILLER_0_145_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15578_ clknet_leaf_20_clk _01153_ VGND VGND VPWR VPWR cpuregs\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14529_ clknet_leaf_137_clk _00187_ VGND VGND VPWR VPWR cpuregs\[13\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_452 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_22_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08050_ _02660_ _02661_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_255 VGND VGND VPWR VPWR picorv32_255/HI eoi[1] sky130_fd_sc_hd__conb_1
Xpicorv32_266 VGND VGND VPWR VPWR picorv32_266/HI eoi[12] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_114_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_277 VGND VGND VPWR VPWR picorv32_277/HI eoi[23] sky130_fd_sc_hd__conb_1
Xpicorv32_288 VGND VGND VPWR VPWR picorv32_288/HI mem_la_addr[0] sky130_fd_sc_hd__conb_1
Xpicorv32_299 VGND VGND VPWR VPWR picorv32_299/HI pcpi_insn[9] sky130_fd_sc_hd__conb_1
X_08952_ _03426_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_102_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07903_ _02491_ _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__or2_1
X_08883_ reg_out\[28\] alu_out_q\[28\] _03176_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07834_ _02428_ _02429_ net187 _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__a211o_1
X_07765_ count_instr\[31\] _01949_ count_cycle\[63\] _01947_ VGND VGND VPWR VPWR _02386_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_100 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09504_ _03894_ _03902_ _03928_ _03964_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07696_ count_instr\[58\] _02052_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_79_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09435_ _03766_ _03897_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_111_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ _03767_ _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08317_ _02441_ _02899_ _02907_ _02608_ VGND VGND VPWR VPWR alu_out\[29\] sky130_fd_sc_hd__a22o_1
XFILLER_0_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_40 _03262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09297_ _02066_ _03396_ _03764_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_51 _03420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_62 _03525_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_73 _03674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08248_ _02801_ _02818_ _02831_ _02838_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__nor4_2
XTAP_TAPCELL_ROW_134_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_84 _04852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_95 _05925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08179_ _02414_ _02581_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10210_ net914 _03263_ _04575_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__mux2_1
X_11190_ _05040_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10141_ _04540_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_120_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput180 net180 VGND VGND VPWR VPWR pcpi_rs1[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput191 net253 VGND VGND VPWR VPWR pcpi_rs1[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10072_ _04502_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__clkbuf_1
X_13900_ _01565_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__buf_6
X_14880_ clknet_leaf_149_clk _00538_ VGND VGND VPWR VPWR cpuregs\[17\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_13831_ _07099_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13762_ _04483_ _03183_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__nor2_4
X_10974_ cpuregs\[17\]\[3\] _04825_ _04995_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__mux2_1
X_15501_ clknet_leaf_90_clk _01086_ VGND VGND VPWR VPWR mem_rdata_q\[24\] sky130_fd_sc_hd__dfxtp_1
X_12713_ _06447_ _06449_ _06451_ _06453_ _05978_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_48_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_520 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13693_ _07026_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15432_ clknet_leaf_126_clk _01022_ VGND VGND VPWR VPWR cpuregs\[18\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12644_ cpuregs\[16\]\[26\] cpuregs\[17\]\[26\] cpuregs\[18\]\[26\] cpuregs\[19\]\[26\]
+ _05921_ _05985_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15363_ clknet_leaf_69_clk _00953_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dfxtp_1
X_12575_ cpuregs\[28\]\[23\] cpuregs\[29\]\[23\] cpuregs\[30\]\[23\] cpuregs\[31\]\[23\]
+ _06191_ _05914_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_463 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14314_ _01783_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__clkbuf_1
X_11526_ _05217_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__inv_2
Xwire241 _06586_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15294_ clknet_leaf_76_clk _00003_ VGND VGND VPWR VPWR is_sltiu_bltu_sltu sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11457_ _05290_ _05293_ _05347_ _05315_ _05348_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__a2111o_1
X_14245_ net663 VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_111_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10408_ net937 _03241_ _04673_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__mux2_1
X_14176_ _01712_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__clkbuf_1
X_11388_ _01903_ _05282_ _05284_ _05285_ _05196_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__a32o_1
X_13127_ _06706_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__clkbuf_1
X_10339_ net1106 _03241_ _04636_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__mux2_1
X_13058_ net1123 _04877_ _06658_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__mux2_1
X_12009_ _05791_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07550_ _02175_ _02176_ _02186_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07481_ _02105_ _02111_ _02121_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09220_ cpuregs\[24\]\[5\] cpuregs\[25\]\[5\] cpuregs\[26\]\[5\] cpuregs\[27\]\[5\]
+ _03458_ _03461_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_372 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09151_ _01992_ _03622_ _03395_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__mux2_1
X_08102_ _02666_ _02684_ _02707_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__nand3_1
XFILLER_0_140_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09082_ cpuregs\[12\]\[2\] cpuregs\[13\]\[2\] cpuregs\[14\]\[2\] cpuregs\[15\]\[2\]
+ _03554_ _03408_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08033_ net200 _02645_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold800 cpuregs\[5\]\[28\] VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 cpuregs\[31\]\[12\] VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold822 cpuregs\[18\]\[13\] VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold833 cpuregs\[10\]\[27\] VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold844 cpuregs\[1\]\[27\] VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold855 cpuregs\[12\]\[25\] VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold866 cpuregs\[12\]\[11\] VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 cpuregs\[4\]\[22\] VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 cpuregs\[4\]\[31\] VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 count_cycle\[18\] VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ cpuregs\[0\]\[29\] cpuregs\[1\]\[29\] cpuregs\[2\]\[29\] cpuregs\[3\]\[29\]
+ _03800_ _03407_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08935_ _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__clkbuf_4
X_08866_ _03347_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__clkbuf_4
X_07817_ _02426_ _02427_ _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__a21oi_1
X_08797_ net678 _03287_ _03249_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__mux2_1
X_07748_ _01943_ _02369_ _02184_ _02370_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_114 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_95_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07679_ net17 _02202_ _02180_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_445 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09418_ _03448_ _03881_ _03468_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__o21a_1
X_10690_ _03240_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__buf_2
XFILLER_0_109_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09349_ cpuregs\[16\]\[9\] cpuregs\[17\]\[9\] cpuregs\[18\]\[9\] cpuregs\[19\]\[9\]
+ _03548_ _03549_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_320 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12360_ _03142_ _06111_ _06115_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11311_ _05194_ reg_pc\[16\] _01843_ _05226_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__o211a_1
X_12291_ _06043_ _06045_ _06047_ _06049_ _03080_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__a221o_2
XFILLER_0_121_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14030_ _01634_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__clkbuf_1
X_11242_ net475 _05175_ _05141_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11173_ _05128_ _05129_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_294 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10124_ _04531_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932_ clknet_leaf_121_clk _00590_ VGND VGND VPWR VPWR count_instr\[41\] sky130_fd_sc_hd__dfxtp_1
X_10055_ _04493_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__clkbuf_1
X_14863_ clknet_leaf_42_clk _00521_ VGND VGND VPWR VPWR cpuregs\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13814_ net715 _06975_ _07086_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14794_ clknet_leaf_54_clk _00452_ VGND VGND VPWR VPWR cpuregs\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13745_ _07054_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10957_ _04989_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_63_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13676_ net742 _06973_ _07014_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__mux2_1
X_10888_ net760 _04875_ _04945_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15415_ clknet_leaf_27_clk _01005_ VGND VGND VPWR VPWR cpuregs\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12627_ cpuregs\[0\]\[26\] cpuregs\[1\]\[26\] cpuregs\[2\]\[26\] cpuregs\[3\]\[26\]
+ _05819_ _03125_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15346_ clknet_leaf_68_clk _00936_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12558_ _06302_ _06304_ _06305_ _03149_ _05815_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_887 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_41_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11509_ _05373_ _05383_ _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__and3_1
X_15277_ clknet_leaf_93_clk _00870_ VGND VGND VPWR VPWR decoded_rd\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold107 count_instr\[63\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ cpuregs\[24\]\[19\] cpuregs\[25\]\[19\] cpuregs\[26\]\[19\] cpuregs\[27\]\[19\]
+ _06074_ _05932_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__mux4_1
Xhold118 net167 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _02346_ VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14228_ _01739_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14159_ cpuregs\[7\]\[26\] _06979_ _01696_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_294 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _03220_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__buf_2
X_08651_ mem_rdata_q\[22\] net15 _03018_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__mux2_1
X_07602_ _02217_ _02220_ _02218_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__a21bo_1
X_08582_ cpuregs\[12\]\[3\] cpuregs\[13\]\[3\] cpuregs\[14\]\[3\] cpuregs\[15\]\[3\]
+ _03092_ _03098_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_626 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07533_ _01944_ _02165_ _02167_ _01928_ _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07464_ _02104_ _02105_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09203_ _03404_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__buf_8
XFILLER_0_146_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07395_ _02023_ _02024_ _02027_ _02039_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__o31a_1
X_09134_ _03436_ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09065_ net182 decoded_imm\[1\] VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__nand2_1
X_08016_ net249 net250 VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold630 cpuregs\[23\]\[22\] VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold641 cpuregs\[7\]\[20\] VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 cpuregs\[4\]\[4\] VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 count_instr\[38\] VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 cpuregs\[12\]\[28\] VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 cpuregs\[19\]\[9\] VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 cpuregs\[13\]\[24\] VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ _03455_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_129_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08918_ _01854_ _03389_ _03392_ net34 VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__o211a_1
X_09898_ _03746_ _04346_ _03603_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08849_ _03331_ _03332_ _03293_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_142_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ net503 _05683_ _05647_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_142_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _04912_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__clkbuf_1
X_11791_ _05639_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_45_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _06926_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__clkbuf_1
X_10742_ _04872_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10673_ cpuregs\[26\]\[3\] _04825_ _04819_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__mux2_1
X_13461_ _06889_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_137_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15200_ clknet_leaf_71_clk alu_out\[13\] VGND VGND VPWR VPWR alu_out_q\[13\] sky130_fd_sc_hd__dfxtp_1
X_12412_ cpuregs\[20\]\[16\] cpuregs\[21\]\[16\] cpuregs\[22\]\[16\] cpuregs\[23\]\[16\]
+ _06065_ _05922_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13392_ net1279 _04817_ _06852_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__mux2_1
X_15131_ clknet_leaf_108_clk _00757_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfxtp_1
X_12343_ _03087_ _06099_ _03153_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_857 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15062_ clknet_leaf_132_clk _00720_ VGND VGND VPWR VPWR count_cycle\[45\] sky130_fd_sc_hd__dfxtp_1
X_12274_ _06033_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_767 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11225_ count_instr\[55\] count_instr\[54\] _05162_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__and3_1
X_14013_ cpuregs\[5\]\[21\] _06969_ _01624_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__mux2_1
X_11156_ _05116_ _05117_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_56_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10107_ _04520_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__clkbuf_1
X_11087_ _05069_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__clkbuf_1
X_15964_ clknet_leaf_138_clk _01536_ VGND VGND VPWR VPWR cpuregs\[10\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_14915_ clknet_leaf_118_clk _00573_ VGND VGND VPWR VPWR count_instr\[24\] sky130_fd_sc_hd__dfxtp_1
X_10038_ latched_rd\[1\] latched_rd\[0\] VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__or2_1
X_15895_ clknet_leaf_133_clk _01467_ VGND VGND VPWR VPWR cpuregs\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14846_ clknet_leaf_147_clk _00504_ VGND VGND VPWR VPWR cpuregs\[20\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14777_ clknet_leaf_157_clk _00435_ VGND VGND VPWR VPWR cpuregs\[16\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11989_ net39 net70 _05774_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13728_ _07045_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13659_ net1357 _06956_ _07003_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07180_ _01845_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15329_ clknet_leaf_77_clk _00919_ VGND VGND VPWR VPWR is_alu_reg_reg sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_76_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_890 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09821_ _04203_ _04271_ _03483_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09752_ _03616_ _04204_ _04205_ _01942_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__o211a_1
X_08703_ reg_pc\[4\] reg_pc\[3\] reg_pc\[2\] VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__and3_1
X_09683_ _02222_ _03617_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__nor2_1
X_08634_ cpuregs\[24\]\[4\] cpuregs\[25\]\[4\] cpuregs\[26\]\[4\] cpuregs\[27\]\[4\]
+ _03150_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_124_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _03038_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07516_ _01845_ _01848_ net22 _01933_ net5 VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__a32o_1
X_08496_ _03024_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__buf_1
XFILLER_0_92_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_119_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07447_ _02081_ _02090_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07378_ reg_pc\[5\] decoded_imm\[5\] VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09117_ cpuregs\[12\]\[3\] cpuregs\[13\]\[3\] cpuregs\[14\]\[3\] cpuregs\[15\]\[3\]
+ _03587_ _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_594 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09048_ _03519_ _03521_ _03431_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold460 cpuregs\[25\]\[1\] VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 cpuregs\[13\]\[5\] VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ cpuregs\[17\]\[20\] _04860_ _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__mux2_1
Xhold482 cpuregs\[10\]\[0\] VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 mem_rdata_q\[8\] VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _06615_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__clkbuf_1
X_14700_ clknet_leaf_24_clk _00358_ VGND VGND VPWR VPWR cpuregs\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11912_ _05721_ _01842_ _05722_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__and3b_1
X_15680_ clknet_leaf_52_clk _01255_ VGND VGND VPWR VPWR cpuregs\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12892_ mem_rdata_q\[31\] mem_rdata_q\[30\] VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__nand2_1
X_14631_ clknet_leaf_130_clk _00289_ VGND VGND VPWR VPWR cpuregs\[21\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_11843_ count_cycle\[37\] _05673_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_138_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_618 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14562_ clknet_leaf_130_clk _00220_ VGND VGND VPWR VPWR cpuregs\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11774_ count_cycle\[13\] count_cycle\[14\] count_cycle\[15\] _05620_ VGND VGND VPWR
+ VPWR _05628_ sky130_fd_sc_hd__and4_4
X_13513_ _06916_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _04818_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__buf_4
X_14493_ clknet_leaf_3_clk _00151_ VGND VGND VPWR VPWR cpuregs\[30\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_13444_ net1144 _04871_ _06874_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10656_ _04814_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10587_ net814 _03374_ _04768_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__mux2_1
X_13375_ _06843_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_152_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15114_ clknet_leaf_74_clk _00740_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12326_ _03134_ _06082_ _03050_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15045_ clknet_leaf_120_clk _00703_ VGND VGND VPWR VPWR count_cycle\[28\] sky130_fd_sc_hd__dfxtp_1
X_12257_ _05912_ _06016_ _03123_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11208_ count_instr\[49\] count_instr\[48\] VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__and2_1
X_12188_ cpuregs\[28\]\[7\] cpuregs\[29\]\[7\] cpuregs\[30\]\[7\] cpuregs\[31\]\[7\]
+ _05895_ _05929_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11139_ net882 _05103_ _05090_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__o21ai_1
X_15947_ clknet_leaf_30_clk _01519_ VGND VGND VPWR VPWR cpuregs\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15878_ clknet_leaf_44_clk _01450_ VGND VGND VPWR VPWR cpuregs\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14829_ clknet_leaf_36_clk _00487_ VGND VGND VPWR VPWR cpuregs\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08350_ net205 _02927_ _02931_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__a21o_2
XFILLER_0_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07301_ cpu_state\[4\] VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_22_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08281_ _02871_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_152_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_152_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_132_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07232_ cpu_state\[3\] is_beq_bne_blt_bge_bltu_bgeu _01859_ _01890_ _01891_ VGND
+ VGND VPWR VPWR _01892_ sky130_fd_sc_hd__a32o_1
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07163_ instr_srai instr_slli instr_srli instr_lhu VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09804_ _03414_ _04255_ _03426_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__o21a_1
Xfanout247 net210 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_4
X_07996_ _02008_ _02611_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__or2_1
X_09735_ cpuregs\[12\]\[21\] cpuregs\[13\]\[21\] cpuregs\[14\]\[21\] cpuregs\[15\]\[21\]
+ _03808_ _03801_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_805 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09666_ cpuregs\[8\]\[19\] cpuregs\[9\]\[19\] cpuregs\[10\]\[19\] cpuregs\[11\]\[19\]
+ _03456_ _03441_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__mux4_1
X_08617_ cpuregs\[8\]\[4\] cpuregs\[9\]\[4\] cpuregs\[10\]\[4\] cpuregs\[11\]\[4\]
+ _03133_ _03134_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__mux4_1
X_09597_ decoded_imm\[16\] _02200_ _04026_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08548_ _03037_ _03067_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_143_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_143_clk sky130_fd_sc_hd__clkbuf_2
X_08479_ _03012_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_1
XFILLER_0_53_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10510_ cpuregs\[14\]\[25\] _03348_ _04731_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11490_ _05379_ _05212_ _05210_ _05208_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_80_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10441_ _04700_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_816 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10372_ _04663_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__clkbuf_1
X_13160_ _01820_ _01894_ _06503_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__or3_2
XFILLER_0_20_315 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12111_ cpuregs\[22\]\[5\] cpuregs\[23\]\[5\] _03096_ VGND VGND VPWR VPWR _05876_
+ sky130_fd_sc_hd__mux2_1
X_13091_ net157 _02509_ _06685_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12042_ mem_do_wdata _05040_ _01955_ _05802_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__and4b_1
Xhold290 cpuregs\[27\]\[16\] VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15801_ clknet_leaf_141_clk _01376_ VGND VGND VPWR VPWR cpuregs\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_13993_ _01615_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_1
X_15732_ clknet_leaf_131_clk _01307_ VGND VGND VPWR VPWR cpuregs\[22\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12944_ _05495_ _01093_ _06587_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ clknet_leaf_5_clk _01238_ VGND VGND VPWR VPWR cpuregs\[29\]\[16\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_130 net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12875_ _05041_ _06560_ _06568_ _06562_ net551 VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__a32o_1
XFILLER_0_158_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_141 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_152 _01945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14614_ clknet_leaf_0_clk _00272_ VGND VGND VPWR VPWR cpuregs\[21\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11826_ net502 _05661_ _05663_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__a21oi_1
*XANTENNA_163 _03435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15594_ clknet_leaf_1_clk _01169_ VGND VGND VPWR VPWR cpuregs\[31\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_174 _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_185 _05358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_196 reg_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14545_ clknet_leaf_34_clk _00203_ VGND VGND VPWR VPWR cpuregs\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_134_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_134_clk sky130_fd_sc_hd__clkbuf_2
X_11757_ count_cycle\[10\] _05613_ _05141_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__o21ai_1
X_10708_ _04849_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14476_ clknet_leaf_27_clk _00134_ VGND VGND VPWR VPWR cpuregs\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11688_ _05251_ _05253_ _05540_ _05288_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_738 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_126_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13427_ cpuregs\[24\]\[17\] _04854_ _06863_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_157_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10639_ net1367 _03322_ _04804_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_654 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13358_ _06834_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12309_ _03143_ _06066_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16077_ net97 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
X_13289_ cpuregs\[18\]\[16\] _04852_ _06791_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__mux2_1
X_15028_ clknet_leaf_132_clk _00686_ VGND VGND VPWR VPWR count_cycle\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07850_ _02468_ _02469_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__and2_1
X_07781_ net215 _02400_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__nand2_1
Xinput3 net417 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
X_09520_ _03746_ _03980_ _03603_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_88_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_704 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09451_ cpuregs\[28\]\[12\] cpuregs\[29\]\[12\] cpuregs\[30\]\[12\] cpuregs\[31\]\[12\]
+ _03598_ _03460_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__mux4_1
X_08402_ reg_next_pc\[6\] reg_out\[6\] _02949_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__mux2_1
X_09382_ _03413_ _03846_ _03418_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_72 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_746 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08333_ _02910_ _02914_ _02919_ _02921_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_125_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_125_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08264_ _02584_ _02856_ _02857_ _02859_ _02430_ VGND VGND VPWR VPWR alu_out\[24\]
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_7_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_105_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07215_ net432 _01876_ _01879_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08195_ _02794_ _02795_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07146_ mem_do_rinst mem_do_prefetch VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07979_ _01978_ _02509_ _02594_ _02596_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__o22a_1
X_09718_ _04167_ _04169_ _04172_ _03575_ _03591_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__a221o_1
X_10990_ _05007_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09649_ _03746_ _04105_ _03603_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_167 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12660_ _03142_ _06398_ _06402_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_139_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _05032_ _05471_ _05237_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_116_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_116_clk sky130_fd_sc_hd__clkbuf_2
X_12591_ cpuregs\[20\]\[24\] cpuregs\[21\]\[24\] cpuregs\[22\]\[24\] cpuregs\[23\]\[24\]
+ _06065_ _03144_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__mux4_1
X_14330_ net912 _03262_ _01789_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__mux2_1
X_11542_ _05269_ _05425_ _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__a21o_1
X_14261_ net632 VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_401 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11473_ _05362_ _05363_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13212_ _06525_ decoded_imm_j\[18\] _06738_ net555 VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__a22o_1
X_10424_ _04691_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_840 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14192_ _01720_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13143_ net154 net116 _06707_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__mux2_1
X_10355_ _04654_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__clkbuf_1
X_10286_ net1012 _03287_ _04611_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__mux2_1
X_13074_ mem_do_rdata mem_do_rinst mem_state\[1\] mem_state\[0\] VGND VGND VPWR VPWR
+ _06675_ sky130_fd_sc_hd__or4b_1
X_12025_ _05799_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__clkbuf_1
X_13976_ _01606_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15715_ clknet_leaf_44_clk _01290_ VGND VGND VPWR VPWR cpuregs\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12927_ _06598_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15646_ clknet_leaf_23_clk _01221_ VGND VGND VPWR VPWR cpuregs\[23\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12858_ _06529_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__buf_2
XFILLER_0_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_618 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11809_ count_cycle\[25\] count_cycle\[26\] _05649_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__and3_1
X_15577_ clknet_leaf_141_clk _01152_ VGND VGND VPWR VPWR cpuregs\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_107_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_107_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_768 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12789_ _03021_ _01062_ _01063_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14528_ clknet_leaf_137_clk _00186_ VGND VGND VPWR VPWR cpuregs\[13\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_464 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14459_ clknet_leaf_10_clk _00117_ VGND VGND VPWR VPWR cpuregs\[12\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_126_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_147 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_256 VGND VGND VPWR VPWR picorv32_256/HI eoi[2] sky130_fd_sc_hd__conb_1
Xpicorv32_267 VGND VGND VPWR VPWR picorv32_267/HI eoi[13] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_114_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_278 VGND VGND VPWR VPWR picorv32_278/HI eoi[24] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_114_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_289 VGND VGND VPWR VPWR picorv32_289/HI mem_la_addr[1] sky130_fd_sc_hd__conb_1
X_08951_ _03425_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07902_ _02495_ _02520_ _02521_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__o21a_1
X_08882_ _03361_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07833_ net246 VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07764_ _02007_ net252 _02201_ _02384_ _01968_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_79_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09503_ decoded_imm\[13\] net175 VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07695_ _02071_ _02315_ _02318_ _02321_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__o31a_1
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09434_ _03765_ _03796_ _03896_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__or3b_1
XFILLER_0_149_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09365_ decoded_imm\[8\] net201 net202 decoded_imm\[9\] VGND VGND VPWR VPWR _03830_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_874 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_90_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08316_ _02905_ _02906_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09296_ _03397_ _03739_ _03763_ _03486_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__a211o_1
*XANTENNA_30 _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_41 _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_52 _03427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_844 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_63 _03547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08247_ _02585_ _02840_ _02843_ VGND VGND VPWR VPWR alu_out\[23\] sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_31_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_74 _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_85 _04854_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_760 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_96 _05927_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08178_ _02222_ net212 _02598_ _02641_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10140_ net1021 _03263_ _04537_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__mux2_1
Xoutput170 net170 VGND VGND VPWR VPWR mem_wstrb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput181 net181 VGND VGND VPWR VPWR pcpi_rs1[19] sky130_fd_sc_hd__clkbuf_4
Xoutput192 net192 VGND VGND VPWR VPWR pcpi_rs1[29] sky130_fd_sc_hd__buf_2
X_10071_ cpuregs\[12\]\[13\] _03268_ _04498_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13830_ _04524_ _04671_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__nor2_4
XFILLER_0_98_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13761_ _07062_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__clkbuf_1
X_10973_ _04998_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__clkbuf_1
X_15500_ clknet_leaf_91_clk _01085_ VGND VGND VPWR VPWR mem_rdata_q\[23\] sky130_fd_sc_hd__dfxtp_1
X_12712_ _03106_ _06452_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13692_ net932 _06989_ _06991_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15431_ clknet_leaf_148_clk _01021_ VGND VGND VPWR VPWR cpuregs\[18\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12643_ _03087_ _06386_ _03153_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_340 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15362_ clknet_leaf_68_clk _00952_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dfxtp_1
X_12574_ _06023_ _06320_ _05840_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313_ cpuregs\[10\]\[4\] _03208_ _01778_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__mux2_1
X_11525_ _05392_ _05401_ _05410_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15293_ clknet_leaf_76_clk _00002_ VGND VGND VPWR VPWR is_slti_blt_slt sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire242 net1417 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14244_ _01747_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11456_ _05323_ _05335_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10407_ _04682_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14175_ net1294 _06927_ _01710_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__mux2_1
X_11387_ _01891_ net361 VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__nand2_4
XFILLER_0_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13126_ net145 net107 _06696_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__mux2_1
X_10338_ _04645_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__clkbuf_1
X_13057_ _06666_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10269_ net1251 _03235_ _04600_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__mux2_1
X_12008_ net48 net79 _05785_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13959_ net1227 _06983_ _01588_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07480_ _02119_ _02120_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_510 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15629_ clknet_leaf_153_clk _01204_ VGND VGND VPWR VPWR cpuregs\[23\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09150_ _03476_ _03608_ _03615_ _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_384 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08101_ _02671_ _02683_ _02707_ _02708_ _02695_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__a32o_1
XFILLER_0_161_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09081_ _00012_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_116_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08032_ _02489_ _02644_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_25_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold801 cpuregs\[3\]\[31\] VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold812 cpuregs\[15\]\[7\] VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 cpuregs\[17\]\[18\] VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold834 cpuregs\[30\]\[16\] VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold845 cpuregs\[3\]\[27\] VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 cpuregs\[11\]\[12\] VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold867 cpuregs\[18\]\[12\] VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 cpuregs\[6\]\[11\] VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 cpuregs\[2\]\[23\] VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ cpuregs\[4\]\[29\] cpuregs\[5\]\[29\] cpuregs\[6\]\[29\] cpuregs\[7\]\[29\]
+ _03800_ _03407_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08934_ _03408_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__buf_8
XFILLER_0_110_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08865_ _03343_ _03346_ _03293_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__mux2_1
X_07816_ _02428_ _02429_ _02430_ _02431_ _02435_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__a221o_1
X_08796_ _03286_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07747_ net22 _02251_ _02179_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07678_ net187 VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_36_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09417_ cpuregs\[28\]\[11\] cpuregs\[29\]\[11\] cpuregs\[30\]\[11\] cpuregs\[31\]\[11\]
+ _03680_ _03443_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09348_ _03807_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09279_ cpuregs\[8\]\[7\] cpuregs\[9\]\[7\] cpuregs\[10\]\[7\] cpuregs\[11\]\[7\]
+ _03640_ _03492_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11310_ _01872_ _05225_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__or2_1
X_12290_ _03149_ _06048_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11241_ _05175_ _05176_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11172_ net1022 net374 _05090_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__o21ai_1
X_10123_ net1050 _03209_ _04526_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ clknet_leaf_114_clk _00589_ VGND VGND VPWR VPWR count_instr\[40\] sky130_fd_sc_hd__dfxtp_1
X_10054_ net1322 _03215_ _04487_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14862_ clknet_leaf_42_clk _00520_ VGND VGND VPWR VPWR cpuregs\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_730 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13813_ _07090_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__clkbuf_1
X_14793_ clknet_leaf_19_clk _00451_ VGND VGND VPWR VPWR cpuregs\[16\]\[31\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13744_ net1327 _06973_ _07050_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__mux2_1
X_10956_ net992 _04875_ _04981_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13675_ _07017_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__clkbuf_1
X_10887_ _04952_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__clkbuf_1
X_15414_ clknet_leaf_27_clk _01004_ VGND VGND VPWR VPWR cpuregs\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12626_ _05925_ _06369_ _03037_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__a21o_1
X_15345_ clknet_leaf_68_clk _00935_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfxtp_1
X_12557_ cpuregs\[16\]\[22\] cpuregs\[17\]\[22\] cpuregs\[18\]\[22\] cpuregs\[19\]\[22\]
+ _05921_ _05985_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11508_ decoded_imm_j\[9\] _05208_ _05359_ _05360_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15276_ clknet_leaf_93_clk _00869_ VGND VGND VPWR VPWR decoded_rd\[3\] sky130_fd_sc_hd__dfxtp_1
X_12488_ _06026_ _06238_ _06193_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__o21a_1
Xhold108 count_instr\[13\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold119 count_instr\[19\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ net638 _06979_ _01732_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11439_ decoded_imm_j\[8\] _05206_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_78_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14158_ _01702_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _06697_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__clkbuf_1
X_14089_ cpuregs\[6\]\[25\] _06977_ _01660_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08650_ _03163_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__clkbuf_1
X_07601_ _02232_ _02233_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__or2b_1
X_08581_ _03090_ _03099_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07532_ _02168_ _02169_ _01955_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07463_ reg_pc\[10\] decoded_imm\[10\] VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09202_ _03476_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07394_ _02023_ _02024_ _02027_ _02038_ _02039_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__o311a_1
XFILLER_0_72_630 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_8_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09133_ cpuregs\[24\]\[3\] cpuregs\[25\]\[3\] cpuregs\[26\]\[3\] cpuregs\[27\]\[3\]
+ _03594_ _03442_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09064_ _01846_ _03396_ _03524_ _03537_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__o22a_1
XFILLER_0_142_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_798 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08015_ _02608_ _02627_ _02629_ _02497_ VGND VGND VPWR VPWR alu_out\[5\] sky130_fd_sc_hd__a22o_1
Xhold620 cpuregs\[24\]\[26\] VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold631 cpuregs\[4\]\[20\] VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 cpuregs\[13\]\[3\] VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold653 cpuregs\[2\]\[16\] VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 cpuregs\[7\]\[23\] VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 cpuregs\[27\]\[20\] VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 cpuregs\[9\]\[1\] VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 cpuregs\[16\]\[0\] VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ cpuregs\[20\]\[28\] cpuregs\[21\]\[28\] cpuregs\[22\]\[28\] cpuregs\[23\]\[28\]
+ _03636_ _03637_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_129_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08917_ instr_sll _03391_ instr_slli cpu_state\[4\] VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_129_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ cpuregs\[24\]\[26\] cpuregs\[25\]\[26\] cpuregs\[26\]\[26\] cpuregs\[27\]\[26\]
+ _03640_ _03492_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_96_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08848_ reg_pc\[23\] _03326_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__xor2_1
X_08779_ reg_pc\[14\] reg_pc\[13\] _03259_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_142_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ cpuregs\[16\]\[22\] _04865_ _04909_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__mux2_1
X_11790_ _05637_ _05625_ _05638_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__and3b_1
XFILLER_0_79_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10741_ cpuregs\[26\]\[25\] _04871_ _04861_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13460_ net799 _04817_ _06888_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10672_ _03201_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12411_ _05879_ _06159_ _06161_ _06163_ _06164_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13391_ _06851_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_20_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_2
X_15130_ clknet_leaf_108_clk _00756_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfxtp_1
X_12342_ cpuregs\[22\]\[13\] cpuregs\[23\]\[13\] _05816_ VGND VGND VPWR VPWR _06099_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15061_ clknet_leaf_113_clk _00719_ VGND VGND VPWR VPWR count_cycle\[44\] sky130_fd_sc_hd__dfxtp_1
X_12273_ net248 _06032_ _05863_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_746 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14012_ _01625_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__clkbuf_1
X_11224_ net505 _05162_ _05164_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11155_ net471 _05112_ _05090_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_56_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10106_ net732 _03381_ _04486_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__mux2_1
X_11086_ _01884_ _05067_ _05068_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__and3_1
X_15963_ clknet_leaf_101_clk _01535_ VGND VGND VPWR VPWR cpuregs\[10\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_87_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_2
X_14914_ clknet_leaf_118_clk _00572_ VGND VGND VPWR VPWR count_instr\[23\] sky130_fd_sc_hd__dfxtp_1
X_10037_ latched_rd\[4\] latched_rd\[2\] latched_rd\[3\] VGND VGND VPWR VPWR _04481_
+ sky130_fd_sc_hd__nand3b_4
X_15894_ clknet_leaf_140_clk _01466_ VGND VGND VPWR VPWR cpuregs\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14845_ clknet_leaf_155_clk _00503_ VGND VGND VPWR VPWR cpuregs\[20\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_98_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14776_ clknet_leaf_151_clk _00434_ VGND VGND VPWR VPWR cpuregs\[16\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11988_ _05780_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13727_ cpuregs\[29\]\[15\] _06956_ _07039_ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__mux2_1
X_10939_ net710 _04858_ _04970_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13658_ _07008_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_82_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12609_ _06138_ _06353_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13589_ _03313_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__buf_2
XFILLER_0_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_836 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15328_ clknet_leaf_77_clk _00918_ VGND VGND VPWR VPWR is_alu_reg_imm sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15259_ clknet_leaf_77_clk _00852_ VGND VGND VPWR VPWR instr_fence sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09820_ net253 _03660_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__nor2_1
X_09751_ _02316_ _03480_ _04092_ _03074_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_78_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_2
X_08702_ reg_pc\[3\] _01971_ reg_pc\[4\] VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09682_ _02290_ _03480_ _04028_ _03074_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08633_ _03052_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _03082_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07515_ net175 VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08495_ mem_rdata_q\[16\] net8 _03018_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07446_ _01943_ _02082_ _02086_ _01927_ _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07377_ reg_pc\[5\] decoded_imm\[5\] VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09116_ _03441_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__buf_8
XFILLER_0_17_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_540 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_346 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09047_ _03403_ _03520_ _03427_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_368 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold450 cpuregs\[29\]\[13\] VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 cpuregs\[20\]\[22\] VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 cpuregs\[17\]\[5\] VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 cpuregs\[18\]\[1\] VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 cpuregs\[3\]\[16\] VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09949_ _04304_ _04305_ _04395_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_5_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_2
X_12960_ net439 _01072_ _06587_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11911_ count_cycle\[57\] _05716_ count_cycle\[58\] VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__a21o_1
X_12891_ mem_rdata_q\[29\] mem_rdata_q\[28\] mem_rdata_q\[19\] mem_rdata_q\[18\] VGND
+ VGND VPWR VPWR _06577_ sky130_fd_sc_hd__or4_1
X_14630_ clknet_leaf_127_clk _00288_ VGND VGND VPWR VPWR cpuregs\[21\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11842_ _05673_ _05674_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14561_ clknet_leaf_145_clk _00219_ VGND VGND VPWR VPWR cpuregs\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_11773_ _05627_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__clkbuf_1
X_13512_ net1349 _04871_ _06910_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _03313_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__clkbuf_4
X_14492_ clknet_leaf_154_clk _00150_ VGND VGND VPWR VPWR cpuregs\[30\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_687 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13443_ _06879_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__clkbuf_1
X_10655_ net847 _03374_ _04804_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_408 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13374_ net823 _04869_ _06838_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10586_ _04777_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15113_ clknet_leaf_105_clk _07138_ VGND VGND VPWR VPWR reg_out\[31\] sky130_fd_sc_hd__dfxtp_1
X_12325_ cpuregs\[6\]\[13\] cpuregs\[7\]\[13\] _03084_ VGND VGND VPWR VPWR _06082_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15044_ clknet_leaf_120_clk _00702_ VGND VGND VPWR VPWR count_cycle\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12256_ cpuregs\[12\]\[10\] cpuregs\[13\]\[10\] cpuregs\[14\]\[10\] cpuregs\[15\]\[10\]
+ _05913_ _05994_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__mux4_1
X_11207_ net458 VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_79_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12187_ _03090_ _05949_ _05927_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_71_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ count_instr\[28\] _05103_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__and2_1
X_11069_ _05055_ _05056_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__nor2_1
X_15946_ clknet_leaf_58_clk _01518_ VGND VGND VPWR VPWR cpuregs\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_0_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_116_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15877_ clknet_leaf_37_clk _01449_ VGND VGND VPWR VPWR cpuregs\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14828_ clknet_leaf_23_clk _00486_ VGND VGND VPWR VPWR cpuregs\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14759_ clknet_leaf_127_clk _00417_ VGND VGND VPWR VPWR cpuregs\[26\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_928 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07300_ count_instr\[0\] _01949_ _01951_ count_cycle\[0\] VGND VGND VPWR VPWR _01952_
+ sky130_fd_sc_hd__a22o_1
X_08280_ _02849_ _02855_ _02864_ _02873_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__o31a_1
XFILLER_0_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07231_ cpu_state\[1\] VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_173 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07162_ instr_sll instr_sub instr_add instr_andi VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09803_ cpuregs\[16\]\[23\] cpuregs\[17\]\[23\] cpuregs\[18\]\[23\] cpuregs\[19\]\[23\]
+ _03673_ _03674_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_161_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout248 net204 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_2
X_07995_ net250 _02610_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__xor2_1
X_09734_ _03557_ _04187_ _03417_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__o21a_1
X_09665_ _04119_ _04120_ _03552_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_828 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08616_ _03063_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__clkbuf_8
X_09596_ _04052_ _04053_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_159_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08547_ cpuregs\[12\]\[2\] cpuregs\[13\]\[2\] cpuregs\[14\]\[2\] cpuregs\[15\]\[2\]
+ _00007_ _00008_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08478_ _02369_ _03011_ _02993_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_544 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_624 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07429_ reg_pc\[8\] decoded_imm\[8\] VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10440_ net934 _03341_ _04695_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10371_ net1086 _03341_ _04658_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12110_ _05873_ _05874_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13090_ _06687_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12041_ net733 _01860_ _01866_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__a21o_1
Xhold280 cpuregs\[18\]\[8\] VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold291 cpuregs\[8\]\[16\] VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15800_ clknet_leaf_132_clk _01375_ VGND VGND VPWR VPWR cpuregs\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_13992_ net768 _06948_ _01613_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__mux2_1
X_15731_ clknet_leaf_146_clk _01306_ VGND VGND VPWR VPWR cpuregs\[22\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12943_ _06606_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__buf_1
XFILLER_0_99_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15662_ clknet_leaf_3_clk _01237_ VGND VGND VPWR VPWR cpuregs\[29\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
*XANTENNA_120 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12874_ _05041_ _06538_ _06568_ _06562_ net635 VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__a32o_1
*XANTENNA_131 net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_142 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14613_ clknet_leaf_0_clk _00271_ VGND VGND VPWR VPWR cpuregs\[21\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11825_ net502 net363 _05622_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__o21ai_1
*XANTENNA_153 _02082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15593_ clknet_leaf_1_clk _01168_ VGND VGND VPWR VPWR cpuregs\[31\]\[10\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_164 _03435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_175 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_186 _05758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
*XANTENNA_197 reg_pc\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14544_ clknet_leaf_32_clk _00202_ VGND VGND VPWR VPWR cpuregs\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11756_ _05615_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_56_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10707_ net863 _04848_ _04840_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__mux2_1
X_14475_ clknet_leaf_53_clk _00133_ VGND VGND VPWR VPWR cpuregs\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11687_ _05253_ _05548_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13426_ _06870_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10638_ _04805_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13357_ cpuregs\[19\]\[16\] _04852_ _06827_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_830 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10569_ net1034 _03314_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12308_ cpuregs\[20\]\[12\] cpuregs\[21\]\[12\] cpuregs\[22\]\[12\] cpuregs\[23\]\[12\]
+ _06065_ _05922_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__mux4_1
X_13288_ _06797_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__clkbuf_1
X_15027_ clknet_leaf_113_clk net532 VGND VGND VPWR VPWR count_cycle\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12239_ cpuregs\[20\]\[9\] cpuregs\[21\]\[9\] cpuregs\[22\]\[9\] cpuregs\[23\]\[9\]
+ _05921_ _05922_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__mux4_1
X_07780_ _02265_ net216 VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__xnor2_1
Xinput4 net482 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
X_15929_ clknet_leaf_129_clk _01501_ VGND VGND VPWR VPWR cpuregs\[0\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09450_ _03414_ _03912_ _03419_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_121_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08401_ _02958_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_1
X_09381_ cpuregs\[24\]\[10\] cpuregs\[25\]\[10\] cpuregs\[26\]\[10\] cpuregs\[27\]\[10\]
+ _03404_ _03408_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08332_ net240 VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08263_ _02431_ _02569_ _02858_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07214_ instr_sw _01874_ _01866_ instr_lw _01878_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08194_ _02785_ _02787_ _02784_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07978_ _01978_ _02509_ _02561_ _02595_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__a31o_1
X_09717_ _04170_ _04171_ _03447_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__mux2_1
X_09648_ cpuregs\[8\]\[18\] cpuregs\[9\]\[18\] cpuregs\[10\]\[18\] cpuregs\[11\]\[18\]
+ _03640_ _03492_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__mux4_1
X_09579_ cpuregs\[28\]\[16\] cpuregs\[29\]\[16\] cpuregs\[30\]\[16\] cpuregs\[31\]\[16\]
+ _03440_ _03451_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_179 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _05233_ _05235_ _05237_ _05457_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_139_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _06177_ _06331_ _06333_ _06335_ _06164_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11541_ _05273_ _05222_ _05426_ _01903_ _05184_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14260_ _01755_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__clkbuf_1
X_11472_ decoded_imm_j\[9\] _05208_ _05353_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_152_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13211_ decoded_imm\[19\] _06752_ _06735_ _06754_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10423_ net1180 _03287_ _04684_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__mux2_1
X_14191_ net935 _06943_ _01710_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_474 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_104_852 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13142_ _06714_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__clkbuf_1
X_10354_ cpuregs\[28\]\[16\] _03287_ _04647_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13073_ mem_do_wdata _01856_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__or2_1
X_10285_ _04617_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__clkbuf_1
X_12024_ net57 net88 _05766_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13975_ net553 _06931_ _01602_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__mux2_1
X_15714_ clknet_leaf_39_clk _01289_ VGND VGND VPWR VPWR cpuregs\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12926_ mem_rdata_q\[29\] net22 _06589_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15645_ clknet_leaf_23_clk _01220_ VGND VGND VPWR VPWR cpuregs\[23\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12857_ _06532_ mem_rdata_q\[13\] _06533_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__and3b_1
XFILLER_0_158_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11808_ net504 _05649_ _05651_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15576_ clknet_leaf_133_clk _01151_ VGND VGND VPWR VPWR cpuregs\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12788_ _06517_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_83_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_190 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_139_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11739_ net508 _05601_ _05603_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14527_ clknet_leaf_97_clk _00185_ VGND VGND VPWR VPWR cpuregs\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14458_ clknet_leaf_11_clk _00116_ VGND VGND VPWR VPWR cpuregs\[12\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13409_ _06861_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14389_ clknet_leaf_12_clk _00052_ VGND VGND VPWR VPWR cpuregs\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_800 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_257 VGND VGND VPWR VPWR picorv32_257/HI eoi[3] sky130_fd_sc_hd__conb_1
XFILLER_0_12_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_268 VGND VGND VPWR VPWR picorv32_268/HI eoi[14] sky130_fd_sc_hd__conb_1
X_08950_ _00015_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_114_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_279 VGND VGND VPWR VPWR picorv32_279/HI eoi[25] sky130_fd_sc_hd__conb_1
X_07901_ _02044_ _02492_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__or2b_1
X_08881_ net1071 _03360_ _03315_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07832_ net188 net220 VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_16_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07763_ net25 _02252_ _02180_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__a21o_1
X_09502_ _03961_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_154_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07694_ _02017_ _02320_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_78_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09433_ _03834_ _03863_ _03864_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ _03829_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08315_ _02458_ _02891_ _02894_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_268 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_20 _03108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09295_ _01943_ _03740_ _03742_ _03488_ _03762_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__a32o_1
*XANTENNA_31 _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
*XANTENNA_42 _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_53 _03438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08246_ _02290_ net218 _02841_ _02842_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_31_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_64 _03549_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
*XANTENNA_75 _03746_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
*XANTENNA_86 _04854_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_97 _05932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_772 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08177_ _02608_ _02775_ _02776_ _02779_ VGND VGND VPWR VPWR alu_out\[17\] sky130_fd_sc_hd__a31o_1
XFILLER_0_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput160 net160 VGND VGND VPWR VPWR mem_wdata[3] sky130_fd_sc_hd__buf_2
Xoutput171 net171 VGND VGND VPWR VPWR pcpi_rs1[0] sky130_fd_sc_hd__clkbuf_4
Xoutput182 net182 VGND VGND VPWR VPWR pcpi_rs1[1] sky130_fd_sc_hd__clkbuf_4
X_10070_ _04501_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_1
Xoutput193 net193 VGND VGND VPWR VPWR pcpi_rs1[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13760_ net1351 _06989_ _07027_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10972_ net634 _04823_ _04995_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__mux2_1
X_12711_ cpuregs\[24\]\[29\] cpuregs\[25\]\[29\] cpuregs\[26\]\[29\] cpuregs\[27\]\[29\]
+ _03150_ _03151_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13691_ _07025_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_680 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12642_ cpuregs\[22\]\[26\] cpuregs\[23\]\[26\] _05979_ VGND VGND VPWR VPWR _06386_
+ sky130_fd_sc_hd__mux2_1
X_15430_ clknet_leaf_149_clk _01020_ VGND VGND VPWR VPWR cpuregs\[18\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_155_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15361_ clknet_leaf_69_clk _00951_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12573_ cpuregs\[16\]\[23\] cpuregs\[17\]\[23\] cpuregs\[18\]\[23\] cpuregs\[19\]\[23\]
+ _05984_ _06068_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_739 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_124_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11524_ _05392_ _05401_ _05410_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__and3_1
X_14312_ _01782_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_61_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15292_ clknet_leaf_78_clk _00884_ VGND VGND VPWR VPWR is_sll_srl_sra sky130_fd_sc_hd__dfxtp_1
Xwire243 _03659_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_4
X_14243_ net702 VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11455_ _05304_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10406_ net1371 _03235_ _04673_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14174_ _01711_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11386_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13125_ _06705_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10337_ cpuregs\[28\]\[8\] _03235_ _04636_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__mux2_1
X_13056_ net1203 _04875_ _06658_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__mux2_1
X_10268_ _04608_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__clkbuf_1
X_12007_ _05790_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10199_ cpuregs\[13\]\[7\] _03228_ _04564_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13958_ _01596_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12909_ _03017_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__buf_4
X_13889_ _01559_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_17_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15628_ clknet_leaf_154_clk _01203_ VGND VGND VPWR VPWR cpuregs\[23\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15559_ clknet_leaf_57_clk _01134_ VGND VGND VPWR VPWR cpuregs\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_08100_ _02680_ _02694_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09080_ _03550_ _03551_ _03552_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08031_ _02492_ _02609_ _02630_ _02573_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__o31a_1
XFILLER_0_141_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_744 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold802 cpuregs\[31\]\[13\] VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold813 count_instr\[21\] VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold824 cpuregs\[11\]\[3\] VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold835 cpuregs\[10\]\[7\] VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 cpuregs\[3\]\[17\] VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 cpuregs\[13\]\[27\] VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold868 cpuregs\[4\]\[28\] VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _04424_ _04425_ _04426_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__o21ai_1
Xhold879 cpuregs\[23\]\[17\] VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ _03407_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08864_ _03344_ _03345_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__nor2_1
X_07815_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__inv_2
X_08795_ _03284_ _03285_ _03261_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__mux2_4
X_07746_ net192 VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07677_ _02300_ _02303_ _01945_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_36_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09416_ _03437_ _03879_ _03426_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09347_ cpuregs\[20\]\[9\] cpuregs\[21\]\[9\] cpuregs\[22\]\[9\] cpuregs\[23\]\[9\]
+ _03438_ _03812_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09278_ _03413_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08229_ _02399_ _02813_ instr_sub VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_783 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11240_ net498 _05172_ _05169_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11171_ count_instr\[38\] _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10122_ _04530_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_42_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14930_ clknet_leaf_114_clk _00588_ VGND VGND VPWR VPWR count_instr\[39\] sky130_fd_sc_hd__dfxtp_1
X_10053_ _04492_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__clkbuf_1
X_14861_ clknet_leaf_37_clk _00519_ VGND VGND VPWR VPWR cpuregs\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_13812_ net1153 _06973_ _07086_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_742 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14792_ clknet_leaf_23_clk _00450_ VGND VGND VPWR VPWR cpuregs\[16\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13743_ _07053_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__clkbuf_1
X_10955_ _04988_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13674_ net989 _06971_ _07014_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__mux2_1
X_10886_ net873 _04873_ _04945_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15413_ clknet_leaf_42_clk _01003_ VGND VGND VPWR VPWR cpuregs\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12625_ cpuregs\[6\]\[26\] cpuregs\[7\]\[26\] _03084_ VGND VGND VPWR VPWR _06369_
+ sky130_fd_sc_hd__mux2_1
X_15344_ clknet_leaf_68_clk _00934_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfxtp_2
X_12556_ _03087_ _06303_ _03153_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_136_571 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11507_ reg_next_pc\[12\] _02999_ _05214_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12487_ cpuregs\[28\]\[19\] cpuregs\[29\]\[19\] cpuregs\[30\]\[19\] cpuregs\[31\]\[19\]
+ _06191_ _05929_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__mux4_1
X_15275_ clknet_leaf_92_clk _00868_ VGND VGND VPWR VPWR decoded_rd\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold109 _00562_ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
X_14226_ _01738_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__clkbuf_1
X_11438_ _05324_ _05323_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_78_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14157_ cpuregs\[7\]\[25\] _06977_ _01696_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11369_ _01890_ _05191_ _05193_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ net136 net98 _06696_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__mux2_1
X_14088_ _01665_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13039_ cpuregs\[1\]\[19\] _04858_ _06647_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07600_ reg_pc\[19\] decoded_imm\[19\] VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_21 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08580_ cpuregs\[8\]\[3\] cpuregs\[9\]\[3\] cpuregs\[10\]\[3\] cpuregs\[11\]\[3\]
+ _03096_ _03098_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__mux4_1
X_07531_ count_instr\[14\] _01949_ count_cycle\[14\] _01951_ VGND VGND VPWR VPWR _02169_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07462_ reg_pc\[10\] decoded_imm\[10\] VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09201_ _02044_ _03481_ _03669_ _03670_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07393_ _02025_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09132_ _03402_ _03602_ _03603_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09063_ reg_pc\[1\] _03488_ _03528_ _03536_ _03486_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__a311o_1
XFILLER_0_25_580 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08014_ _02496_ _02581_ _02628_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__a21o_1
Xhold610 cpuregs\[20\]\[8\] VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 cpuregs\[17\]\[16\] VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_130_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold632 cpuregs\[29\]\[6\] VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 cpuregs\[22\]\[4\] VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 cpuregs\[26\]\[20\] VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 cpuregs\[23\]\[11\] VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold676 cpuregs\[30\]\[25\] VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 cpuregs\[21\]\[29\] VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 cpuregs\[11\]\[31\] VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _03434_ _04407_ _04409_ _04411_ _03490_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08916_ instr_srl instr_srli _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_129_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _04343_ _04344_ _03579_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__mux2_1
X_08847_ reg_out\[23\] alu_out_q\[23\] _03175_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_108_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08778_ reg_pc\[13\] _03259_ reg_pc\[14\] VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_142_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _02304_ _02312_ _02350_ _02352_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_0_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _03347_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_756 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_95_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10671_ _04824_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_137_357 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_806 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12410_ _00011_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__buf_4
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ _04485_ _04744_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__nor2_4
XFILLER_0_62_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12341_ _05872_ _06097_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15060_ clknet_leaf_132_clk _00718_ VGND VGND VPWR VPWR count_cycle\[43\] sky130_fd_sc_hd__dfxtp_1
X_12272_ _05901_ _06020_ _06031_ _05904_ decoded_imm\[10\] VGND VGND VPWR VPWR _06032_
+ sky130_fd_sc_hd__a32o_2
X_14011_ net1051 _06966_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11223_ count_instr\[54\] _05162_ _05141_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11154_ count_instr\[33\] count_instr\[32\] count_instr\[31\] _05109_ VGND VGND VPWR
+ VPWR _05116_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ _04519_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11085_ count_instr\[12\] _05065_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__nand2_1
X_15962_ clknet_leaf_135_clk _01534_ VGND VGND VPWR VPWR cpuregs\[10\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_14913_ clknet_leaf_119_clk _00571_ VGND VGND VPWR VPWR count_instr\[22\] sky130_fd_sc_hd__dfxtp_1
X_10036_ _03396_ _04461_ _04479_ _04480_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__a31o_1
X_15893_ clknet_leaf_15_clk _01465_ VGND VGND VPWR VPWR cpuregs\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14844_ clknet_leaf_152_clk _00502_ VGND VGND VPWR VPWR cpuregs\[20\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14775_ clknet_leaf_151_clk _00433_ VGND VGND VPWR VPWR cpuregs\[16\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11987_ net38 net69 _05774_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13726_ _07044_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__clkbuf_1
X_10938_ _04979_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_650 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13657_ cpuregs\[23\]\[14\] _06954_ _07003_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__mux2_1
X_10869_ net875 _04856_ _04934_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12608_ cpuregs\[8\]\[25\] cpuregs\[9\]\[25\] cpuregs\[10\]\[25\] cpuregs\[11\]\[25\]
+ _06061_ _03137_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__mux4_1
X_13588_ _06965_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15327_ clknet_leaf_20_clk _00917_ VGND VGND VPWR VPWR cpuregs\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_390 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12539_ _05925_ _06286_ _03050_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15258_ clknet_leaf_112_clk _00851_ VGND VGND VPWR VPWR instr_rdinstr sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14209_ _01729_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__clkbuf_1
X_15189_ clknet_leaf_70_clk alu_out\[2\] VGND VGND VPWR VPWR alu_out_q\[2\] sky130_fd_sc_hd__dfxtp_1
X_09750_ _02277_ _03770_ _04203_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__o21ba_1
X_08701_ reg_out\[4\] alu_out_q\[4\] latched_stalu VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__mux2_1
X_09681_ _03476_ _04136_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08632_ _03046_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__buf_8
XFILLER_0_146_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08563_ _03037_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07514_ _02151_ _02152_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08494_ _03023_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07445_ _02087_ _02088_ _01954_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__o21a_2
XFILLER_0_91_203 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_92_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07376_ _02003_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09115_ _03586_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__buf_8
XFILLER_0_143_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09046_ cpuregs\[8\]\[1\] cpuregs\[9\]\[1\] cpuregs\[10\]\[1\] cpuregs\[11\]\[1\]
+ _03494_ _03497_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_678 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold440 cpuregs\[9\]\[0\] VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 cpuregs\[3\]\[4\] VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 cpuregs\[14\]\[29\] VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 cpuregs\[22\]\[25\] VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 cpuregs\[9\]\[8\] VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 net52 VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__dlygate4sd3_1
X_09948_ _04337_ _04384_ _04385_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_5_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _02306_ _03617_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__nor2_1
X_11910_ _05706_ _05713_ _05720_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__and3_1
X_12890_ net443 net564 _06575_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__nor3_1
XFILLER_0_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11841_ net520 _05670_ _05647_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__o21ai_1
X_11772_ _05624_ _05625_ _05626_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__and3b_1
X_14560_ clknet_leaf_142_clk _00218_ VGND VGND VPWR VPWR cpuregs\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10723_ _04859_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__clkbuf_1
X_13511_ _06915_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14491_ clknet_leaf_2_clk _00149_ VGND VGND VPWR VPWR cpuregs\[30\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13442_ net1003 _04869_ _06874_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10654_ _04813_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_82_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13373_ _06842_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10585_ net749 _03367_ _04768_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__mux2_1
X_15112_ clknet_leaf_105_clk _07137_ VGND VGND VPWR VPWR reg_out\[30\] sky130_fd_sc_hd__dfxtp_1
X_12324_ _05871_ _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15043_ clknet_leaf_120_clk _00701_ VGND VGND VPWR VPWR count_cycle\[26\] sky130_fd_sc_hd__dfxtp_1
X_12255_ _06012_ _06013_ _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11206_ _05152_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__clkbuf_1
X_12186_ cpuregs\[16\]\[7\] cpuregs\[17\]\[7\] cpuregs\[18\]\[7\] cpuregs\[19\]\[7\]
+ _05948_ _05925_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11137_ _05103_ _05104_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11068_ net765 _05053_ _05044_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__o21ai_1
X_15945_ clknet_leaf_36_clk _01517_ VGND VGND VPWR VPWR cpuregs\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_10019_ _04462_ _04463_ _03414_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__mux2_1
X_15876_ clknet_leaf_26_clk _01448_ VGND VGND VPWR VPWR cpuregs\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14827_ clknet_leaf_52_clk _00485_ VGND VGND VPWR VPWR cpuregs\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_59_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14758_ clknet_leaf_148_clk _00416_ VGND VGND VPWR VPWR cpuregs\[26\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_406 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13709_ _07035_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_597 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14689_ clknet_leaf_147_clk _00347_ VGND VGND VPWR VPWR cpuregs\[27\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07230_ _01889_ decoder_trigger VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__nand2_4
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_88 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_143_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07161_ _00001_ _01825_ _01826_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_70_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09802_ _03647_ _04253_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout249 net124 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_4
X_07994_ _02573_ _02609_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__nand2_1
X_09733_ cpuregs\[8\]\[21\] cpuregs\[9\]\[21\] cpuregs\[10\]\[21\] cpuregs\[11\]\[21\]
+ _03586_ _03449_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__mux4_1
X_09664_ cpuregs\[0\]\[19\] cpuregs\[1\]\[19\] cpuregs\[2\]\[19\] cpuregs\[3\]\[19\]
+ _03808_ _03801_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__mux4_1
X_08615_ _03051_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__clkbuf_8
X_09595_ decoded_imm\[17\] _02213_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_159_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ cpuregs\[8\]\[2\] cpuregs\[9\]\[2\] cpuregs\[10\]\[2\] cpuregs\[11\]\[2\]
+ _03046_ _03052_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__mux4_1
X_08477_ reg_next_pc\[29\] reg_out\[29\] _02991_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07428_ _02019_ _02057_ _02072_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_21_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07359_ _01958_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_111 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_61_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10370_ _04662_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_894 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_143_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09029_ cpuregs\[24\]\[1\] cpuregs\[25\]\[1\] cpuregs\[26\]\[1\] cpuregs\[27\]\[1\]
+ _03406_ _03410_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12040_ _02558_ _03672_ _05802_ _05804_ _05812_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__a41o_1
Xhold270 cpuregs\[21\]\[19\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_385 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold281 cpuregs\[31\]\[14\] VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 reg_next_pc\[9\] VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13991_ _01614_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15730_ clknet_leaf_155_clk _01305_ VGND VGND VPWR VPWR cpuregs\[22\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12942_ mem_rdata_q\[31\] net430 _06589_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ clknet_leaf_143_clk _01236_ VGND VGND VPWR VPWR cpuregs\[29\]\[14\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_110 decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12873_ _06567_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__clkbuf_2
*XANTENNA_121 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_132 net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14612_ clknet_leaf_2_clk _00270_ VGND VGND VPWR VPWR cpuregs\[21\]\[10\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_143 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11824_ net362 _05662_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__nor2_1
X_15592_ clknet_leaf_33_clk _01167_ VGND VGND VPWR VPWR cpuregs\[31\]\[9\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_154 _02251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_165 _03443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_176 _04672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_187 _05871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
*XANTENNA_198 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14543_ clknet_leaf_41_clk _00201_ VGND VGND VPWR VPWR cpuregs\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11755_ _05613_ _05113_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_101_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10706_ _03274_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_707 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14474_ clknet_leaf_45_clk _00132_ VGND VGND VPWR VPWR cpuregs\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11686_ _05418_ net483 _05358_ _05559_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13425_ net658 _04852_ _06863_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__mux2_1
X_10637_ net1310 _03314_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_106_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_179 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10568_ _04745_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13356_ _06833_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12307_ _03046_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__clkbuf_8
X_13287_ net1290 _04850_ _06791_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__mux2_1
X_10499_ _04708_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15026_ clknet_leaf_113_clk _00684_ VGND VGND VPWR VPWR count_cycle\[9\] sky130_fd_sc_hd__dfxtp_1
X_12238_ _05879_ _05993_ _05996_ _05998_ _03104_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__a221o_2
X_12169_ cpuregs\[24\]\[6\] cpuregs\[25\]\[6\] cpuregs\[26\]\[6\] cpuregs\[27\]\[6\]
+ _03095_ _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__mux4_1
Xinput5 net492 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_15928_ clknet_leaf_141_clk _01500_ VGND VGND VPWR VPWR cpuregs\[0\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_88_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15859_ clknet_leaf_7_clk _01431_ VGND VGND VPWR VPWR cpuregs\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08400_ _02030_ _02957_ _02951_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__mux2_1
X_09380_ _03843_ _03844_ _03807_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__mux2_1
X_08331_ _02910_ _02914_ _02919_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08262_ _02306_ net246 _02618_ _02562_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07213_ _01877_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08193_ net181 _02793_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07977_ _02562_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__clkbuf_4
X_09716_ cpuregs\[0\]\[20\] cpuregs\[1\]\[20\] cpuregs\[2\]\[20\] cpuregs\[3\]\[20\]
+ _03457_ _03595_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09647_ _03454_ _04103_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09578_ _03500_ _04036_ _03468_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _03045_ _03048_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_139_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11540_ _05222_ _05414_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11471_ _05359_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10422_ _04690_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__clkbuf_1
X_13210_ _06525_ decoded_imm_j\[19\] _06738_ net541 VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__a22o_1
X_14190_ _01719_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10353_ _04653_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13141_ net153 net115 _06707_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13072_ mem_do_wdata _06672_ _06673_ net514 VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__a2bb2o_1
X_10284_ net584 _03282_ _04611_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__mux2_1
X_12023_ _05798_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13974_ _01605_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__clkbuf_1
X_15713_ clknet_leaf_28_clk _01288_ VGND VGND VPWR VPWR cpuregs\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12925_ _06597_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_103_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15644_ clknet_leaf_130_clk _01219_ VGND VGND VPWR VPWR cpuregs\[23\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12856_ _06546_ _06560_ _06559_ _06530_ net491 VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11807_ net1408 _05649_ _05622_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_83_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ clknet_leaf_135_clk _01150_ VGND VGND VPWR VPWR cpuregs\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12787_ mem_rdata_q\[1\] net12 _01857_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14526_ clknet_leaf_97_clk _00184_ VGND VGND VPWR VPWR cpuregs\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11738_ count_cycle\[4\] _05601_ _05141_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14457_ clknet_leaf_10_clk _00115_ VGND VGND VPWR VPWR cpuregs\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11669_ _05495_ _05246_ _05534_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13408_ net1363 _04835_ _06852_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__mux2_1
X_14388_ clknet_leaf_17_clk _00051_ VGND VGND VPWR VPWR cpuregs\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_626 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_106_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_469 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13339_ _06824_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__clkbuf_1
Xpicorv32_258 VGND VGND VPWR VPWR picorv32_258/HI eoi[4] sky130_fd_sc_hd__conb_1
Xpicorv32_269 VGND VGND VPWR VPWR picorv32_269/HI eoi[15] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_114_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_20_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15009_ clknet_leaf_112_clk _00667_ VGND VGND VPWR VPWR reg_next_pc\[24\] sky130_fd_sc_hd__dfxtp_1
X_07900_ _02030_ _02518_ _02519_ _02008_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__o22a_1
X_08880_ _03359_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07831_ net189 net221 VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__or2b_1
X_07762_ _02018_ _02374_ _02383_ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__o21a_1
X_09501_ decoded_imm\[14\] net176 VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__nand2_1
X_07693_ _02014_ count_cycle\[57\] count_cycle\[25\] _01951_ _02319_ VGND VGND VPWR
+ VPWR _02320_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09432_ _03893_ _03894_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09363_ _02099_ _03828_ _03395_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__mux2_1
X_08314_ _02903_ _02904_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__nor2_1
X_09294_ _03574_ _03751_ _03761_ _03526_ reg_pc\[7\] VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__a32o_1
*XANTENNA_10 _01967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
*XANTENNA_21 _03124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_32 _03201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_43 _03286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08245_ _02290_ net218 _02561_ _02595_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__a31o_1
*XANTENNA_54 _03446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_65 _03586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_76 _03800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_87 _04858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_98 _05948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08176_ _02777_ _02778_ _02418_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput150 net150 VGND VGND VPWR VPWR mem_wdata[23] sky130_fd_sc_hd__buf_2
Xoutput161 net161 VGND VGND VPWR VPWR mem_wdata[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput172 net172 VGND VGND VPWR VPWR pcpi_rs1[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput183 net183 VGND VGND VPWR VPWR pcpi_rs1[20] sky130_fd_sc_hd__buf_2
Xoutput194 net194 VGND VGND VPWR VPWR pcpi_rs1[30] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_902 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_98_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10971_ _04997_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__clkbuf_1
X_12710_ _05912_ _06450_ _06193_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__o21a_1
X_13690_ net1167 _06987_ _06991_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12641_ _05872_ _06384_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15360_ clknet_leaf_68_clk _00950_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dfxtp_1
X_12572_ _06142_ _06318_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14311_ cpuregs\[10\]\[3\] _03201_ _01778_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _05408_ _05409_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15291_ clknet_leaf_78_clk _00883_ VGND VGND VPWR VPWR is_sb_sh_sw sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_740 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire244 net245 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_2
X_14242_ _01746_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__clkbuf_1
X_11454_ decoded_imm_j\[7\] _05204_ _05332_ _05334_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_150_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10405_ _04681_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11385_ _05191_ _05195_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__and2_1
X_14173_ net923 _06923_ _01710_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13124_ net144 net106 _06696_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__mux2_1
X_10336_ _04644_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_13055_ _06665_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__clkbuf_1
X_10267_ net1066 _03228_ _04600_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__mux2_1
X_12006_ net47 net78 _05785_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__mux2_1
X_10198_ _04571_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13957_ net697 _06981_ _01588_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__mux2_1
X_12908_ _06588_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13888_ net1094 _06981_ _01551_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15627_ clknet_leaf_0_clk _01202_ VGND VGND VPWR VPWR cpuregs\[23\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12839_ _06519_ _06526_ _06552_ _06513_ net707 VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__a32o_1
XFILLER_0_158_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_56_320 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_130_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15558_ clknet_leaf_36_clk _01133_ VGND VGND VPWR VPWR cpuregs\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_14509_ clknet_leaf_39_clk _00167_ VGND VGND VPWR VPWR cpuregs\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15489_ clknet_leaf_86_clk _01074_ VGND VGND VPWR VPWR mem_rdata_q\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08030_ _02608_ _02639_ _02640_ _02643_ _02493_ VGND VGND VPWR VPWR alu_out\[6\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_116_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 mem_rdata[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold803 cpuregs\[13\]\[28\] VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_890 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold814 cpuregs\[24\]\[22\] VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold825 cpuregs\[29\]\[5\] VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold836 net59 VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold847 cpuregs\[8\]\[28\] VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 cpuregs\[31\]\[17\] VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 cpuregs\[24\]\[19\] VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _04424_ _04425_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__or3_1
XFILLER_0_149_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08932_ _00013_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08863_ reg_pc\[25\] _03338_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__and2_1
X_07814_ _02432_ _02433_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__nand2_1
X_08794_ reg_pc\[16\] _03279_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07745_ _02366_ _02367_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__xnor2_1
X_07676_ _02300_ _02303_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09415_ cpuregs\[16\]\[11\] cpuregs\[17\]\[11\] cpuregs\[18\]\[11\] cpuregs\[19\]\[11\]
+ _03673_ _03674_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09346_ _00013_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__buf_6
XFILLER_0_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_632 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09277_ _03743_ _03744_ _03579_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08228_ _02397_ _02569_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_745 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_16_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08159_ net178 _02761_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11170_ _05125_ _05123_ net372 _05052_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__a211oi_1
X_10121_ cpuregs\[30\]\[3\] _03202_ _04526_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10052_ cpuregs\[12\]\[4\] _03209_ _04487_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__mux2_1
X_14860_ clknet_leaf_28_clk _00518_ VGND VGND VPWR VPWR cpuregs\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_13811_ _07089_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__clkbuf_1
X_14791_ clknet_leaf_125_clk _00449_ VGND VGND VPWR VPWR cpuregs\[16\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13742_ cpuregs\[29\]\[22\] _06971_ _07050_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__mux2_1
X_10954_ net811 _04873_ _04981_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13673_ _07016_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__clkbuf_1
X_10885_ _04951_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15412_ clknet_leaf_42_clk _01002_ VGND VGND VPWR VPWR cpuregs\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12624_ _05871_ _06367_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__and2_1
X_15343_ clknet_leaf_68_clk _00933_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dfxtp_2
X_12555_ cpuregs\[22\]\[22\] cpuregs\[23\]\[22\] _05816_ VGND VGND VPWR VPWR _06303_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11506_ _05353_ _05362_ _05373_ _05383_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__and4bb_1
X_15274_ clknet_leaf_93_clk _00867_ VGND VGND VPWR VPWR decoded_rd\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12486_ _06023_ _06236_ _05840_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14225_ net793 _06977_ _01732_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__mux2_1
X_11437_ _05258_ net845 _05239_ _05330_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14156_ _01701_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__clkbuf_1
X_11368_ _05263_ net496 _05266_ _05267_ _05257_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_111_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13107_ _06684_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10319_ _04485_ _04522_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__nor2_4
X_14087_ net911 _06975_ _01660_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__mux2_1
X_11299_ _05188_ reg_pc\[13\] VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__or2_1
X_13038_ _06656_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14989_ clknet_leaf_83_clk _00647_ VGND VGND VPWR VPWR reg_next_pc\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_33 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07530_ count_instr\[46\] _01946_ _01947_ count_cycle\[46\] VGND VGND VPWR VPWR _02168_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07461_ _02019_ _02093_ _02103_ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_815 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_57_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_159_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09200_ _03482_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__clkbuf_4
X_07392_ _02037_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09131_ _03418_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09062_ _01854_ _03531_ _03532_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_594 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08013_ _02030_ net249 _02561_ _02563_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold600 cpuregs\[20\]\[16\] VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold611 cpuregs\[16\]\[14\] VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold622 cpuregs\[27\]\[6\] VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 cpuregs\[20\]\[27\] VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold644 cpuregs\[24\]\[24\] VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold655 cpuregs\[27\]\[22\] VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 cpuregs\[3\]\[11\] VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 cpuregs\[16\]\[13\] VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 cpuregs\[30\]\[31\] VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 cpuregs\[16\]\[19\] VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _03455_ _04410_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08915_ instr_sra instr_srai VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_129_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ cpuregs\[16\]\[26\] cpuregs\[17\]\[26\] cpuregs\[18\]\[26\] cpuregs\[19\]\[26\]
+ _03719_ _03450_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_129_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _03330_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08777_ reg_out\[14\] alu_out_q\[14\] _03174_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _02310_ _02328_ _02350_ _02351_ _02335_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_0_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07659_ _02270_ _02274_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10670_ net1089 _04823_ _04819_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_818 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09329_ decoded_imm\[9\] net202 VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_643 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_8_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12340_ cpuregs\[20\]\[13\] cpuregs\[21\]\[13\] _05979_ VGND VGND VPWR VPWR _06097_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12271_ _06022_ _06025_ _06028_ _06030_ _03080_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__a221o_2
XFILLER_0_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14010_ _01601_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__buf_4
X_11222_ _05162_ _05163_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11153_ _05115_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__clkbuf_1
X_10104_ cpuregs\[12\]\[29\] _03374_ _04509_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11084_ count_instr\[12\] _05065_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__or2_1
X_15961_ clknet_leaf_139_clk _01533_ VGND VGND VPWR VPWR cpuregs\[10\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14912_ clknet_leaf_119_clk _00570_ VGND VGND VPWR VPWR count_instr\[21\] sky130_fd_sc_hd__dfxtp_1
X_10035_ _02380_ _03486_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__and2_1
X_15892_ clknet_leaf_16_clk _01464_ VGND VGND VPWR VPWR cpuregs\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_14843_ clknet_leaf_160_clk _00501_ VGND VGND VPWR VPWR cpuregs\[20\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14774_ clknet_leaf_158_clk _00432_ VGND VGND VPWR VPWR cpuregs\[16\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ _05779_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_595 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13725_ net659 _06954_ _07039_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10937_ net1048 _04856_ _04970_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13656_ _07007_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__clkbuf_1
X_10868_ _04942_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12607_ _06058_ _06351_ _06182_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13587_ cpuregs\[31\]\[19\] _06964_ _06946_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10799_ cpuregs\[16\]\[17\] _04854_ _04898_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15326_ clknet_leaf_58_clk _00916_ VGND VGND VPWR VPWR cpuregs\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12538_ cpuregs\[6\]\[22\] cpuregs\[7\]\[22\] _03084_ VGND VGND VPWR VPWR _06286_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15257_ clknet_leaf_112_clk _00850_ VGND VGND VPWR VPWR instr_rdcycleh sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12469_ cpuregs\[16\]\[18\] cpuregs\[17\]\[18\] cpuregs\[18\]\[18\] cpuregs\[19\]\[18\]
+ _05921_ _05985_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14208_ net1230 _06960_ _01721_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15188_ clknet_leaf_71_clk alu_out\[1\] VGND VGND VPWR VPWR alu_out_q\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14139_ _01692_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08700_ _03203_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__clkbuf_1
X_09680_ _03473_ _04126_ _04135_ _03526_ reg_pc\[19\] VGND VGND VPWR VPWR _04136_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_146_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08631_ _03045_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08562_ _03054_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07513_ _02134_ _02136_ _02133_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_155_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_155_clk sky130_fd_sc_hd__clkbuf_2
X_08493_ decoded_imm_j\[15\] _01077_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__mux2_1
X_07444_ count_instr\[8\] instr_rdinstr count_cycle\[8\] _01950_ VGND VGND VPWR VPWR
+ _02088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07375_ net1413 _02013_ count_cycle\[5\] _02020_ _02021_ VGND VGND VPWR VPWR _02022_
+ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_40_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09114_ _00012_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__buf_8
XFILLER_0_115_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09045_ _03493_ _03515_ _03518_ _03415_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold430 cpuregs\[30\]\[20\] VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 cpuregs\[31\]\[24\] VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 cpuregs\[20\]\[26\] VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 cpuregs\[17\]\[26\] VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 cpuregs\[26\]\[24\] VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 cpuregs\[11\]\[22\] VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 cpuregs\[31\]\[9\] VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__dlygate4sd3_1
X_09947_ _02340_ _03770_ _04328_ _03670_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_5_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _02449_ _03770_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__nor2_1
X_08829_ net617 _03314_ _03315_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__mux2_1
X_11840_ net501 count_cycle\[35\] count_cycle\[36\] _05667_ VGND VGND VPWR VPWR _05673_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_67_212 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_95_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11771_ count_cycle\[13\] _05620_ count_cycle\[14\] VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_146_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_146_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_138_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13510_ cpuregs\[9\]\[24\] _04869_ _06910_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__mux2_1
X_10722_ net692 _04858_ _04840_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_716 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14490_ clknet_leaf_5_clk _00148_ VGND VGND VPWR VPWR cpuregs\[30\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_749 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_604 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13441_ _06878_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_492 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10653_ net1059 _03367_ _04804_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13372_ net1372 _04867_ _06838_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__mux2_1
X_10584_ _04776_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__clkbuf_1
X_15111_ clknet_leaf_103_clk _07135_ VGND VGND VPWR VPWR reg_out\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12323_ cpuregs\[4\]\[13\] cpuregs\[5\]\[13\] _03062_ VGND VGND VPWR VPWR _06080_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_575 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15042_ clknet_leaf_120_clk _00700_ VGND VGND VPWR VPWR count_cycle\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12254_ _03037_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_75_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11205_ _01884_ _05150_ _05151_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12185_ _03051_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__buf_8
X_11136_ net534 _05100_ _05090_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__o21ai_1
X_11067_ count_instr\[7\] count_instr\[6\] _05051_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__and3_1
X_15944_ clknet_leaf_36_clk _01516_ VGND VGND VPWR VPWR cpuregs\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_10018_ cpuregs\[20\]\[30\] cpuregs\[21\]\[30\] cpuregs\[22\]\[30\] cpuregs\[23\]\[30\]
+ _03673_ _03674_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__mux4_1
X_15875_ clknet_leaf_51_clk _01447_ VGND VGND VPWR VPWR cpuregs\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ clknet_leaf_54_clk _00484_ VGND VGND VPWR VPWR cpuregs\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_14757_ clknet_leaf_150_clk _00415_ VGND VGND VPWR VPWR cpuregs\[26\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_137_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_137_clk sky130_fd_sc_hd__clkbuf_2
X_11969_ _05770_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__clkbuf_1
X_13708_ net991 _06937_ _07028_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_127_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14688_ clknet_leaf_147_clk _00346_ VGND VGND VPWR VPWR cpuregs\[27\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13639_ _06998_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_486 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_816 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07160_ instr_sb instr_lw instr_lh instr_jalr VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__or4_1
XFILLER_0_143_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15309_ clknet_leaf_18_clk _00899_ VGND VGND VPWR VPWR cpuregs\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_136_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09801_ cpuregs\[20\]\[23\] cpuregs\[21\]\[23\] cpuregs\[22\]\[23\] cpuregs\[23\]\[23\]
+ _03516_ _03409_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07993_ net97 net108 net251 net119 VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__or4_4
X_09732_ _04184_ _04185_ _03552_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__mux2_1
X_09663_ cpuregs\[4\]\[19\] cpuregs\[5\]\[19\] cpuregs\[6\]\[19\] cpuregs\[7\]\[19\]
+ _03808_ _03801_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__mux4_1
X_08614_ _03045_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__clkbuf_8
X_09594_ decoded_imm\[17\] _02213_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__nand2_1
X_08545_ _03061_ _03064_ _03034_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_128_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_128_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08476_ _03010_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_1
XFILLER_0_92_513 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_453 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07427_ _02058_ _02064_ _02070_ _02071_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_21_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07358_ _02001_ _02004_ _02005_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07289_ net1 net130 _01938_ _01940_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__a22o_1
X_09028_ _03403_ _03491_ _03501_ _03420_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_130_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold260 net164 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 count_cycle\[38\] VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold282 cpuregs\[23\]\[1\] VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 instr_sh VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13990_ cpuregs\[5\]\[10\] _06945_ _01613_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__mux2_1
X_12941_ _06605_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15660_ clknet_leaf_143_clk _01235_ VGND VGND VPWR VPWR cpuregs\[29\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_100 _05984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12872_ is_alu_reg_reg _06528_ net242 VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__and3_1
*XANTENNA_111 mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_122 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14611_ clknet_leaf_30_clk _00269_ VGND VGND VPWR VPWR cpuregs\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11823_ net507 _05658_ _05647_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__o21ai_1
*XANTENNA_133 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_119_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_119_clk sky130_fd_sc_hd__clkbuf_2
*XANTENNA_144 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15591_ clknet_leaf_55_clk _01166_ VGND VGND VPWR VPWR cpuregs\[31\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_908 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_155 _03045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_166 _03449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
*XANTENNA_177 _04782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14542_ clknet_leaf_43_clk _00200_ VGND VGND VPWR VPWR cpuregs\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11754_ count_cycle\[9\] _05611_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_188 _05886_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_199 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _04847_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__clkbuf_1
X_14473_ clknet_leaf_59_clk _00131_ VGND VGND VPWR VPWR cpuregs\[12\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11685_ _05263_ _05558_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13424_ _06869_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__clkbuf_1
X_10636_ _04781_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_529 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13355_ cpuregs\[19\]\[15\] _04850_ _06827_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10567_ _04767_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ _05879_ _06057_ _06060_ _06063_ _03104_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__a221o_2
X_13286_ _06796_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10498_ _04730_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__clkbuf_1
X_15025_ clknet_leaf_113_clk _00683_ VGND VGND VPWR VPWR count_cycle\[8\] sky130_fd_sc_hd__dfxtp_1
X_12237_ _03106_ _05997_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__or2_1
X_12168_ _03052_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__buf_4
X_11119_ count_instr\[22\] count_instr\[21\] _05087_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__and3_1
X_12099_ _05866_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__clkbuf_1
X_15927_ clknet_leaf_133_clk _01499_ VGND VGND VPWR VPWR cpuregs\[0\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xinput6 net460 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_88_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15858_ clknet_leaf_6_clk _01430_ VGND VGND VPWR VPWR cpuregs\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14809_ clknet_leaf_160_clk _00467_ VGND VGND VPWR VPWR cpuregs\[25\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15789_ clknet_leaf_142_clk _01364_ VGND VGND VPWR VPWR cpuregs\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08330_ _02394_ _02918_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_604 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08261_ _02849_ _02855_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07212_ cpu_state\[1\] net34 VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__nand2_4
XFILLER_0_160_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08192_ net213 _02792_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__xor2_2
XFILLER_0_116_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_144_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_796 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_65_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07976_ _01978_ _02509_ _02593_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__a21oi_1
X_09715_ cpuregs\[4\]\[20\] cpuregs\[5\]\[20\] cpuregs\[6\]\[20\] cpuregs\[7\]\[20\]
+ _03457_ _03464_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09646_ cpuregs\[12\]\[18\] cpuregs\[13\]\[18\] cpuregs\[14\]\[18\] cpuregs\[15\]\[18\]
+ _03582_ _03716_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_153_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09577_ cpuregs\[24\]\[16\] cpuregs\[25\]\[16\] cpuregs\[26\]\[16\] cpuregs\[27\]\[16\]
+ _03636_ _03637_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08528_ cpuregs\[24\]\[2\] cpuregs\[25\]\[2\] cpuregs\[26\]\[2\] cpuregs\[27\]\[2\]
+ _03046_ _03047_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_139_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08459_ _02998_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_108_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11470_ _05360_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10421_ net872 _03282_ _04684_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_752 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13140_ _06713_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10352_ cpuregs\[28\]\[15\] _03282_ _04647_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13071_ _05766_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10283_ _04616_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__clkbuf_1
X_12022_ net56 net87 _05766_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13973_ cpuregs\[5\]\[2\] _06929_ _01602_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__mux2_1
X_12924_ decoded_imm_j\[8\] _01090_ _03169_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__mux2_1
X_15712_ clknet_leaf_53_clk _01287_ VGND VGND VPWR VPWR cpuregs\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15643_ clknet_leaf_129_clk _01218_ VGND VGND VPWR VPWR cpuregs\[23\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12855_ _06532_ _06536_ _06533_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__nor3_1
XFILLER_0_29_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11806_ _05649_ _05650_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_83_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15574_ clknet_leaf_140_clk _01149_ VGND VGND VPWR VPWR cpuregs\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _06516_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__clkbuf_1
X_14525_ clknet_leaf_13_clk _00183_ VGND VGND VPWR VPWR cpuregs\[13\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11737_ _05601_ _05602_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_710 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_126_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_911 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14456_ clknet_leaf_17_clk _00114_ VGND VGND VPWR VPWR cpuregs\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11668_ _05494_ _05249_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_12_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _06860_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__clkbuf_1
X_10619_ _04795_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14387_ clknet_leaf_13_clk _00050_ VGND VGND VPWR VPWR cpuregs\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11599_ _05031_ reg_next_pc\[20\] VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13338_ cpuregs\[19\]\[7\] _04833_ _06816_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpicorv32_259 VGND VGND VPWR VPWR picorv32_259/HI eoi[5] sky130_fd_sc_hd__conb_1
X_13269_ _06787_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15008_ clknet_leaf_110_clk _00666_ VGND VGND VPWR VPWR reg_next_pc\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07830_ net190 VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07761_ _01970_ _02379_ _02382_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__a21o_1
X_09500_ decoded_imm\[14\] net176 VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__or2_1
X_07692_ count_instr\[57\] instr_rdinstrh _01949_ count_instr\[25\] VGND VGND VPWR
+ VPWR _02319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09431_ decoded_imm\[12\] net174 VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_96 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09362_ _03651_ _03798_ _03799_ _03823_ _03827_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__a311o_1
XFILLER_0_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08313_ _02369_ _02901_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09293_ _03753_ _03755_ _03757_ _03759_ _03760_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_11 _01967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_22 _03134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_33 _03208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08244_ _02290_ net218 _02593_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_229 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_44 _03286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_55 _03446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_66 _03588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_77 _03801_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_88 _04875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08175_ _02417_ _02568_ _02595_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
*XANTENNA_99 _05969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput140 net140 VGND VGND VPWR VPWR mem_wdata[14] sky130_fd_sc_hd__clkbuf_4
Xoutput151 net151 VGND VGND VPWR VPWR mem_wdata[24] sky130_fd_sc_hd__clkbuf_4
Xoutput162 net162 VGND VGND VPWR VPWR mem_wdata[5] sky130_fd_sc_hd__clkbuf_4
Xoutput173 net173 VGND VGND VPWR VPWR pcpi_rs1[11] sky130_fd_sc_hd__clkbuf_4
Xoutput184 net184 VGND VGND VPWR VPWR pcpi_rs1[21] sky130_fd_sc_hd__buf_2
Xoutput195 net252 VGND VGND VPWR VPWR pcpi_rs1[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07959_ _02576_ _02577_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10970_ net655 _04821_ _04995_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__mux2_1
X_09629_ _04082_ _04055_ _04085_ _04052_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_468 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ cpuregs\[20\]\[26\] cpuregs\[21\]\[26\] _05979_ VGND VGND VPWR VPWR _06384_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12571_ cpuregs\[20\]\[23\] cpuregs\[21\]\[23\] cpuregs\[22\]\[23\] cpuregs\[23\]\[23\]
+ _06065_ _03144_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_50_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_93_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14310_ _01781_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__clkbuf_1
X_11522_ decoded_imm_j\[14\] _05219_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15290_ clknet_leaf_78_clk _00882_ VGND VGND VPWR VPWR is_jalr_addi_slti_sltiu_xori_ori_andi
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_702 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire245 _03117_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_2
X_14241_ net606 VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11453_ decoded_imm_j\[9\] _05208_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10404_ net888 _03228_ _04673_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14172_ _01709_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__buf_6
X_11384_ _05191_ _05195_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13123_ _06704_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10335_ net1309 _03228_ _04636_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13054_ net711 _04873_ _06658_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__mux2_1
X_10266_ _04607_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__clkbuf_1
X_12005_ _05789_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10197_ net893 _03221_ _04564_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13956_ _01595_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12907_ decoded_imm_j\[4\] _01086_ _06587_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__mux2_1
X_13887_ _01558_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ clknet_leaf_1_clk _01201_ VGND VGND VPWR VPWR cpuregs\[23\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12838_ _01074_ _01075_ _01076_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__nor3_1
XFILLER_0_29_535 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_389 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_56_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15557_ clknet_leaf_27_clk _01132_ VGND VGND VPWR VPWR cpuregs\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12769_ _01970_ _05185_ _01894_ _03176_ _01843_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14508_ clknet_leaf_23_clk _00166_ VGND VGND VPWR VPWR cpuregs\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15488_ clknet_leaf_93_clk _01073_ VGND VGND VPWR VPWR mem_rdata_q\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_25_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_613 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput20 net426 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_116_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_201 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14439_ clknet_leaf_95_clk _00097_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dfxtp_1
Xinput31 net428 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_130_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold804 cpuregs\[5\]\[22\] VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 cpuregs\[22\]\[6\] VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold826 cpuregs\[10\]\[30\] VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold837 cpuregs\[12\]\[27\] VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold848 cpuregs\[2\]\[26\] VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09980_ _04399_ _04400_ _04401_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__o21a_1
Xhold859 cpuregs\[3\]\[3\] VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08931_ _03405_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08862_ reg_pc\[25\] _03338_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__nor2_1
X_07813_ net190 net222 VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__or2_1
X_08793_ reg_out\[16\] alu_out_q\[16\] _03175_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07744_ _02353_ _02356_ _02355_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_144_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07675_ _02301_ _02302_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09414_ _03647_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09345_ _03547_ _03804_ _03806_ _03810_ _03489_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_32_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_90_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09276_ cpuregs\[0\]\[7\] cpuregs\[1\]\[7\] cpuregs\[2\]\[7\] cpuregs\[3\]\[7\] _03439_
+ _03450_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_43_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08227_ _02277_ net217 _02598_ _02641_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08158_ net178 _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08089_ _02696_ _02697_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10120_ _04529_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_99_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_2
X_10051_ _04491_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13810_ net1321 _06971_ _07086_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__mux2_1
X_14790_ clknet_leaf_126_clk _00448_ VGND VGND VPWR VPWR cpuregs\[16\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_13741_ _07052_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10953_ _04987_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13672_ cpuregs\[23\]\[21\] _06969_ _07014_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__mux2_1
X_10884_ net802 _04871_ _04945_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12623_ cpuregs\[4\]\[26\] cpuregs\[5\]\[26\] _03051_ VGND VGND VPWR VPWR _06367_
+ sky130_fd_sc_hd__mux2_1
X_15411_ clknet_leaf_37_clk _01001_ VGND VGND VPWR VPWR cpuregs\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_155_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_81_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_93_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15342_ clknet_leaf_68_clk _00932_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dfxtp_1
X_12554_ _05872_ _06301_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_551 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_124_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11505_ _05391_ _05392_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15273_ clknet_leaf_93_clk _00866_ VGND VGND VPWR VPWR decoded_rd\[0\] sky130_fd_sc_hd__dfxtp_1
X_12485_ cpuregs\[16\]\[19\] cpuregs\[17\]\[19\] cpuregs\[18\]\[19\] cpuregs\[19\]\[19\]
+ _05948_ _06068_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__mux4_1
XFILLER_0_123_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_532 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14224_ _01737_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__clkbuf_1
X_11436_ _05269_ _05325_ _05326_ _05329_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14155_ net1231 _06975_ _01696_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11367_ _05187_ _05265_ _05193_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13106_ _06695_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _04634_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__clkbuf_1
X_14086_ _01664_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__clkbuf_1
X_11298_ reg_next_pc\[13\] _03265_ _02946_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__mux2_2
XFILLER_0_119_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13037_ cpuregs\[1\]\[18\] _04856_ _06647_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__mux2_1
X_10249_ cpuregs\[13\]\[31\] _03386_ _04563_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14988_ clknet_leaf_83_clk _00646_ VGND VGND VPWR VPWR reg_next_pc\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13939_ _01586_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__clkbuf_1
X_07460_ _02058_ _02098_ _02102_ _02071_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_827 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_119_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15609_ clknet_leaf_144_clk _01184_ VGND VGND VPWR VPWR cpuregs\[31\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_07391_ reg_pc\[6\] decoded_imm\[6\] VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_14_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_2
X_09130_ cpuregs\[28\]\[3\] cpuregs\[29\]\[3\] cpuregs\[30\]\[3\] cpuregs\[31\]\[3\]
+ _03601_ _03492_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09061_ _03482_ _03533_ _03534_ _01953_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08012_ _02621_ _02626_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__xnor2_1
Xhold601 cpuregs\[10\]\[18\] VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold612 cpuregs\[9\]\[17\] VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 cpuregs\[19\]\[0\] VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 cpuregs\[2\]\[9\] VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 cpuregs\[5\]\[9\] VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 cpuregs\[21\]\[11\] VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold667 cpuregs\[10\]\[5\] VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09963_ cpuregs\[12\]\[28\] cpuregs\[13\]\[28\] cpuregs\[14\]\[28\] cpuregs\[15\]\[28\]
+ _03458_ _03461_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__mux4_1
Xhold678 cpuregs\[14\]\[8\] VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 cpuregs\[20\]\[18\] VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ cpu_state\[2\] cpu_state\[4\] VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09894_ cpuregs\[20\]\[26\] cpuregs\[21\]\[26\] cpuregs\[22\]\[26\] cpuregs\[23\]\[26\]
+ _03587_ _03588_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_129_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ net844 _03329_ _03315_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__mux2_1
X_08776_ _03269_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__clkbuf_1
X_07727_ _02326_ _02336_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_0_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_427 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07658_ _02285_ _02286_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
X_07589_ net10 _02202_ _02180_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__a21o_1
X_09328_ decoded_imm\[9\] net202 VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_655 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_145_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_793 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09259_ cpuregs\[0\]\[6\] cpuregs\[1\]\[6\] cpuregs\[2\]\[6\] cpuregs\[3\]\[6\] _03719_
+ _03450_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12270_ _03149_ _06029_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11221_ net511 _05160_ _05133_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11152_ _05112_ _05113_ _05114_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__and3b_1
X_10103_ _04518_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__clkbuf_1
X_11083_ _05065_ _05066_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__nor2_1
X_15960_ clknet_leaf_141_clk _01532_ VGND VGND VPWR VPWR cpuregs\[10\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14911_ clknet_leaf_119_clk _00569_ VGND VGND VPWR VPWR count_instr\[20\] sky130_fd_sc_hd__dfxtp_1
X_10034_ reg_pc\[30\] _03528_ _04478_ _03626_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__a211o_1
X_15891_ clknet_leaf_5_clk _01463_ VGND VGND VPWR VPWR cpuregs\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14842_ clknet_leaf_160_clk _00500_ VGND VGND VPWR VPWR cpuregs\[20\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14773_ clknet_leaf_159_clk _00431_ VGND VGND VPWR VPWR cpuregs\[16\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11985_ net37 net68 _05774_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_574 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_85_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10936_ _04978_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__clkbuf_1
X_13724_ _07043_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__clkbuf_1
X_13655_ net1342 _06952_ _07003_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__mux2_1
X_10867_ net966 _04854_ _04934_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12606_ cpuregs\[12\]\[25\] cpuregs\[13\]\[25\] cpuregs\[14\]\[25\] cpuregs\[15\]\[25\]
+ _03133_ _03134_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13586_ _03306_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__buf_2
X_10798_ _04905_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15325_ clknet_leaf_133_clk _00915_ VGND VGND VPWR VPWR cpuregs\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12537_ _05871_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_595 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_880 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12468_ _03087_ _06219_ _03153_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__a21o_1
X_15256_ clknet_leaf_87_clk _00849_ VGND VGND VPWR VPWR instr_rdcycle sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_151_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14207_ _01728_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_93_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11419_ decoded_imm_j\[6\] _05201_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_93_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15187_ clknet_leaf_71_clk alu_out\[0\] VGND VGND VPWR VPWR alu_out_q\[0\] sky130_fd_sc_hd__dfxtp_1
X_12399_ _06132_ _06141_ _06152_ _06153_ decoded_imm\[15\] VGND VGND VPWR VPWR _06154_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14138_ net848 _06958_ _01685_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14069_ _01655_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_3_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_2
X_08630_ _03143_ _03145_ _03147_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08561_ _03033_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07512_ _02149_ _02150_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08492_ _03021_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__buf_4
XFILLER_0_159_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07443_ count_instr\[40\] instr_rdinstrh instr_rdcycleh count_cycle\[40\] VGND VGND
+ VPWR VPWR _02087_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07374_ count_instr\[5\] _01965_ count_cycle\[37\] _02014_ VGND VGND VPWR VPWR _02021_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09113_ _03581_ _03584_ _03467_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_40_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_463 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_115_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09044_ _03410_ _03517_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold420 count_cycle\[7\] VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 cpuregs\[11\]\[10\] VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold442 cpuregs\[5\]\[17\] VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 net58 VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 cpuregs\[19\]\[24\] VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 cpuregs\[25\]\[15\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 reg_next_pc\[7\] VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 cpuregs\[26\]\[31\] VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__dlygate4sd3_1
X_09946_ _04329_ _04392_ _03670_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_55_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _03475_ _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__and2_1
X_08828_ _03184_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08759_ _03254_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11770_ _01839_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_544 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_49_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10721_ _03306_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ cpuregs\[24\]\[23\] _04867_ _06874_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__mux2_1
X_10652_ _04812_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_97_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_860 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_178 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13371_ _06841_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__clkbuf_1
X_10583_ net1254 _03360_ _04768_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_880 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_134_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15110_ clknet_leaf_103_clk _07134_ VGND VGND VPWR VPWR reg_out\[28\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12322_ _06079_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_39_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15041_ clknet_leaf_122_clk _00699_ VGND VGND VPWR VPWR count_cycle\[24\] sky130_fd_sc_hd__dfxtp_1
X_12253_ cpuregs\[0\]\[10\] cpuregs\[1\]\[10\] cpuregs\[2\]\[10\] cpuregs\[3\]\[10\]
+ _05908_ _05909_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_75_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11204_ net1401 _05148_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12184_ _03143_ _05946_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__or2_1
X_11135_ count_instr\[27\] count_instr\[26\] _05095_ _05098_ VGND VGND VPWR VPWR _05103_
+ sky130_fd_sc_hd__and4_1
X_11066_ _05053_ _05054_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__nor2_1
X_15943_ clknet_leaf_38_clk _01515_ VGND VGND VPWR VPWR cpuregs\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_10017_ cpuregs\[16\]\[30\] cpuregs\[17\]\[30\] cpuregs\[18\]\[30\] cpuregs\[19\]\[30\]
+ _03673_ _03674_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15874_ clknet_leaf_51_clk _01446_ VGND VGND VPWR VPWR cpuregs\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14825_ clknet_leaf_19_clk _00483_ VGND VGND VPWR VPWR cpuregs\[25\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14756_ clknet_leaf_150_clk _00414_ VGND VGND VPWR VPWR cpuregs\[26\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11968_ net1195 net90 _05767_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13707_ _07034_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10919_ _04969_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__clkbuf_1
X_14687_ clknet_leaf_128_clk _00345_ VGND VGND VPWR VPWR cpuregs\[27\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_11899_ _05706_ _05713_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13638_ cpuregs\[23\]\[5\] _06935_ _06992_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13569_ net1161 _06952_ _06946_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_828 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_143_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_699 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_125_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15308_ clknet_leaf_8_clk _00898_ VGND VGND VPWR VPWR cpuregs\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15239_ clknet_leaf_76_clk _00832_ VGND VGND VPWR VPWR instr_xori sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_382 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09800_ _03427_ _04247_ _04249_ _04251_ _03591_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__a221o_1
X_07992_ net240 VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09731_ cpuregs\[0\]\[21\] cpuregs\[1\]\[21\] cpuregs\[2\]\[21\] cpuregs\[3\]\[21\]
+ _03800_ _03407_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09662_ _04116_ _04117_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__xnor2_1
X_08613_ _03128_ _03130_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__nor2_1
X_09593_ _03396_ _04032_ _04050_ _04051_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_49_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08544_ cpuregs\[0\]\[2\] cpuregs\[1\]\[2\] cpuregs\[2\]\[2\] cpuregs\[3\]\[2\] _03062_
+ _03063_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__mux4_1
XFILLER_0_159_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08475_ net253 _03009_ _02993_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_622 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07426_ _01955_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07357_ _02001_ _02004_ _01945_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07288_ _01939_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09027_ _03493_ _03495_ _03499_ _03500_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold250 cpuregs\[3\]\[0\] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold261 cpuregs\[17\]\[8\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold272 cpuregs\[28\]\[21\] VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 cpuregs\[9\]\[10\] VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 cpuregs\[14\]\[2\] VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09929_ _03436_ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12940_ decoded_imm_j\[19\] _01081_ _06587_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _06546_ _06565_ _06566_ _06562_ instr_sub VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__a32o_1
*XANTENNA_101 _06761_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_112 mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14610_ clknet_leaf_55_clk _00268_ VGND VGND VPWR VPWR cpuregs\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_123 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11822_ count_cycle\[28\] count_cycle\[29\] count_cycle\[30\] _05655_ VGND VGND VPWR
+ VPWR _05661_ sky130_fd_sc_hd__and4_4
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_134 net212 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15590_ clknet_leaf_35_clk _01165_ VGND VGND VPWR VPWR cpuregs\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_145 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_156 _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_167 _03449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11753_ count_cycle\[7\] count_cycle\[8\] count_cycle\[9\] _05607_ VGND VGND VPWR
+ VPWR _05613_ sky130_fd_sc_hd__and4_4
*XANTENNA_178 _04782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14541_ clknet_leaf_39_clk _00199_ VGND VGND VPWR VPWR cpuregs\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_189 _05925_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10704_ net1075 _04846_ _04840_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _01903_ _05548_ _05556_ _05264_ _05557_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__a221o_1
X_14472_ clknet_leaf_59_clk _00130_ VGND VGND VPWR VPWR cpuregs\[12\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_37_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13423_ net1219 _04850_ _06863_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__mux2_1
X_10635_ _04803_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13354_ _06832_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_800 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10566_ net657 _03307_ _04757_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12305_ _03106_ _06062_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__or2_1
X_13285_ net1107 _04848_ _06791_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_488 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10497_ net782 _03307_ _04720_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__mux2_1
X_15024_ clknet_leaf_113_clk _00682_ VGND VGND VPWR VPWR count_cycle\[7\] sky130_fd_sc_hd__dfxtp_1
X_12236_ cpuregs\[8\]\[9\] cpuregs\[9\]\[9\] cpuregs\[10\]\[9\] cpuregs\[11\]\[9\]
+ _03150_ _05917_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_20_875 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12167_ _03083_ _05930_ _03081_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__o21a_1
X_11118_ _05089_ _05091_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__nor2_1
X_12098_ _02509_ _05865_ _05863_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15926_ clknet_leaf_145_clk _01498_ VGND VGND VPWR VPWR cpuregs\[0\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_11049_ count_instr\[2\] net994 _05041_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 mem_rdata[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_88_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ clknet_leaf_9_clk _01429_ VGND VGND VPWR VPWR cpuregs\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14808_ clknet_leaf_153_clk _00466_ VGND VGND VPWR VPWR cpuregs\[25\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15788_ clknet_leaf_16_clk _01363_ VGND VGND VPWR VPWR cpuregs\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14739_ clknet_leaf_29_clk _00397_ VGND VGND VPWR VPWR cpuregs\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_46_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08260_ _02849_ _02855_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07211_ _01865_ _01873_ _01875_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08191_ _02656_ _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07975_ instr_xor instr_xori VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__nor2_4
X_09714_ _03746_ _04168_ _03467_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__o21a_1
X_09645_ _03433_ _04097_ _04099_ _04101_ _03760_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__a221o_1
X_09576_ _04033_ _04034_ _03414_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08527_ _00008_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08458_ _02290_ _02997_ _02993_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07409_ _01949_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__buf_4
XFILLER_0_80_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08389_ reg_next_pc\[2\] reg_out\[2\] _02949_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10420_ _04689_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_764 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10351_ _04652_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13070_ _02951_ _05767_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__nand2_1
X_10282_ cpuregs\[2\]\[14\] _03275_ _04611_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12021_ _05797_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13972_ _01604_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__clkbuf_1
X_15711_ clknet_leaf_54_clk _01286_ VGND VGND VPWR VPWR cpuregs\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12923_ _06596_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_103_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15642_ clknet_leaf_153_clk _01217_ VGND VGND VPWR VPWR cpuregs\[23\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12854_ _06546_ _06534_ _06559_ _06530_ net440 VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__a32o_1
X_11805_ net797 _05646_ _05647_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15573_ clknet_leaf_140_clk _01148_ VGND VGND VPWR VPWR cpuregs\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12785_ mem_rdata_q\[0\] net1 _01857_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14524_ clknet_leaf_18_clk _00182_ VGND VGND VPWR VPWR cpuregs\[13\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11736_ net528 _05598_ _05169_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_154_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14455_ clknet_leaf_13_clk _00113_ VGND VGND VPWR VPWR cpuregs\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_923 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11667_ _05249_ _05528_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ net1201 _04833_ _06852_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10618_ cpuregs\[15\]\[11\] _03255_ _04793_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__mux2_1
X_14386_ clknet_leaf_15_clk _00049_ VGND VGND VPWR VPWR cpuregs\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11598_ _05235_ _05478_ _05300_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10549_ _04758_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13337_ _06823_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13268_ cpuregs\[18\]\[6\] _04831_ _06780_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15007_ clknet_leaf_112_clk _00665_ VGND VGND VPWR VPWR reg_next_pc\[22\] sky130_fd_sc_hd__dfxtp_1
X_12219_ _05872_ _05980_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13199_ net574 _06742_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07760_ _02065_ _02380_ _02201_ _02381_ _01955_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__a221o_1
X_15909_ clknet_leaf_39_clk _01481_ VGND VGND VPWR VPWR cpuregs\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_07691_ _01977_ _02316_ _02201_ _02317_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__a22o_1
X_09430_ decoded_imm\[12\] net174 VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09361_ _03616_ _03825_ _03826_ _01942_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__o211a_1
X_08312_ _02902_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__inv_2
X_09292_ _03430_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_12 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_901 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_23 _03137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08243_ _02838_ _02839_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__xnor2_1
*XANTENNA_34 _03208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_45 _03295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_457 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_56 _03474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_67 _03588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_78 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08174_ _02213_ net211 _02618_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_134_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_89 _04886_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput130 net130 VGND VGND VPWR VPWR mem_la_wstrb[0] sky130_fd_sc_hd__buf_2
Xoutput141 net141 VGND VGND VPWR VPWR mem_wdata[15] sky130_fd_sc_hd__clkbuf_4
Xoutput152 net152 VGND VGND VPWR VPWR mem_wdata[25] sky130_fd_sc_hd__buf_2
XFILLER_0_11_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput163 net163 VGND VGND VPWR VPWR mem_wdata[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput174 net174 VGND VGND VPWR VPWR pcpi_rs1[12] sky130_fd_sc_hd__clkbuf_4
Xoutput185 net185 VGND VGND VPWR VPWR pcpi_rs1[22] sky130_fd_sc_hd__buf_2
Xoutput196 net196 VGND VGND VPWR VPWR pcpi_rs1[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_149_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07958_ net182 _02574_ _02575_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__or3_1
X_07889_ net119 VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__clkbuf_4
X_09628_ _04083_ _04084_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ _03895_ _03930_ _03963_ _04012_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_65_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_322 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12570_ _06177_ _06312_ _06314_ _06316_ _06164_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11521_ _05407_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_347 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11452_ net361 _05208_ _05338_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__and3_1
X_14240_ _01745_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10403_ _04680_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__clkbuf_1
X_14171_ _03180_ _04485_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__nor2_2
XFILLER_0_116_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11383_ _05280_ _05272_ _05278_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__a21bo_1
X_13122_ net143 net105 _06696_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10334_ _04643_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__clkbuf_1
X_13053_ _06664_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__clkbuf_1
X_10265_ net996 _03221_ _04600_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__mux2_1
X_12004_ net761 net77 _05785_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10196_ _04570_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_21_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13955_ net921 _06979_ _01588_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__mux2_1
X_12906_ _03021_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__buf_4
X_13886_ cpuregs\[22\]\[26\] _06979_ _01551_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ clknet_leaf_0_clk _01200_ VGND VGND VPWR VPWR cpuregs\[23\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12837_ _06551_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__buf_1
XFILLER_0_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15556_ clknet_leaf_38_clk _01131_ VGND VGND VPWR VPWR cpuregs\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_344 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12768_ latched_store _01888_ _06502_ _06505_ _05358_ VGND VGND VPWR VPWR _00806_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14507_ clknet_leaf_56_clk _00165_ VGND VGND VPWR VPWR cpuregs\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11719_ _05261_ _05584_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__or2_1
X_15487_ clknet_leaf_93_clk _01072_ VGND VGND VPWR VPWR mem_rdata_q\[10\] sky130_fd_sc_hd__dfxtp_1
X_12699_ _06438_ _06439_ _03082_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput10 net416 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
X_14438_ clknet_leaf_96_clk _00096_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_116_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_625 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xinput21 net423 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_116_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput32 net424 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_126_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_40_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14369_ net1208 _03385_ _01777_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__mux2_1
Xhold805 cpuregs\[12\]\[9\] VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 cpuregs\[18\]\[10\] VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 cpuregs\[31\]\[18\] VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold838 cpuregs\[2\]\[20\] VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold849 cpuregs\[10\]\[31\] VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08930_ _03404_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__buf_8
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08861_ reg_out\[25\] alu_out_q\[25\] _03176_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__mux2_1
X_07812_ net190 net222 VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__nand2_1
X_08792_ _03283_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__clkbuf_1
X_07743_ _02364_ _02365_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07674_ reg_pc\[24\] decoded_imm\[24\] VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_144_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09413_ cpuregs\[20\]\[11\] cpuregs\[21\]\[11\] cpuregs\[22\]\[11\] cpuregs\[23\]\[11\]
+ _03516_ _03674_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09344_ _03807_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09275_ cpuregs\[4\]\[7\] cpuregs\[5\]\[7\] cpuregs\[6\]\[7\] cpuregs\[7\]\[7\] _03439_
+ _03450_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08226_ _02608_ _02820_ _02821_ _02824_ VGND VGND VPWR VPWR alu_out\[21\] sky130_fd_sc_hd__a31o_2
XFILLER_0_145_574 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08157_ net247 _02760_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08088_ _02680_ _02687_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10050_ cpuregs\[12\]\[3\] _03202_ _04487_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13740_ cpuregs\[29\]\[21\] _06969_ _07050_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10952_ cpuregs\[20\]\[25\] _04871_ _04981_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13671_ _07015_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__clkbuf_1
X_10883_ _04950_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15410_ clknet_leaf_29_clk _01000_ VGND VGND VPWR VPWR cpuregs\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12622_ _06366_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15341_ clknet_leaf_49_clk _00931_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dfxtp_1
X_12553_ cpuregs\[20\]\[22\] cpuregs\[21\]\[22\] _05979_ VGND VGND VPWR VPWR _06301_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11504_ decoded_imm_j\[13\] _05217_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__nand2_1
X_15272_ clknet_leaf_107_clk _00865_ VGND VGND VPWR VPWR decoded_imm_j\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12484_ _06142_ _06234_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14223_ cpuregs\[8\]\[24\] _06975_ _01732_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_544 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11435_ _05327_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14154_ _01700_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__clkbuf_1
X_11366_ _05187_ _05265_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13105_ net166 net128 _06685_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__mux2_1
X_10317_ net713 _03386_ _04599_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__mux2_1
X_14085_ net999 _06973_ _01660_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__mux2_1
X_11297_ _05194_ net1221 _01843_ _05216_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13036_ _06655_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__clkbuf_1
X_10248_ _04597_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10179_ net1047 _03386_ _04525_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__mux2_1
X_14987_ clknet_leaf_83_clk _00645_ VGND VGND VPWR VPWR reg_next_pc\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13938_ net1338 _06962_ _01577_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13869_ cpuregs\[22\]\[18\] _06962_ _07111_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15608_ clknet_leaf_122_clk _01183_ VGND VGND VPWR VPWR cpuregs\[31\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_07390_ _02019_ _02022_ _02036_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15539_ clknet_leaf_22_clk _01124_ VGND VGND VPWR VPWR cpuregs\[24\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09060_ _02030_ _03480_ _03074_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__a21o_1
X_08011_ _02624_ _02625_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold602 cpuregs\[18\]\[5\] VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold613 cpuregs\[27\]\[1\] VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 cpuregs\[26\]\[22\] VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold635 _05037_ VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 cpuregs\[1\]\[23\] VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 cpuregs\[19\]\[14\] VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 reg_next_pc\[4\] VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 cpuregs\[17\]\[28\] VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ _03415_ _04408_ _03420_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__o21a_1
X_08913_ _01862_ _01869_ _01898_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__o21ai_2
X_09893_ _01958_ _04334_ _04336_ _03651_ _04341_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__clkbuf_4
X_08775_ net1335 _03268_ _03249_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__mux2_1
X_07726_ _02327_ _02335_ _02336_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07657_ reg_pc\[23\] decoded_imm\[23\] VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_839 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07588_ net180 VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__buf_4
XFILLER_0_63_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09327_ _02082_ _03624_ _03793_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_552 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09258_ cpuregs\[4\]\[6\] cpuregs\[5\]\[6\] cpuregs\[6\]\[6\] cpuregs\[7\]\[6\] _03719_
+ _03450_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08209_ _02801_ _02808_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__nand2_1
X_09189_ net243 VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11220_ count_instr\[53\] count_instr\[52\] count_instr\[51\] _05156_ VGND VGND VPWR
+ VPWR _05162_ sky130_fd_sc_hd__and4_4
XFILLER_0_114_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11151_ count_instr\[31\] net377 count_instr\[32\] VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__a21o_1
X_10102_ net1033 _03367_ _04509_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__mux2_1
X_11082_ net679 _05063_ _05044_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_8_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910_ clknet_leaf_123_clk _00568_ VGND VGND VPWR VPWR count_instr\[19\] sky130_fd_sc_hd__dfxtp_1
X_10033_ _03474_ _04469_ _04477_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__and3_1
X_15890_ clknet_leaf_4_clk _01462_ VGND VGND VPWR VPWR cpuregs\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_14841_ clknet_leaf_1_clk _00499_ VGND VGND VPWR VPWR cpuregs\[20\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_14772_ clknet_leaf_158_clk _00430_ VGND VGND VPWR VPWR cpuregs\[16\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11984_ _05778_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__clkbuf_1
X_13723_ net809 _06952_ _07039_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10935_ net1143 _04854_ _04970_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_828 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13654_ _07006_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__clkbuf_1
X_10866_ _04941_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12605_ _06348_ _06349_ _03082_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__mux2_2
X_13585_ _06963_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__clkbuf_1
X_10797_ net1378 _04852_ _04898_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15324_ clknet_leaf_135_clk _00914_ VGND VGND VPWR VPWR cpuregs\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12536_ cpuregs\[4\]\[22\] cpuregs\[5\]\[22\] _03051_ VGND VGND VPWR VPWR _06284_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15255_ clknet_leaf_79_clk _00848_ VGND VGND VPWR VPWR instr_srai sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12467_ cpuregs\[22\]\[18\] cpuregs\[23\]\[18\] _05816_ VGND VGND VPWR VPWR _06219_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14206_ net650 _06958_ _01721_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11418_ decoded_imm_j\[6\] _05201_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15186_ clknet_leaf_72_clk _00811_ VGND VGND VPWR VPWR latched_is_lb sky130_fd_sc_hd__dfxtp_1
X_12398_ _01918_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_93_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14137_ _01691_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11349_ reg_next_pc\[28\] _03362_ _02948_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__mux2_2
X_14068_ net1085 _06956_ _01649_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__mux2_1
X_13019_ _06646_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__clkbuf_1
X_08560_ reg_sh\[3\] net1405 _01915_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_124_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07511_ reg_pc\[13\] decoded_imm\[13\] VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08491_ _03020_ _01861_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__nor2_8
XFILLER_0_71_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07442_ _02083_ _02084_ _02085_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07373_ _01951_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09112_ cpuregs\[8\]\[3\] cpuregs\[9\]\[3\] cpuregs\[10\]\[3\] cpuregs\[11\]\[3\]
+ _03582_ _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_40_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_820 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09043_ cpuregs\[12\]\[1\] cpuregs\[13\]\[1\] _03516_ VGND VGND VPWR VPWR _03517_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold410 cpuregs\[18\]\[0\] VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 cpuregs\[16\]\[4\] VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 cpuregs\[10\]\[19\] VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 cpuregs\[25\]\[25\] VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 reg_next_pc\[26\] VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold465 count_cycle\[60\] VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 cpuregs\[9\]\[9\] VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 cpuregs\[24\]\[28\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold498 cpuregs\[13\]\[13\] VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09945_ net252 _03390_ _03660_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_55_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _03472_ _04316_ _04325_ _03525_ reg_pc\[25\] VGND VGND VPWR VPWR _04326_
+ sky130_fd_sc_hd__a32o_1
X_08827_ _03313_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__clkbuf_4
X_08758_ _03173_ _03251_ _03252_ _03253_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__a22o_4
X_07709_ _02018_ _02324_ _02334_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08689_ _03193_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__buf_2
X_10720_ _04857_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_138_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10651_ net1137 _03360_ _04804_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10582_ _04775_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__clkbuf_1
X_13370_ net850 _04865_ _06838_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12321_ _02463_ _06078_ _06052_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15040_ clknet_leaf_122_clk _00698_ VGND VGND VPWR VPWR count_cycle\[23\] sky130_fd_sc_hd__dfxtp_1
X_12252_ cpuregs\[4\]\[10\] cpuregs\[5\]\[10\] cpuregs\[6\]\[10\] cpuregs\[7\]\[10\]
+ _06011_ _03097_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_75_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_536 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11203_ count_instr\[48\] _05148_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__or2_1
X_12183_ cpuregs\[20\]\[7\] cpuregs\[21\]\[7\] cpuregs\[22\]\[7\] cpuregs\[23\]\[7\]
+ _05921_ _05922_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__mux4_1
X_11134_ _05102_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__clkbuf_1
X_11065_ count_instr\[6\] _05051_ _05044_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__o21ai_1
X_15942_ clknet_leaf_26_clk _01514_ VGND VGND VPWR VPWR cpuregs\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_10016_ _03397_ _04456_ _04457_ _04460_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__a31o_1
X_15873_ clknet_leaf_22_clk _01445_ VGND VGND VPWR VPWR cpuregs\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_14824_ clknet_leaf_23_clk _00482_ VGND VGND VPWR VPWR cpuregs\[25\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ clknet_leaf_125_clk _00413_ VGND VGND VPWR VPWR cpuregs\[26\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11967_ _05769_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13706_ net1184 _06935_ _07028_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_258 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10918_ net1318 _04837_ _04959_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14686_ clknet_leaf_147_clk _00344_ VGND VGND VPWR VPWR cpuregs\[27\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11898_ count_cycle\[53\] count_cycle\[54\] VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13637_ _06997_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10849_ _04932_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13568_ _03267_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__buf_2
XFILLER_0_109_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15307_ clknet_leaf_8_clk _00897_ VGND VGND VPWR VPWR cpuregs\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12519_ _06058_ _06267_ _06182_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13499_ net1323 _04858_ _06899_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15238_ clknet_leaf_76_clk _00831_ VGND VGND VPWR VPWR instr_sltiu sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_50_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15169_ clknet_leaf_51_clk _00794_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_22_394 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07991_ _02515_ _02600_ _02607_ _02585_ VGND VGND VPWR VPWR alu_out\[3\] sky130_fd_sc_hd__a22o_1
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ cpuregs\[4\]\[21\] cpuregs\[5\]\[21\] cpuregs\[6\]\[21\] cpuregs\[7\]\[21\]
+ _03800_ _03801_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__mux4_1
X_09661_ decoded_imm\[18\] _02222_ _04089_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__a21oi_1
X_08612_ cpuregs\[0\]\[4\] cpuregs\[1\]\[4\] cpuregs\[2\]\[4\] cpuregs\[3\]\[4\] _03107_
+ _03129_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09592_ _02200_ _03486_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08543_ _03039_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08474_ reg_next_pc\[28\] reg_out\[28\] _02991_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07425_ _02065_ _02066_ _02069_ _01927_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07356_ _02002_ _02003_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07287_ mem_wordsize\[2\] _01880_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_154_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09026_ _03413_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__buf_6
XFILLER_0_5_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold240 cpuregs\[7\]\[15\] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 cpuregs\[0\]\[6\] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 cpuregs\[5\]\[12\] VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold273 cpuregs\[0\]\[11\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 cpuregs\[23\]\[2\] VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 cpuregs\[0\]\[20\] VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09928_ cpuregs\[24\]\[27\] cpuregs\[25\]\[27\] cpuregs\[26\]\[27\] cpuregs\[27\]\[27\]
+ _03594_ _03442_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_70_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09859_ cpuregs\[4\]\[25\] cpuregs\[5\]\[25\] cpuregs\[6\]\[25\] cpuregs\[7\]\[25\]
+ _03800_ _03407_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_29_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ mem_rdata_q\[31\] mem_rdata_q\[29\] _06563_ mem_rdata_q\[30\] VGND VGND VPWR
+ VPWR _06566_ sky130_fd_sc_hd__nor4b_4
XFILLER_0_99_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_102 _06888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11821_ _05660_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__clkbuf_1
*XANTENNA_113 mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_124 net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_135 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_146 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_157 _03095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14540_ clknet_leaf_26_clk _00198_ VGND VGND VPWR VPWR cpuregs\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11752_ _05611_ _05612_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__nor2_1
*XANTENNA_168 _03474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_179 _04846_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10703_ _03267_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_101_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ clknet_leaf_98_clk _00129_ VGND VGND VPWR VPWR cpuregs\[12\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _05273_ _05541_ _05251_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_154_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13422_ _06868_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10634_ net1135 _03307_ _04793_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_64_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13353_ net1016 _04848_ _06827_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__mux2_1
X_10565_ _04766_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__clkbuf_1
X_12304_ cpuregs\[8\]\[12\] cpuregs\[9\]\[12\] cpuregs\[10\]\[12\] cpuregs\[11\]\[12\]
+ _06061_ _05917_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13284_ _06795_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__clkbuf_1
X_10496_ _04729_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15023_ clknet_leaf_111_clk _00681_ VGND VGND VPWR VPWR count_cycle\[6\] sky130_fd_sc_hd__dfxtp_1
X_12235_ _05912_ _05995_ _03123_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_887 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12166_ cpuregs\[28\]\[6\] cpuregs\[29\]\[6\] cpuregs\[30\]\[6\] cpuregs\[31\]\[6\]
+ _05895_ _05929_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__mux4_1
X_11117_ net1172 _05087_ _05090_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__o21ai_1
X_12097_ decoded_imm\[2\] _03071_ _01906_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__mux2_1
X_15925_ clknet_leaf_16_clk _01497_ VGND VGND VPWR VPWR cpuregs\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11048_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__buf_4
Xinput8 net421 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_88_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15856_ clknet_leaf_16_clk _01428_ VGND VGND VPWR VPWR cpuregs\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807_ clknet_leaf_153_clk _00465_ VGND VGND VPWR VPWR cpuregs\[25\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15787_ clknet_leaf_4_clk _01362_ VGND VGND VPWR VPWR cpuregs\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12999_ _06635_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_158_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14738_ clknet_leaf_55_clk _00396_ VGND VGND VPWR VPWR cpuregs\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_129_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14669_ clknet_leaf_37_clk _00327_ VGND VGND VPWR VPWR cpuregs\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07210_ instr_sw instr_sh instr_sb _01874_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__or4b_1
XFILLER_0_116_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08190_ net212 net211 net247 _02759_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__or4_1
XFILLER_0_144_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_100_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07974_ _02590_ _02591_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__xor2_1
X_09713_ cpuregs\[8\]\[20\] cpuregs\[9\]\[20\] cpuregs\[10\]\[20\] cpuregs\[11\]\[20\]
+ _03601_ _03583_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__mux4_1
X_09644_ _03454_ _04100_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__or2_1
X_09575_ cpuregs\[20\]\[16\] cpuregs\[21\]\[16\] cpuregs\[22\]\[16\] cpuregs\[23\]\[16\]
+ _03673_ _03674_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08526_ _00007_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_67_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08457_ reg_next_pc\[23\] reg_out\[23\] _02991_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07408_ count_instr\[39\] _02052_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__and2_1
X_08388_ _02948_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__buf_4
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07339_ _01971_ decoded_imm\[2\] VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_150_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10350_ net656 _03275_ _04647_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_104_878 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09009_ _01846_ _02008_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__mux2_1
X_10281_ _04615_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ net54 net85 _05766_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__mux2_1
X_13971_ cpuregs\[5\]\[1\] _06927_ _01602_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__mux2_1
X_15710_ clknet_leaf_20_clk _01285_ VGND VGND VPWR VPWR cpuregs\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_607 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12922_ mem_rdata_q\[28\] net21 _06589_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__mux2_1
X_15641_ clknet_leaf_153_clk _01216_ VGND VGND VPWR VPWR cpuregs\[23\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ _06558_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_85_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11804_ count_cycle\[22\] count_cycle\[23\] count_cycle\[24\] _05640_ VGND VGND VPWR
+ VPWR _05649_ sky130_fd_sc_hd__and4_4
X_15572_ clknet_leaf_133_clk _01147_ VGND VGND VPWR VPWR cpuregs\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12784_ _06515_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_83_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ clknet_leaf_10_clk _00181_ VGND VGND VPWR VPWR cpuregs\[13\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_11735_ count_cycle\[0\] count_cycle\[1\] count_cycle\[2\] count_cycle\[3\] VGND
+ VGND VPWR VPWR _05601_ sky130_fd_sc_hd__and4_4
XFILLER_0_127_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14454_ clknet_leaf_13_clk _00112_ VGND VGND VPWR VPWR cpuregs\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11666_ _05288_ _05540_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_935 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _06859_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__clkbuf_1
X_10617_ _04794_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__clkbuf_1
X_14385_ clknet_leaf_8_clk _00048_ VGND VGND VPWR VPWR cpuregs\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11597_ _05470_ _05472_ _05477_ _05367_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13336_ cpuregs\[19\]\[6\] _04831_ _06816_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__mux2_1
X_10548_ net1148 _03248_ _04757_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_94_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13267_ _06786_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__clkbuf_1
X_10479_ cpuregs\[14\]\[10\] _03248_ _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15006_ clknet_leaf_109_clk _00664_ VGND VGND VPWR VPWR reg_next_pc\[21\] sky130_fd_sc_hd__dfxtp_1
X_12218_ cpuregs\[20\]\[8\] cpuregs\[21\]\[8\] _05979_ VGND VGND VPWR VPWR _05980_
+ sky130_fd_sc_hd__mux2_1
X_13198_ decoded_imm\[25\] _06740_ _06737_ _06747_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__o22a_1
X_12149_ _03062_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15908_ clknet_leaf_26_clk _01480_ VGND VGND VPWR VPWR cpuregs\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_07690_ net18 _02252_ _02180_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__a21o_1
X_15839_ clknet_leaf_132_clk _01411_ VGND VGND VPWR VPWR cpuregs\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09360_ _02154_ _03480_ _03709_ _03074_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08311_ _02369_ _02901_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_857 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09291_ _03436_ _03758_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_138_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
*XANTENNA_13 _01978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08242_ _02831_ _02833_ _02829_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_24 _03143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_35 _03230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_46 _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_57 _03489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_68 _03588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08173_ _02762_ _02766_ _02774_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__a21o_1
*XANTENNA_79 _04818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_104_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput120 net120 VGND VGND VPWR VPWR mem_la_wdata[30] sky130_fd_sc_hd__clkbuf_4
Xoutput131 net131 VGND VGND VPWR VPWR mem_la_wstrb[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput142 net142 VGND VGND VPWR VPWR mem_wdata[16] sky130_fd_sc_hd__clkbuf_4
Xoutput153 net153 VGND VGND VPWR VPWR mem_wdata[26] sky130_fd_sc_hd__clkbuf_4
Xoutput164 net164 VGND VGND VPWR VPWR mem_wdata[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput175 net175 VGND VGND VPWR VPWR pcpi_rs1[13] sky130_fd_sc_hd__clkbuf_4
Xoutput186 net186 VGND VGND VPWR VPWR pcpi_rs1[23] sky130_fd_sc_hd__clkbuf_4
Xoutput197 net197 VGND VGND VPWR VPWR pcpi_rs1[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_149_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07957_ _02574_ _02575_ net182 VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07888_ _01931_ _02507_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__or2_1
X_09627_ decoded_imm\[18\] net180 VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__nand2_1
X_09558_ _04017_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08509_ decoded_imm_j\[19\] _01081_ _03022_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09489_ _03475_ _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_654 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_148_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11520_ decoded_imm_j\[14\] _05219_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_827 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11451_ _01842_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10402_ net851 _03221_ _04673_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__mux2_1
X_14170_ _01708_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__clkbuf_1
X_11382_ decoded_imm_j\[2\] _05191_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13121_ _06703_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10333_ net886 _03221_ _04636_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__mux2_1
X_13052_ cpuregs\[1\]\[25\] _04871_ _06658_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10264_ _04606_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__clkbuf_1
X_12003_ _05788_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__clkbuf_1
X_10195_ net830 _03215_ _04564_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__mux2_1
X_13954_ _01594_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__clkbuf_1
X_12905_ _02013_ _06553_ _06582_ net239 VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__a22o_1
X_13885_ _01557_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ clknet_leaf_30_clk _01199_ VGND VGND VPWR VPWR cpuregs\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12836_ _06532_ net6 _03017_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_8_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15555_ clknet_leaf_44_clk _01130_ VGND VGND VPWR VPWR cpuregs\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12767_ _01945_ _02558_ _06504_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14506_ clknet_leaf_54_clk _00164_ VGND VGND VPWR VPWR cpuregs\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11718_ _05263_ net539 _05358_ _05588_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__o211a_1
X_15486_ clknet_leaf_92_clk _01071_ VGND VGND VPWR VPWR mem_rdata_q\[9\] sky130_fd_sc_hd__dfxtp_1
X_12698_ cpuregs\[0\]\[29\] cpuregs\[1\]\[29\] cpuregs\[2\]\[29\] cpuregs\[3\]\[29\]
+ _03091_ _05829_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_553 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_65_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14437_ clknet_leaf_96_clk _00095_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dfxtp_4
X_11649_ _05289_ _05520_ _05521_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__a31o_1
Xinput11 net419 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_116_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput22 net413 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput33 mem_ready VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14368_ _01811_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_491 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_40_724 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold806 cpuregs\[28\]\[17\] VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 cpuregs\[9\]\[16\] VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold828 cpuregs\[8\]\[19\] VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ _06813_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold839 cpuregs\[18\]\[7\] VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__dlygate4sd3_1
X_14299_ net560 VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08860_ _03342_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__clkbuf_1
X_07811_ net187 net246 VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__nand2_1
X_08791_ net582 _03282_ _03249_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__mux2_1
X_07742_ reg_pc\[29\] decoded_imm\[29\] VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__nand2_1
X_07673_ reg_pc\[24\] decoded_imm\[24\] VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_144_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09412_ _03427_ _03871_ _03873_ _03875_ _03490_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_36_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09343_ cpuregs\[12\]\[9\] cpuregs\[13\]\[9\] cpuregs\[14\]\[9\] cpuregs\[15\]\[9\]
+ _03808_ _03801_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09274_ _03482_ _03741_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08225_ _02265_ net216 _02822_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__o22a_1
XFILLER_0_160_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_586 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08156_ _02757_ _02759_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08087_ _02694_ _02695_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08989_ _03459_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10951_ _04986_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13670_ net1259 _06966_ _07014_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__mux2_1
X_10882_ net827 _04869_ _04945_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12621_ net220 _06365_ _06282_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_159_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15340_ clknet_leaf_49_clk _00930_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dfxtp_2
X_12552_ _06297_ _06298_ _06299_ _05873_ _03113_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11503_ decoded_imm_j\[13\] _05217_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15271_ clknet_leaf_105_clk _00864_ VGND VGND VPWR VPWR decoded_imm_j\[19\] sky130_fd_sc_hd__dfxtp_1
X_12483_ cpuregs\[20\]\[19\] cpuregs\[21\]\[19\] cpuregs\[22\]\[19\] cpuregs\[23\]\[19\]
+ _06065_ _03144_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14222_ _01736_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11434_ _05204_ _05312_ _01903_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14153_ net1023 _06973_ _01696_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_100_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_100_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_78_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11365_ decoded_imm_j\[1\] _05264_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__nand2_1
X_13104_ _06694_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__clkbuf_1
X_10316_ _04633_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14084_ _01663_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__clkbuf_1
X_11296_ _05031_ _05215_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__nand2_1
X_13035_ net1053 _04854_ _06647_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__mux2_1
X_10247_ net665 _03381_ _04563_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10178_ _04559_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14986_ clknet_leaf_82_clk _00644_ VGND VGND VPWR VPWR reg_next_pc\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13937_ _01585_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13868_ _01548_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15607_ clknet_leaf_129_clk _01182_ VGND VGND VPWR VPWR cpuregs\[31\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12819_ _01901_ decoder_pseudo_trigger VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__or2_4
XFILLER_0_9_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13799_ net1205 _06960_ _07075_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__mux2_1
X_15538_ clknet_leaf_125_clk _01123_ VGND VGND VPWR VPWR cpuregs\[24\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_151_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_564 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15469_ clknet_leaf_125_clk _01059_ VGND VGND VPWR VPWR cpuregs\[19\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08010_ _02030_ _02623_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__or2_1
Xhold603 cpuregs\[3\]\[8\] VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold614 cpuregs\[21\]\[26\] VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_111_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold625 cpuregs\[11\]\[18\] VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold636 _05042_ VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold647 cpuregs\[1\]\[14\] VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_50 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold658 cpuregs\[12\]\[6\] VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ cpuregs\[8\]\[28\] cpuregs\[9\]\[28\] cpuregs\[10\]\[28\] cpuregs\[11\]\[28\]
+ _03641_ _03642_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold669 cpuregs\[30\]\[9\] VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__dlygate4sd3_1
X_08912_ _03387_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09892_ _04337_ _04340_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08843_ _03324_ _03327_ _03293_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_146_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08774_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__clkbuf_4
X_07725_ count_cycle\[28\] _02020_ _02347_ _02348_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_158_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_158_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07656_ reg_pc\[23\] decoded_imm\[23\] VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07587_ _02219_ _02220_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09326_ _03672_ _03769_ _03774_ _03792_ _03665_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__o311a_1
XFILLER_0_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_118_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09257_ _03436_ _03725_ _03467_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08208_ _02756_ net237 _02807_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_178 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09188_ instr_srl instr_srli _03390_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__nor3_1
X_08139_ net177 _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11150_ _01839_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__clkbuf_4
X_10101_ _04517_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_464 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11081_ count_instr\[11\] count_instr\[10\] _05062_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ _04471_ _04473_ _04476_ _03427_ _03490_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__a221o_1
X_14840_ clknet_leaf_153_clk _00498_ VGND VGND VPWR VPWR cpuregs\[20\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_14771_ clknet_leaf_29_clk _00429_ VGND VGND VPWR VPWR cpuregs\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_149_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_149_clk sky130_fd_sc_hd__clkbuf_2
X_11983_ net36 net67 _05774_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__mux2_1
X_13722_ _07042_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__clkbuf_1
X_10934_ _04977_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_85_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13653_ cpuregs\[23\]\[12\] _06950_ _07003_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10865_ net646 _04852_ _04934_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12604_ cpuregs\[0\]\[25\] cpuregs\[1\]\[25\] cpuregs\[2\]\[25\] cpuregs\[3\]\[25\]
+ _06055_ _05829_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_94_771 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13584_ net1186 _06962_ _06946_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__mux2_1
X_10796_ _04904_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15323_ clknet_leaf_20_clk _00913_ VGND VGND VPWR VPWR cpuregs\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12535_ _06283_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15254_ clknet_leaf_76_clk _00847_ VGND VGND VPWR VPWR instr_and sky130_fd_sc_hd__dfxtp_1
X_12466_ _05872_ _06217_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14205_ _01727_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__clkbuf_1
X_11417_ _05199_ _05201_ _05296_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15185_ clknet_leaf_72_clk _00810_ VGND VGND VPWR VPWR latched_is_lh sky130_fd_sc_hd__dfxtp_1
X_12397_ _06144_ _06146_ _06148_ _06150_ _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__a221o_2
XFILLER_0_2_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14136_ net599 _06956_ _01685_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__mux2_1
X_11348_ _05227_ _05251_ _05252_ _05224_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14067_ _01654_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__clkbuf_1
X_11279_ reg_next_pc\[7\] _02999_ _05203_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__a21o_2
X_13018_ net929 _04837_ _06636_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__mux2_1
X_14969_ clknet_leaf_105_clk _00627_ VGND VGND VPWR VPWR reg_pc\[15\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_124_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07510_ reg_pc\[13\] decoded_imm\[13\] VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_141_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08490_ mem_do_rinst VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07441_ latched_is_lb _02069_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__and2_2
XFILLER_0_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07372_ _02018_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09111_ _03408_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_40_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09042_ _03404_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__buf_8
XFILLER_0_5_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_41_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold400 cpuregs\[17\]\[31\] VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold411 cpuregs\[7\]\[3\] VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 decoded_imm\[31\] VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 cpuregs\[1\]\[3\] VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 cpuregs\[20\]\[28\] VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold455 cpuregs\[27\]\[29\] VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 cpuregs\[11\]\[9\] VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 cpuregs\[14\]\[26\] VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold488 cpuregs\[15\]\[29\] VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ _04391_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__clkbuf_1
Xhold499 cpuregs\[15\]\[9\] VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _04318_ _04320_ _04322_ _04324_ _03429_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_5_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _03309_ _03312_ _03293_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__mux2_2
X_08757_ reg_pc\[11\] _03245_ _03172_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__a21oi_1
X_07708_ _02058_ _02330_ _02333_ _01968_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_727 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08688_ _03191_ _03192_ _03172_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__mux2_2
X_07639_ reg_pc\[22\] decoded_imm\[22\] VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10650_ _04811_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09309_ _03403_ _03775_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_350 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10581_ net741 _03355_ _04768_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__mux2_1
X_12320_ _05901_ _06064_ _06077_ _05904_ decoded_imm\[12\] VGND VGND VPWR VPWR _06078_
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12251_ _05907_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_375 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11202_ _05148_ _05149_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_548 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12182_ _05879_ _05940_ _05942_ _05944_ _03104_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__a221o_2
X_11133_ _05100_ _01884_ _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__and3b_1
X_11064_ count_instr\[6\] _05051_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__and2_1
X_15941_ clknet_leaf_37_clk _01513_ VGND VGND VPWR VPWR cpuregs\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_10015_ _01943_ _04458_ _04459_ _03476_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__a31o_1
X_15872_ clknet_leaf_22_clk _01444_ VGND VGND VPWR VPWR cpuregs\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_14823_ clknet_leaf_127_clk _00481_ VGND VGND VPWR VPWR cpuregs\[25\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14754_ clknet_leaf_126_clk _00412_ VGND VGND VPWR VPWR cpuregs\[26\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11966_ net812 net89 _05767_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_401 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10917_ _04968_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__clkbuf_1
X_13705_ _07033_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__clkbuf_1
X_14685_ clknet_leaf_156_clk _00343_ VGND VGND VPWR VPWR cpuregs\[27\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_626 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11897_ net454 VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_719 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_132_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_445 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13636_ net1244 _06933_ _06992_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__mux2_1
X_10848_ net1119 _04835_ _04923_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13567_ _06951_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10779_ _04895_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15306_ clknet_leaf_11_clk _00896_ VGND VGND VPWR VPWR cpuregs\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_12518_ cpuregs\[12\]\[21\] cpuregs\[13\]\[21\] cpuregs\[14\]\[21\] cpuregs\[15\]\[21\]
+ _03133_ _05994_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__mux4_1
X_13498_ _06908_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12449_ _05871_ _06200_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__and2_1
X_15237_ clknet_leaf_77_clk _00830_ VGND VGND VPWR VPWR instr_slti sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15168_ clknet_leaf_51_clk _00793_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14119_ net1345 _06939_ _01674_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__mux2_1
X_15099_ clknet_leaf_100_clk _07122_ VGND VGND VPWR VPWR reg_out\[17\] sky130_fd_sc_hd__dfxtp_1
X_07990_ _02605_ _02606_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_54 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09660_ _04114_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_105_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08611_ _03047_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__clkbuf_8
X_09591_ reg_pc\[16\] _03528_ _04049_ _03626_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__a211o_1
X_08542_ _03038_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__buf_6
XFILLER_0_82_64 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_159_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08473_ _03008_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
XFILLER_0_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_423 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_148_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07424_ net30 net130 _02068_ _01940_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_123 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_46_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_114_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07355_ reg_pc\[4\] decoded_imm\[4\] VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07286_ _01935_ _01936_ _01937_ net8 VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_154_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ _03497_ _03498_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_57_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold230 cpuregs\[10\]\[15\] VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 reg_next_pc\[22\] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 cpuregs\[0\]\[14\] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 cpuregs\[28\]\[25\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 cpuregs\[5\]\[4\] VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 cpuregs\[3\]\[5\] VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 cpuregs\[17\]\[1\] VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ _03402_ _04374_ _03603_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_70_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_123_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09858_ _04304_ _04305_ _04306_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08809_ reg_pc\[18\] _03291_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _04239_ _04240_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_29_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _05658_ _05625_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__and3b_1
XFILLER_0_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_103 _07028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_114 reg_next_pc\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_125 net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_136 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_147 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11751_ net623 _05609_ _05169_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__o21ai_1
*XANTENNA_158 _03173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_169 _03547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_80_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_2
X_10702_ _04845_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__clkbuf_1
X_14470_ clknet_leaf_97_clk _00128_ VGND VGND VPWR VPWR cpuregs\[12\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11682_ _05551_ _05555_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_101_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_132_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13421_ net1314 _04848_ _06863_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__mux2_1
X_10633_ _04802_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13352_ _06831_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__clkbuf_1
X_10564_ net1330 _03302_ _04757_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_651 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_51_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12303_ _03046_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__clkbuf_8
X_13283_ net1181 _04846_ _06791_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10495_ net808 _03302_ _04720_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15022_ clknet_leaf_111_clk _00680_ VGND VGND VPWR VPWR count_cycle\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12234_ cpuregs\[12\]\[9\] cpuregs\[13\]\[9\] cpuregs\[14\]\[9\] cpuregs\[15\]\[9\]
+ _05913_ _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12165_ _03063_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__buf_4
XFILLER_0_130_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_899 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11116_ _05040_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__clkbuf_4
X_12096_ _05864_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15924_ clknet_leaf_143_clk _01496_ VGND VGND VPWR VPWR cpuregs\[0\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11047_ _01839_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__buf_4
XFILLER_0_36_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 net409 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_88_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ clknet_leaf_16_clk _01427_ VGND VGND VPWR VPWR cpuregs\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_88_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14806_ clknet_leaf_156_clk _00464_ VGND VGND VPWR VPWR cpuregs\[25\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ clknet_leaf_7_clk _01361_ VGND VGND VPWR VPWR cpuregs\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12998_ _04483_ _04562_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__nor2_2
XFILLER_0_148_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14737_ clknet_leaf_36_clk _00395_ VGND VGND VPWR VPWR cpuregs\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11949_ _04453_ _04457_ _05753_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_71_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_143_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14668_ clknet_leaf_27_clk _00326_ VGND VGND VPWR VPWR cpuregs\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_404 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13619_ _06986_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14599_ clknet_leaf_131_clk _00257_ VGND VGND VPWR VPWR cpuregs\[28\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07973_ _02566_ _02577_ _02576_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_52_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09712_ _03454_ _04166_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__or2_1
X_09643_ cpuregs\[28\]\[18\] cpuregs\[29\]\[18\] cpuregs\[30\]\[18\] cpuregs\[31\]\[18\]
+ _03598_ _03716_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__mux4_1
X_09574_ cpuregs\[16\]\[16\] cpuregs\[17\]\[16\] cpuregs\[18\]\[16\] cpuregs\[19\]\[16\]
+ _03673_ _03674_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__mux4_1
X_08525_ _00009_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08456_ _02996_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07407_ _01946_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__buf_2
X_08387_ _02947_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07338_ reg_pc\[3\] decoded_imm\[3\] VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07269_ _01907_ _01923_ _01916_ _01838_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__and4b_1
X_09008_ _03482_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10280_ net938 _03268_ _04611_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13970_ _01603_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__clkbuf_1
X_12921_ _06595_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_619 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_87_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15640_ clknet_leaf_122_clk _01215_ VGND VGND VPWR VPWR cpuregs\[23\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12852_ is_alu_reg_imm _06528_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__and2_1
X_11803_ _05646_ _05648_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_140_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15571_ clknet_leaf_140_clk _01146_ VGND VGND VPWR VPWR cpuregs\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12783_ mem_rdata_q\[2\] net23 _03017_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_83_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _05600_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__clkbuf_1
X_14522_ clknet_leaf_10_clk _00180_ VGND VGND VPWR VPWR cpuregs\[13\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_83_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11665_ _05249_ _05528_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__nor2_1
X_14453_ clknet_leaf_31_clk _00111_ VGND VGND VPWR VPWR cpuregs\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10616_ cpuregs\[15\]\[10\] _03248_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__mux2_1
X_13404_ cpuregs\[24\]\[6\] _04831_ _06852_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ clknet_leaf_11_clk _00047_ VGND VGND VPWR VPWR cpuregs\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11596_ _05475_ _05476_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_446 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_106_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13335_ _06822_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__clkbuf_1
X_10547_ _04745_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__buf_4
XFILLER_0_106_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13266_ net961 _04829_ _06780_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__mux2_1
X_10478_ _04708_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_114_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15005_ clknet_leaf_106_clk _00663_ VGND VGND VPWR VPWR reg_next_pc\[20\] sky130_fd_sc_hd__dfxtp_1
X_12217_ _03038_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__buf_4
X_13197_ mem_rdata_q\[25\] _06742_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12148_ _03082_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12079_ cpuregs\[0\]\[1\] cpuregs\[1\]\[1\] cpuregs\[2\]\[1\] cpuregs\[3\]\[1\] _03091_
+ _03125_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__mux4_1
X_15907_ clknet_leaf_50_clk _01479_ VGND VGND VPWR VPWR cpuregs\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15838_ clknet_leaf_129_clk _01410_ VGND VGND VPWR VPWR cpuregs\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15769_ clknet_leaf_141_clk _01344_ VGND VGND VPWR VPWR cpuregs\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_44_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08310_ net224 _02900_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09290_ cpuregs\[24\]\[7\] cpuregs\[25\]\[7\] cpuregs\[26\]\[7\] cpuregs\[27\]\[7\]
+ _03463_ _03464_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08241_ net186 _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__xnor2_2
*XANTENNA_14 _02057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_25 _03143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_700 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_16_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_36 _03248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_47 _03329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
*XANTENNA_58 _03492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ _02762_ _02766_ _02774_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__nand3_1
XFILLER_0_133_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_69 _03588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_552 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_125_470 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput110 net110 VGND VGND VPWR VPWR mem_la_wdata[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput121 net121 VGND VGND VPWR VPWR mem_la_wdata[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput132 net132 VGND VGND VPWR VPWR mem_la_wstrb[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput143 net143 VGND VGND VPWR VPWR mem_wdata[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput154 net154 VGND VGND VPWR VPWR mem_wdata[27] sky130_fd_sc_hd__clkbuf_4
Xoutput165 net165 VGND VGND VPWR VPWR mem_wdata[8] sky130_fd_sc_hd__clkbuf_4
Xoutput176 net176 VGND VGND VPWR VPWR pcpi_rs1[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput187 net187 VGND VGND VPWR VPWR pcpi_rs1[24] sky130_fd_sc_hd__clkbuf_4
Xoutput198 net198 VGND VGND VPWR VPWR pcpi_rs1[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_149_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07956_ _02572_ net97 net108 VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__and3_1
X_07887_ net97 VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09626_ decoded_imm\[18\] net180 VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__or2_1
X_09557_ _02177_ _04016_ _03395_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_65_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08508_ _03030_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__buf_1
X_09488_ _03472_ _03940_ _03949_ _03526_ reg_pc\[13\] VGND VGND VPWR VPWR _03950_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08439_ _02984_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_1
XFILLER_0_93_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11450_ _05258_ net523 _05239_ _05342_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__o211a_1
Xwire237 _02803_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_1
X_10401_ _04679_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__clkbuf_1
X_11381_ decoded_imm_j\[2\] _05191_ _05275_ _05278_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13120_ net1154 net104 _06696_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10332_ _04642_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_298 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13051_ _06663_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_484 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10263_ net596 _03215_ _04600_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__mux2_1
X_12002_ net512 net76 _05785_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__mux2_1
X_10194_ _04569_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_89_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13953_ cpuregs\[4\]\[25\] _06977_ _01588_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__mux2_1
X_12904_ net444 _06530_ _06535_ net241 VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13884_ net832 _06977_ _01551_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15623_ clknet_leaf_25_clk _01198_ VGND VGND VPWR VPWR cpuregs\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _06550_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__buf_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15554_ clknet_leaf_37_clk _01129_ VGND VGND VPWR VPWR cpuregs\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12766_ _01927_ _01894_ _03389_ _06503_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__or4_1
X_14505_ clknet_leaf_18_clk _00163_ VGND VGND VPWR VPWR cpuregs\[30\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_11717_ _05285_ _05260_ _05587_ _05300_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__a22o_1
X_12697_ cpuregs\[4\]\[29\] cpuregs\[5\]\[29\] cpuregs\[6\]\[29\] cpuregs\[7\]\[29\]
+ _05908_ _06156_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__mux4_1
X_15485_ clknet_leaf_92_clk _01070_ VGND VGND VPWR VPWR mem_rdata_q\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11648_ _05244_ _05522_ _05524_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__a21oi_1
X_14436_ clknet_leaf_96_clk _00094_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_154_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 net408 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_116_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput23 net986 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_116_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput34 resetn VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
X_11579_ decoded_imm_j\[19\] _05233_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__and2_1
X_14367_ net1185 _03380_ _01777_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold807 cpuregs\[30\]\[6\] VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold818 cpuregs\[22\]\[29\] VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ cpuregs\[18\]\[30\] _04881_ _06779_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__mux2_1
Xhold829 count_instr\[31\] VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ _01774_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13249_ _06763_ decoded_imm_j\[2\] _06732_ mem_rdata_q\[9\] _06540_ VGND VGND VPWR
+ VPWR _06776_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07810_ net187 net246 VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__or2_1
X_08790_ _03281_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07741_ reg_pc\[29\] decoded_imm\[29\] VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__nor2_1
X_07672_ _02247_ _02297_ _02298_ _02299_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09411_ _03647_ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_36_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_36_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09342_ _00012_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_47_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_64 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_87_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09273_ _02044_ _02082_ _03617_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_828 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08224_ _02265_ net216 _02598_ _02563_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_598 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08155_ _02657_ _02700_ _02758_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__or3_4
XFILLER_0_126_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08086_ net173 _02693_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08988_ _03456_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__buf_6
X_07939_ instr_and instr_andi VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__or2_1
X_10950_ net723 _04869_ _04981_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09609_ _03647_ _04066_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__or2_1
X_10881_ _04949_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12620_ _05900_ _06355_ _06364_ _01918_ decoded_imm\[25\] VGND VGND VPWR VPWR _06365_
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_80_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12551_ cpuregs\[28\]\[22\] cpuregs\[29\]\[22\] _03085_ VGND VGND VPWR VPWR _06299_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_666 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11502_ _05258_ reg_next_pc\[12\] _05343_ _05390_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12482_ _06177_ _06228_ _06230_ _06232_ _06164_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__a221o_1
X_15270_ clknet_leaf_86_clk _00863_ VGND VGND VPWR VPWR decoded_imm_j\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14221_ cpuregs\[8\]\[23\] _06973_ _01732_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__mux2_1
X_11433_ _05204_ _05312_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14152_ _01699_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11364_ _01889_ _01901_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__nor2_2
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10315_ net951 _03381_ _04599_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__mux2_1
X_13103_ net165 net127 _06685_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__mux2_1
X_14083_ cpuregs\[6\]\[22\] _06971_ _01660_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__mux2_1
X_11295_ reg_next_pc\[12\] _02999_ _05214_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_111_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13034_ _06654_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__clkbuf_1
X_10246_ _04596_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10177_ net785 _03381_ _04525_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__mux2_1
X_14985_ clknet_leaf_105_clk _00643_ VGND VGND VPWR VPWR reg_pc\[31\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_161_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13936_ net1042 _06960_ _01577_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13867_ cpuregs\[22\]\[17\] _06960_ _07111_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15606_ clknet_leaf_145_clk _01181_ VGND VGND VPWR VPWR cpuregs\[31\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12818_ net883 _06530_ _06539_ _05804_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13798_ _07082_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15537_ clknet_leaf_126_clk _01122_ VGND VGND VPWR VPWR cpuregs\[24\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12749_ cpuregs\[8\]\[31\] cpuregs\[9\]\[31\] cpuregs\[10\]\[31\] cpuregs\[11\]\[31\]
+ _05970_ _03137_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_115_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15468_ clknet_leaf_148_clk _01058_ VGND VGND VPWR VPWR cpuregs\[19\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_576 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_738 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14419_ clknet_leaf_62_clk _00077_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dfxtp_4
X_15399_ clknet_leaf_87_clk _00989_ VGND VGND VPWR VPWR decoded_imm\[9\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_69_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold604 cpuregs\[15\]\[0\] VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 cpuregs\[19\]\[31\] VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 cpuregs\[27\]\[13\] VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold637 cpuregs\[2\]\[6\] VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 cpuregs\[25\]\[20\] VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09960_ _04405_ _04406_ _03647_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold659 cpuregs\[29\]\[1\] VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08911_ net1057 _03386_ _03184_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09891_ _04305_ _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_31 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08842_ _03325_ _03326_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_146_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _03265_ _03266_ _03261_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__mux2_2
X_07724_ count_instr\[28\] _01965_ count_cycle\[60\] _02055_ VGND VGND VPWR VPWR _02348_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ _02055_ count_cycle\[55\] count_cycle\[23\] _02020_ _02283_ VGND VGND VPWR
+ VPWR _02284_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_791 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07586_ _02209_ _02211_ _02208_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09325_ _03474_ _03782_ _03790_ _03791_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09256_ cpuregs\[8\]\[6\] cpuregs\[9\]\[6\] cpuregs\[10\]\[6\] cpuregs\[11\]\[6\]
+ _03463_ _03464_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08207_ _02805_ _02806_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09187_ _01847_ _02082_ _03479_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08138_ net209 _02742_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08069_ net248 _02678_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__xnor2_1
X_10100_ net1196 _03360_ _04509_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__mux2_1
X_11080_ _05063_ _05064_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _04474_ _04475_ _03647_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ clknet_leaf_55_clk _00428_ VGND VGND VPWR VPWR cpuregs\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11982_ _05777_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__clkbuf_1
X_13721_ net1191 _06950_ _07039_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__mux2_1
X_10933_ net959 _04852_ _04970_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13652_ _07005_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__clkbuf_1
X_10864_ _04940_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12603_ cpuregs\[4\]\[25\] cpuregs\[5\]\[25\] cpuregs\[6\]\[25\] cpuregs\[7\]\[25\]
+ _05908_ _06156_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10795_ cpuregs\[16\]\[15\] _04850_ _04898_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__mux2_1
X_13583_ _03301_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__buf_2
XFILLER_0_155_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_783 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_176 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15322_ clknet_leaf_139_clk _00912_ VGND VGND VPWR VPWR cpuregs\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12534_ net216 _06281_ _06282_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__mux2_1
X_15253_ clknet_leaf_76_clk _00846_ VGND VGND VPWR VPWR instr_or sky130_fd_sc_hd__dfxtp_1
X_12465_ cpuregs\[20\]\[18\] cpuregs\[21\]\[18\] _05979_ VGND VGND VPWR VPWR _06217_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14204_ net1084 _06956_ _01721_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__mux2_1
X_11416_ _05258_ net571 _05239_ _05311_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12396_ _03033_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__buf_4
X_15184_ clknet_leaf_82_clk _00809_ VGND VGND VPWR VPWR decoder_pseudo_trigger sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_544 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14135_ _01690_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__clkbuf_1
X_11347_ _05231_ reg_pc\[27\] VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_18_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14066_ cpuregs\[6\]\[14\] _06954_ _01649_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__mux2_1
X_11278_ _02945_ _03226_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10229_ net1041 _03322_ _04586_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__mux2_1
X_13017_ _06645_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14968_ clknet_leaf_107_clk _00626_ VGND VGND VPWR VPWR reg_pc\[14\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_124_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13919_ net1246 _06943_ _01566_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14899_ clknet_leaf_113_clk _00557_ VGND VGND VPWR VPWR count_instr\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07440_ _01845_ _01848_ net17 net31 _01933_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07371_ _02006_ _02012_ _02016_ _02018_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__o22a_1
XFILLER_0_147_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09110_ _03554_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__buf_6
XFILLER_0_128_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09041_ cpuregs\[14\]\[1\] cpuregs\[15\]\[1\] _03406_ VGND VGND VPWR VPWR _03515_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold401 cpuregs\[25\]\[27\] VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold412 cpuregs\[27\]\[24\] VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 cpuregs\[14\]\[19\] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 cpuregs\[8\]\[25\] VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 cpuregs\[8\]\[29\] VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold456 cpuregs\[2\]\[4\] VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 cpuregs\[13\]\[9\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 cpuregs\[24\]\[27\] VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold489 cpuregs\[7\]\[16\] VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _02340_ _04390_ _03394_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _03435_ _04323_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_5_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _03310_ _03311_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__nor2_1
X_08756_ reg_pc\[11\] _03245_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__or2_1
X_07707_ _01943_ _02331_ _02184_ _02332_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08687_ reg_out\[2\] alu_out_q\[2\] latched_stalu VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_739 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_95_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07638_ _02019_ _02259_ _02268_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_569 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07569_ _02198_ _02199_ _02204_ _02071_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_24_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09308_ cpuregs\[12\]\[8\] cpuregs\[13\]\[8\] cpuregs\[14\]\[8\] cpuregs\[15\]\[8\]
+ _03494_ _03497_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__mux4_1
X_10580_ _04774_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09239_ _01978_ _02112_ _03479_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12250_ _06010_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11201_ net1241 _05146_ _05133_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_352 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12181_ _03106_ _05943_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11132_ _05095_ _05098_ count_instr\[26\] VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__a21o_1
Xhold990 cpuregs\[9\]\[25\] VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ _05049_ _05047_ _05051_ _05052_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__a211oi_1
X_15940_ clknet_leaf_26_clk _01512_ VGND VGND VPWR VPWR cpuregs\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_10014_ _02369_ _03770_ _04380_ _03616_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__a211o_1
X_15871_ clknet_leaf_132_clk _01443_ VGND VGND VPWR VPWR cpuregs\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14822_ clknet_leaf_126_clk _00480_ VGND VGND VPWR VPWR cpuregs\[25\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ clknet_leaf_147_clk _00411_ VGND VGND VPWR VPWR cpuregs\[26\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11965_ _05768_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_739 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13704_ net1096 _06933_ _07028_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__mux2_1
X_10916_ net969 _04835_ _04959_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__mux2_1
X_14684_ clknet_leaf_157_clk _00342_ VGND VGND VPWR VPWR cpuregs\[27\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11896_ _05711_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_638 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_208 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13635_ _06996_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__clkbuf_1
X_10847_ _04931_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13566_ net1170 _06950_ _06946_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10778_ net1381 _04833_ _04887_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__mux2_1
X_15305_ clknet_leaf_32_clk _00895_ VGND VGND VPWR VPWR cpuregs\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12517_ _06264_ _06265_ _06014_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13497_ net1308 _04856_ _06899_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15236_ clknet_leaf_76_clk _00829_ VGND VGND VPWR VPWR instr_addi sky130_fd_sc_hd__dfxtp_1
X_12448_ cpuregs\[4\]\[18\] cpuregs\[5\]\[18\] _03062_ VGND VGND VPWR VPWR _06200_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15167_ clknet_leaf_56_clk _00792_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12379_ cpuregs\[0\]\[15\] cpuregs\[1\]\[15\] cpuregs\[2\]\[15\] cpuregs\[3\]\[15\]
+ _06055_ _05909_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__mux4_1
X_14118_ _01681_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15098_ clknet_leaf_100_clk _07121_ VGND VGND VPWR VPWR reg_out\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14049_ net1257 _06937_ _01638_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08610_ _03045_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__clkbuf_8
X_09590_ _03474_ _04040_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08541_ _03042_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08472_ _02340_ _03007_ _02993_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_65_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_94 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07423_ net16 _01937_ _02067_ _01935_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07354_ reg_pc\[4\] decoded_imm\[4\] VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_18_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07285_ _01931_ mem_wordsize\[2\] _01844_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_154_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09024_ cpuregs\[20\]\[1\] cpuregs\[21\]\[1\] _03405_ VGND VGND VPWR VPWR _03498_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_516 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_130_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 cpuregs\[4\]\[12\] VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_374 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold231 cpuregs\[21\]\[2\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 cpuregs\[21\]\[1\] VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 cpuregs\[1\]\[5\] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 count_cycle\[8\] VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 cpuregs\[17\]\[2\] VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 cpuregs\[3\]\[15\] VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 cpuregs\[28\]\[14\] VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ cpuregs\[28\]\[27\] cpuregs\[29\]\[27\] cpuregs\[30\]\[27\] cpuregs\[31\]\[27\]
+ _03601_ _03492_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_70_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _04304_ _04305_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__nand3_1
X_08808_ reg_out\[18\] alu_out_q\[18\] _03175_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__mux2_1
X_09788_ decoded_imm\[23\] net186 VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_29_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_104 _07064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08739_ reg_out\[9\] alu_out_q\[9\] _03174_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__mux2_1
*XANTENNA_115 reg_pc\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_126 net186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_137 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_148 net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11750_ count_cycle\[7\] count_cycle\[8\] _05607_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__and3_1
*XANTENNA_159 _03192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10701_ net717 _04844_ _04840_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_912 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11681_ _05553_ _05554_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_101_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13420_ _06867_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10632_ net774 _03302_ _04793_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10563_ _04765_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__clkbuf_1
X_13351_ net907 _04846_ _06827_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_134_663 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12302_ _06058_ _06059_ _03123_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13282_ _06794_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__clkbuf_1
X_10494_ _04728_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15021_ clknet_leaf_111_clk _00679_ VGND VGND VPWR VPWR count_cycle\[4\] sky130_fd_sc_hd__dfxtp_1
X_12233_ _03063_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_195 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12164_ _03090_ _05926_ _05927_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11115_ count_instr\[21\] _05087_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__and2_1
X_12095_ _02503_ _05861_ _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__mux2_1
X_15923_ clknet_leaf_1_clk _01495_ VGND VGND VPWR VPWR cpuregs\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_11046_ count_instr\[2\] _05037_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15854_ clknet_leaf_5_clk _01426_ VGND VGND VPWR VPWR cpuregs\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_88_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ clknet_leaf_160_clk _00463_ VGND VGND VPWR VPWR cpuregs\[25\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ clknet_leaf_8_clk _01360_ VGND VGND VPWR VPWR cpuregs\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12997_ _05041_ _06526_ _06629_ _06513_ _05804_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14736_ clknet_leaf_30_clk _00394_ VGND VGND VPWR VPWR cpuregs\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11948_ decoded_imm\[31\] net252 VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14667_ clknet_leaf_46_clk _00325_ VGND VGND VPWR VPWR cpuregs\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11879_ count_cycle\[48\] count_cycle\[49\] VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13618_ cpuregs\[31\]\[29\] _06985_ _06967_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14598_ clknet_leaf_128_clk _00256_ VGND VGND VPWR VPWR cpuregs\[28\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_764 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13549_ _03227_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__buf_2
XFILLER_0_27_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15219_ clknet_leaf_78_clk _00812_ VGND VGND VPWR VPWR instr_lui sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07972_ _02588_ _02589_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09711_ cpuregs\[12\]\[20\] cpuregs\[13\]\[20\] cpuregs\[14\]\[20\] cpuregs\[15\]\[20\]
+ _03582_ _03716_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09642_ _03414_ _04098_ _03419_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__o21a_1
X_09573_ _03397_ _04027_ _04031_ _03672_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08524_ _03042_ _03043_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08455_ _02277_ _02995_ _02993_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_766 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07406_ _01951_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08386_ _02946_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07337_ reg_pc\[3\] decoded_imm\[3\] VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_151_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07268_ _01840_ is_sb_sh_sw _01906_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09007_ _01895_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__buf_2
XFILLER_0_130_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07199_ mem_do_wdata cpu_state\[5\] _01862_ _01863_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__a31o_1
X_09909_ _04352_ _04354_ _04357_ _03575_ _03591_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a221o_1
X_12920_ decoded_imm_j\[7\] _01089_ _03169_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__mux2_1
X_12851_ instr_sh _06554_ _06539_ net647 VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_103_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ net1069 _05643_ _05647_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__o21ai_1
X_15570_ clknet_leaf_15_clk _01145_ VGND VGND VPWR VPWR cpuregs\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12782_ _06514_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__buf_1
XFILLER_0_69_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14521_ clknet_leaf_10_clk _00179_ VGND VGND VPWR VPWR cpuregs\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _05598_ _05113_ _05599_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_83_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14452_ clknet_leaf_11_clk _00110_ VGND VGND VPWR VPWR cpuregs\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11664_ _05418_ net489 _05343_ _05539_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13403_ _06858_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10615_ _04781_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_12_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14383_ clknet_leaf_31_clk _00046_ VGND VGND VPWR VPWR cpuregs\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11595_ _05463_ _05465_ _05461_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_460 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13334_ net708 _04829_ _06816_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_458 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10546_ _04756_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13265_ _06785_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__clkbuf_1
X_10477_ _04719_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__clkbuf_1
X_15004_ clknet_leaf_106_clk _00662_ VGND VGND VPWR VPWR reg_next_pc\[19\] sky130_fd_sc_hd__dfxtp_1
X_12216_ _03033_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_114_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13196_ decoded_imm\[26\] _06740_ _06737_ _06746_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_131_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12147_ _05906_ _05910_ _03124_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12078_ _05845_ _05846_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__nor2_1
X_11029_ _05027_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__clkbuf_1
X_15906_ clknet_leaf_48_clk _01478_ VGND VGND VPWR VPWR cpuregs\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15837_ clknet_leaf_17_clk _01409_ VGND VGND VPWR VPWR cpuregs\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15768_ clknet_leaf_132_clk _01343_ VGND VGND VPWR VPWR cpuregs\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14719_ clknet_leaf_97_clk _00377_ VGND VGND VPWR VPWR cpuregs\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15699_ clknet_leaf_145_clk _01274_ VGND VGND VPWR VPWR cpuregs\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08240_ net218 _02836_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_625 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_15 _02099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_26 _03149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_829 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_37 _03255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_48 _03348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08171_ _02771_ _02773_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_59 _03492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_482 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput100 net100 VGND VGND VPWR VPWR mem_la_wdata[12] sky130_fd_sc_hd__clkbuf_4
Xoutput111 net111 VGND VGND VPWR VPWR mem_la_wdata[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput122 net251 VGND VGND VPWR VPWR mem_la_wdata[3] sky130_fd_sc_hd__clkbuf_4
Xoutput133 net133 VGND VGND VPWR VPWR mem_la_wstrb[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput144 net144 VGND VGND VPWR VPWR mem_wdata[18] sky130_fd_sc_hd__clkbuf_4
Xoutput155 net155 VGND VGND VPWR VPWR mem_wdata[28] sky130_fd_sc_hd__clkbuf_4
Xoutput166 net166 VGND VGND VPWR VPWR mem_wdata[9] sky130_fd_sc_hd__clkbuf_4
Xoutput177 net177 VGND VGND VPWR VPWR pcpi_rs1[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput188 net188 VGND VGND VPWR VPWR pcpi_rs1[25] sky130_fd_sc_hd__buf_2
XFILLER_0_11_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput199 net199 VGND VGND VPWR VPWR pcpi_rs1[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_149_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07955_ _02573_ net97 _02503_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__a21oi_1
X_07886_ _02504_ _02505_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__nand2_1
X_09625_ decoded_imm\[17\] net179 VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__nor2_1
X_09556_ _03476_ _04006_ _04009_ _04015_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__a211o_1
X_08507_ mem_rdata_q\[19\] net11 _03018_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09487_ _03942_ _03944_ _03946_ _03948_ _03429_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__a221o_2
XFILLER_0_93_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08438_ _02213_ _02983_ _02971_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_202 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08369_ net249 net216 _01932_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__mux2_1
Xwire238 _02548_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10400_ cpuregs\[21\]\[5\] _03215_ _04673_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11380_ _05276_ _05277_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_586 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10331_ net879 _03215_ _04636_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__mux2_1
X_13050_ net1063 _04869_ _06658_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__mux2_1
X_10262_ _04605_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12001_ _05787_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__clkbuf_1
X_10193_ net954 _03209_ _04564_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13952_ _01593_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12903_ _05036_ _06584_ _06571_ _06585_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__nor4_1
X_13883_ _01556_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__clkbuf_1
X_15622_ clknet_leaf_36_clk _01197_ VGND VGND VPWR VPWR cpuregs\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12834_ mem_rdata_q\[13\] net5 _03017_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ clknet_leaf_27_clk _01128_ VGND VGND VPWR VPWR cpuregs\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12765_ cpu_state\[3\] _01891_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14504_ clknet_leaf_24_clk _00162_ VGND VGND VPWR VPWR cpuregs\[30\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11716_ _01889_ _05583_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__o21ai_1
X_15484_ clknet_leaf_91_clk _01069_ VGND VGND VPWR VPWR mem_rdata_q\[7\] sky130_fd_sc_hd__dfxtp_1
X_12696_ _06437_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14435_ clknet_leaf_96_clk _00093_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11647_ _05288_ _05523_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__or2_1
Xinput13 net410 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_116_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_851 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xinput24 net411 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_116_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14366_ _01810_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_133_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11578_ _05263_ net784 _05358_ _05459_ _05460_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_24_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13317_ _06812_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__clkbuf_1
Xhold808 cpuregs\[23\]\[30\] VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold819 count_instr\[18\] VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ net972 _03189_ _04746_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__mux2_1
X_14297_ net734 VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13248_ mem_rdata_q\[22\] _06627_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13179_ _06734_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__clkbuf_4
X_07740_ count_cycle\[29\] _02020_ _02361_ _02362_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__a211o_1
X_07671_ _02270_ _02285_ _02286_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__o21bai_1
X_09410_ cpuregs\[12\]\[11\] cpuregs\[13\]\[11\] cpuregs\[14\]\[11\] cpuregs\[15\]\[11\]
+ _03516_ _03409_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_144_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09341_ _03400_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09272_ _02125_ _03481_ _03661_ _03075_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08223_ _02265_ net216 _02593_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08154_ net209 net208 net207 net206 VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__or4_1
XFILLER_0_160_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08085_ net173 _02693_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08987_ cpuregs\[28\]\[0\] cpuregs\[29\]\[0\] cpuregs\[30\]\[0\] cpuregs\[31\]\[0\]
+ _03458_ _03461_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__mux4_1
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07938_ _02551_ _02553_ _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__or3_2
XFILLER_0_97_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07869_ net126 VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_3_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09608_ cpuregs\[20\]\[17\] cpuregs\[21\]\[17\] cpuregs\[22\]\[17\] cpuregs\[23\]\[17\]
+ _03516_ _03409_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10880_ net1147 _04867_ _04945_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09539_ cpuregs\[16\]\[15\] cpuregs\[17\]\[15\] cpuregs\[18\]\[15\] cpuregs\[19\]\[15\]
+ _03598_ _03460_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_80_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12550_ _05974_ cpuregs\[30\]\[22\] _05896_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_678 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_108_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11501_ _05285_ _05216_ _05389_ _05300_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__a22o_1
X_12481_ _06138_ _06231_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14220_ _01735_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__clkbuf_1
X_11432_ _05273_ _05204_ _05184_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14151_ cpuregs\[7\]\[22\] _06971_ _01696_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11363_ _05031_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_78_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13102_ _06693_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__clkbuf_1
X_10314_ _04632_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_95_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14082_ _01662_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__clkbuf_1
X_11294_ _02946_ _03257_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ net1072 _04852_ _06647_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__mux2_1
X_10245_ net1122 _03374_ _04586_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10176_ _04558_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14984_ clknet_leaf_86_clk _00642_ VGND VGND VPWR VPWR reg_pc\[30\] sky130_fd_sc_hd__dfxtp_2
X_13935_ _01584_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_161_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13866_ _01547_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__clkbuf_1
X_15605_ clknet_leaf_144_clk _01180_ VGND VGND VPWR VPWR cpuregs\[31\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12817_ _06528_ _06538_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13797_ net853 _06958_ _07075_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__mux2_1
X_15536_ clknet_leaf_150_clk _01121_ VGND VGND VPWR VPWR cpuregs\[24\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12748_ _03143_ _06486_ _06182_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__o21a_1
XFILLER_0_155_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15467_ clknet_leaf_151_clk _01057_ VGND VGND VPWR VPWR cpuregs\[19\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12679_ _06419_ _06420_ _03082_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14418_ clknet_leaf_62_clk _00076_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dfxtp_4
X_15398_ clknet_leaf_87_clk _00988_ VGND VGND VPWR VPWR decoded_imm\[10\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_142_558 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14349_ cpuregs\[10\]\[21\] _03321_ _01800_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__mux2_1
Xhold605 cpuregs\[18\]\[24\] VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 cpuregs\[11\]\[1\] VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 mem_rdata[2] VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 cpuregs\[31\]\[10\] VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 count_instr\[41\] VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08910_ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_792 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09890_ _04282_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08841_ reg_pc\[22\] reg_pc\[21\] _03311_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ reg_pc\[13\] _03259_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07723_ count_instr\[60\] _02052_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07654_ count_instr\[55\] _01946_ _02054_ net518 VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07585_ _02217_ _02218_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09324_ reg_pc\[8\] _03527_ _03625_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09255_ _03593_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08206_ _02762_ _02771_ _02772_ _02802_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__a211o_1
XFILLER_0_141_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09186_ _03074_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__buf_2
XFILLER_0_161_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08137_ _02466_ _02727_ _02573_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08068_ _02482_ _02476_ _02657_ _02573_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__o31a_1
XFILLER_0_12_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10030_ cpuregs\[0\]\[30\] cpuregs\[1\]\[30\] cpuregs\[2\]\[30\] cpuregs\[3\]\[30\]
+ _03673_ _03451_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_8_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11981_ net35 net66 _05774_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__mux2_1
X_13720_ _07041_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__clkbuf_1
X_10932_ _04976_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13651_ net1024 _06948_ _07003_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__mux2_1
X_10863_ net834 _04850_ _04934_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12602_ _06347_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13582_ _06961_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__clkbuf_1
X_10794_ _04903_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15321_ clknet_leaf_132_clk _00911_ VGND VGND VPWR VPWR cpuregs\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_795 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_155_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12533_ _05862_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15252_ clknet_leaf_80_clk _00845_ VGND VGND VPWR VPWR instr_sra sky130_fd_sc_hd__dfxtp_1
X_12464_ _06213_ _06214_ _06215_ _05873_ _03113_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14203_ _01726_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11415_ _05309_ _05310_ _05185_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__a21o_1
X_15183_ clknet_leaf_82_clk _00808_ VGND VGND VPWR VPWR latched_branch sky130_fd_sc_hd__dfxtp_2
X_12395_ _06073_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_22_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14134_ cpuregs\[7\]\[14\] _06954_ _01685_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11346_ reg_next_pc\[27\] _03357_ _02948_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14065_ _01653_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__clkbuf_1
X_11277_ _05186_ _05201_ _05202_ _01885_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__o211a_1
X_13016_ net1065 _04835_ _06636_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__mux2_1
X_10228_ _04587_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10159_ net1080 _03322_ _04548_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14967_ clknet_leaf_105_clk _00625_ VGND VGND VPWR VPWR reg_pc\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_77_707 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_89_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13918_ _01575_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_141_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14898_ clknet_leaf_112_clk _00556_ VGND VGND VPWR VPWR count_instr\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13849_ _07109_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07370_ _02017_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_604 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_57_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15519_ clknet_leaf_156_clk _01104_ VGND VGND VPWR VPWR cpuregs\[24\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_40_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09040_ _03510_ _03512_ _03513_ _03403_ _03420_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold402 net46 VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold413 cpuregs\[16\]\[21\] VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 cpuregs\[11\]\[25\] VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 cpuregs\[10\]\[29\] VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 cpuregs\[23\]\[28\] VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 cpuregs\[11\]\[0\] VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 cpuregs\[25\]\[24\] VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _03476_ _04379_ _04383_ _04389_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__a211o_1
Xhold479 cpuregs\[30\]\[24\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09873_ cpuregs\[24\]\[25\] cpuregs\[25\]\[25\] cpuregs\[26\]\[25\] cpuregs\[27\]\[25\]
+ _03808_ _03812_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_55_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ reg_pc\[20\] reg_pc\[19\] _03299_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__and3_1
X_08755_ reg_out\[11\] alu_out_q\[11\] _03174_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__mux2_2
X_07706_ net19 _02202_ _02179_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__a21o_1
X_08686_ _01971_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07637_ _02058_ _02264_ _02267_ _01968_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07568_ _02065_ _02200_ _02201_ _02203_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09307_ _03670_ _03772_ _03773_ _01943_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07499_ net174 VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_683 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09238_ _03704_ _03706_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09169_ _03404_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__buf_6
XFILLER_0_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11200_ count_instr\[47\] _05146_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12180_ cpuregs\[8\]\[7\] cpuregs\[9\]\[7\] cpuregs\[10\]\[7\] cpuregs\[11\]\[7\]
+ _03150_ _05917_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_364 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11131_ count_instr\[26\] _05095_ _05098_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold980 cpuregs\[5\]\[24\] VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 cpuregs\[24\]\[20\] VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ _05036_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__buf_4
XFILLER_0_101_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10013_ _04381_ _04392_ _03483_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__o21ai_1
X_15870_ clknet_leaf_129_clk _01442_ VGND VGND VPWR VPWR cpuregs\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_14821_ clknet_leaf_150_clk _00479_ VGND VGND VPWR VPWR cpuregs\[25\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ clknet_leaf_149_clk _00410_ VGND VGND VPWR VPWR cpuregs\[26\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ net1292 net86 _05767_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13703_ _07032_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__clkbuf_1
X_10915_ _04967_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__clkbuf_1
X_14683_ clknet_leaf_160_clk _00341_ VGND VGND VPWR VPWR cpuregs\[27\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_11895_ _01884_ _05709_ _05710_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__and3_1
X_13634_ cpuregs\[23\]\[3\] _06931_ _06992_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__mux2_1
X_10846_ net1139 _04833_ _04923_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13565_ _03262_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__clkbuf_4
X_10777_ _04894_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15304_ clknet_leaf_56_clk _00894_ VGND VGND VPWR VPWR cpuregs\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12516_ cpuregs\[0\]\[21\] cpuregs\[1\]\[21\] cpuregs\[2\]\[21\] cpuregs\[3\]\[21\]
+ _06055_ _05829_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13496_ _06907_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__clkbuf_1
X_15235_ clknet_leaf_77_clk net648 VGND VGND VPWR VPWR instr_sh sky130_fd_sc_hd__dfxtp_1
X_12447_ _06199_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_686 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15166_ clknet_leaf_51_clk _00791_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dfxtp_4
X_12378_ cpuregs\[4\]\[15\] cpuregs\[5\]\[15\] cpuregs\[6\]\[15\] cpuregs\[7\]\[15\]
+ _06011_ _03097_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14117_ cpuregs\[7\]\[6\] _06937_ _01674_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__mux2_1
X_11329_ _01842_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15097_ clknet_leaf_100_clk _07120_ VGND VGND VPWR VPWR reg_out\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14048_ _01644_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08540_ _03050_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__or2_1
X_08471_ reg_next_pc\[27\] reg_out\[27\] _02991_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07422_ net7 net25 _01844_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07353_ _01988_ _01975_ _01986_ _02000_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__o31a_1
XFILLER_0_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_61_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07284_ net31 net17 _01845_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09023_ _03496_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_131_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold210 net61 VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold221 cpuregs\[2\]\[0\] VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold232 cpuregs\[7\]\[4\] VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold243 instr_slli VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 cpuregs\[0\]\[5\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold265 instr_xori VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 instr_sll VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 cpuregs\[25\]\[16\] VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09925_ _03581_ _04372_ _03547_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__o21a_1
Xhold298 cpuregs\[27\]\[19\] VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ decoded_imm\[24\] _02306_ _04282_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_0_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08807_ _03296_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_37_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09787_ decoded_imm\[23\] net186 VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _03236_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
*XANTENNA_105 _07100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_116 reg_pc\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_127 net186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_138 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08669_ _03175_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__buf_4
*XANTENNA_149 _01674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10700_ _03262_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11680_ _05530_ _05532_ _05533_ _05543_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_924 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10631_ _04801_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13350_ _06830_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__clkbuf_1
X_10562_ net1109 _03295_ _04757_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_404 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12301_ cpuregs\[12\]\[12\] cpuregs\[13\]\[12\] cpuregs\[14\]\[12\] cpuregs\[15\]\[12\]
+ _05913_ _05994_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__mux4_1
X_13281_ net1226 _04844_ _06791_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10493_ cpuregs\[14\]\[17\] _03295_ _04720_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__mux2_1
X_15020_ clknet_leaf_111_clk _00678_ VGND VGND VPWR VPWR count_cycle\[3\] sky130_fd_sc_hd__dfxtp_1
X_12232_ _05991_ _05992_ _03124_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12163_ _03034_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__buf_4
XFILLER_0_130_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11114_ _05087_ _05088_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__nor2_1
X_12094_ _05862_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__buf_4
X_15922_ clknet_leaf_6_clk _01494_ VGND VGND VPWR VPWR cpuregs\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11045_ net494 _05033_ _05038_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15853_ clknet_leaf_7_clk _01425_ VGND VGND VPWR VPWR cpuregs\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_88_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ clknet_leaf_159_clk _00462_ VGND VGND VPWR VPWR cpuregs\[25\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15784_ clknet_leaf_32_clk _01359_ VGND VGND VPWR VPWR cpuregs\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ net1133 _06626_ _06632_ _06634_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_857 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11947_ _01953_ _03770_ _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__and3_1
X_14735_ clknet_leaf_43_clk _00393_ VGND VGND VPWR VPWR cpuregs\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14666_ clknet_leaf_45_clk _00324_ VGND VGND VPWR VPWR cpuregs\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11878_ net479 _05695_ _05698_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13617_ _03373_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_918 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10829_ _04921_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__clkbuf_1
X_14597_ clknet_leaf_144_clk _00255_ VGND VGND VPWR VPWR cpuregs\[28\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_916 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13548_ _06938_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_631 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_15_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_501 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13479_ _06898_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_623 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15218_ clknet_leaf_71_clk alu_out\[31\] VGND VGND VPWR VPWR alu_out_q\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15149_ clknet_leaf_70_clk _00774_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_2_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07971_ net193 _02587_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__or2_1
X_09710_ _03433_ _04160_ _04162_ _04164_ _03760_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09641_ cpuregs\[24\]\[18\] cpuregs\[25\]\[18\] cpuregs\[26\]\[18\] cpuregs\[27\]\[18\]
+ _03640_ _03496_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__mux4_1
X_09572_ _03483_ _03952_ _04028_ _04030_ _01958_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__o311a_1
XFILLER_0_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08523_ cpuregs\[16\]\[2\] cpuregs\[17\]\[2\] cpuregs\[18\]\[2\] cpuregs\[19\]\[2\]
+ _03038_ _03039_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08454_ reg_next_pc\[22\] reg_out\[22\] _02991_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07405_ _02043_ _02048_ _02050_ _02018_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__o22a_1
XFILLER_0_148_778 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08385_ _02945_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__clkbuf_4
X_07336_ _01970_ _01974_ _01976_ _01985_ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07267_ net1409 _01921_ _01922_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09006_ _03480_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07198_ mem_do_rdata cpu_state\[6\] _01862_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09908_ _04355_ _04356_ _03579_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__mux2_1
X_09839_ cpuregs\[0\]\[24\] cpuregs\[1\]\[24\] cpuregs\[2\]\[24\] cpuregs\[3\]\[24\]
+ _03641_ _03642_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12850_ net673 _06554_ _06535_ net647 VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _05040_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__clkbuf_4
X_12781_ mem_rdata_q\[3\] net26 _03017_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__mux2_1
X_14520_ clknet_leaf_17_clk _00178_ VGND VGND VPWR VPWR cpuregs\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11732_ count_cycle\[0\] count_cycle\[1\] count_cycle\[2\] VGND VGND VPWR VPWR _05599_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_83_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14451_ clknet_leaf_31_clk _00109_ VGND VGND VPWR VPWR cpuregs\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_54_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11663_ _05537_ _05538_ _05185_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13402_ net946 _04829_ _06852_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__mux2_1
X_10614_ _04792_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14382_ clknet_leaf_58_clk _00045_ VGND VGND VPWR VPWR cpuregs\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11594_ _05473_ _05474_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13333_ _06821_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10545_ cpuregs\[27\]\[9\] _03241_ _04746_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_130_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_130_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13264_ net722 _04827_ _06780_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__mux2_1
X_10476_ net1260 _03241_ _04709_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__mux2_1
X_15003_ clknet_leaf_107_clk _00661_ VGND VGND VPWR VPWR reg_next_pc\[18\] sky130_fd_sc_hd__dfxtp_1
X_12215_ _05973_ _05975_ _05976_ _05873_ _03113_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_114_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13195_ mem_rdata_q\[26\] _06742_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12146_ cpuregs\[0\]\[6\] cpuregs\[1\]\[6\] cpuregs\[2\]\[6\] cpuregs\[3\]\[6\] _05908_
+ _05909_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_63_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12077_ cpuregs\[4\]\[1\] cpuregs\[5\]\[1\] cpuregs\[6\]\[1\] cpuregs\[7\]\[1\] _03107_
+ _03108_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__mux4_1
X_11028_ net1281 _04879_ _05017_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__mux2_1
X_15905_ clknet_leaf_21_clk _01477_ VGND VGND VPWR VPWR cpuregs\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15836_ clknet_leaf_142_clk _01408_ VGND VGND VPWR VPWR cpuregs\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15767_ clknet_leaf_134_clk _01342_ VGND VGND VPWR VPWR cpuregs\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12979_ _06624_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
X_14718_ clknet_leaf_21_clk _00376_ VGND VGND VPWR VPWR cpuregs\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_72_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15698_ clknet_leaf_3_clk _01273_ VGND VGND VPWR VPWR cpuregs\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14649_ clknet_leaf_10_clk _00307_ VGND VGND VPWR VPWR cpuregs\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_16 _02949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_637 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_27 _03150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_38 _03257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08170_ _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__inv_2
*XANTENNA_49 _03402_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_121_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_121_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_113_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_634 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_125_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput101 net101 VGND VGND VPWR VPWR mem_la_wdata[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput112 net112 VGND VGND VPWR VPWR mem_la_wdata[23] sky130_fd_sc_hd__buf_2
XFILLER_0_51_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput123 net123 VGND VGND VPWR VPWR mem_la_wdata[4] sky130_fd_sc_hd__clkbuf_4
Xoutput134 net134 VGND VGND VPWR VPWR mem_valid sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput145 net145 VGND VGND VPWR VPWR mem_wdata[19] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_81_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput156 net156 VGND VGND VPWR VPWR mem_wdata[29] sky130_fd_sc_hd__clkbuf_4
Xoutput167 net167 VGND VGND VPWR VPWR mem_wstrb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput178 net178 VGND VGND VPWR VPWR pcpi_rs1[16] sky130_fd_sc_hd__clkbuf_4
Xoutput189 net189 VGND VGND VPWR VPWR pcpi_rs1[26] sky130_fd_sc_hd__buf_2
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07954_ _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_149_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07885_ _01844_ _02503_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__nand2_1
X_09624_ _04057_ _04076_ _04081_ _03396_ _02213_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__o32a_1
X_09555_ _04013_ _04014_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_90_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08506_ _03029_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__clkbuf_1
X_09486_ _03435_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_65_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_827 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08437_ reg_next_pc\[17\] reg_out\[17\] _02969_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__mux2_2
XFILLER_0_135_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08368_ _02940_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_1
XFILLER_0_160_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_212 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xwire239 _06583_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_1
X_07319_ _01969_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_908 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_112_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_112_clk sky130_fd_sc_hd__clkbuf_2
X_08299_ net223 _02890_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__xor2_1
XFILLER_0_132_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10330_ _04641_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10261_ net815 _03209_ _04600_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__mux2_1
X_12000_ net519 net75 _05785_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__mux2_1
X_10192_ _04568_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__clkbuf_1
X_13951_ net744 _06975_ _01588_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12902_ mem_rdata_q\[4\] mem_rdata_q\[5\] mem_rdata_q\[6\] mem_rdata_q\[3\] VGND
+ VGND VPWR VPWR _06585_ sky130_fd_sc_hd__or4b_1
X_13882_ net753 _06975_ _01551_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_129_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15621_ clknet_leaf_33_clk _01196_ VGND VGND VPWR VPWR cpuregs\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12833_ _06549_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__buf_1
XFILLER_0_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12764_ _05185_ _02071_ _01840_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__a21oi_1
X_15552_ clknet_leaf_51_clk _01127_ VGND VGND VPWR VPWR cpuregs\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14503_ clknet_leaf_130_clk _00161_ VGND VGND VPWR VPWR cpuregs\[30\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11715_ _05367_ _05584_ _05585_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__or3b_1
X_15483_ clknet_leaf_83_clk _01068_ VGND VGND VPWR VPWR mem_rdata_q\[6\] sky130_fd_sc_hd__dfxtp_1
X_12695_ net223 _06436_ _06282_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__mux2_1
X_11646_ _05244_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__nor2_1
X_14434_ clknet_leaf_60_clk _00092_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_126_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput14 net485 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ net794 _03373_ _01800_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__mux2_1
Xinput25 mem_rdata[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_103_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_103_clk sky130_fd_sc_hd__clkbuf_2
X_11577_ _05184_ _05230_ _05449_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_133_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_554 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13316_ cpuregs\[18\]\[29\] _04879_ _06802_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10528_ _04747_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__clkbuf_1
X_14296_ _01773_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__clkbuf_1
Xhold809 cpuregs\[6\]\[18\] VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13247_ net689 _06531_ _06773_ _06774_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__o22a_1
X_10459_ _04710_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13178_ mem_rdata_q\[31\] _06733_ _06540_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__a21o_1
X_12129_ cpuregs\[12\]\[5\] cpuregs\[13\]\[5\] cpuregs\[14\]\[5\] cpuregs\[15\]\[5\]
+ _03096_ _03098_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__mux4_1
X_07670_ _02260_ _02271_ _02272_ _02287_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_144_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15819_ clknet_leaf_32_clk _01391_ VGND VGND VPWR VPWR cpuregs\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09340_ _03557_ _03805_ _03417_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_36_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09271_ _03736_ _03738_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_715 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08222_ _02818_ _02819_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_60_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08153_ _02656_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__buf_2
XFILLER_0_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08084_ net205 _02692_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08986_ _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__clkbuf_8
X_07937_ net238 _02554_ _02556_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__o21a_1
X_07868_ _02477_ _02478_ _02481_ _02487_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09607_ _03427_ _04060_ _04062_ _04064_ _03490_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__a221o_2
X_07799_ _02417_ _02418_ net247 VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__a21bo_1
X_09538_ _03593_ _03997_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09469_ _03894_ _03902_ _03930_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11500_ _05289_ _05384_ _05385_ _05386_ _05388_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__a32o_1
X_12480_ cpuregs\[8\]\[19\] cpuregs\[9\]\[19\] cpuregs\[10\]\[19\] cpuregs\[11\]\[19\]
+ _06061_ _05917_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11431_ _05323_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14150_ _01698_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_885 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11362_ _05185_ _05261_ _05262_ _05257_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_78_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13101_ net619 _02489_ _06685_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ cpuregs\[2\]\[29\] _03374_ _04622_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14081_ net1336 _06969_ _01660_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11293_ _05194_ reg_pc\[11\] _01843_ _05213_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_95_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13032_ _06653_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__clkbuf_1
X_10244_ _04595_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__clkbuf_1
X_10175_ net1061 _03374_ _04548_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__mux2_1
X_14983_ clknet_leaf_106_clk _00641_ VGND VGND VPWR VPWR reg_pc\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13934_ net1029 _06958_ _01577_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_161_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13865_ net1393 _06958_ _07111_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15604_ clknet_leaf_121_clk _01179_ VGND VGND VPWR VPWR cpuregs\[31\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12816_ _06532_ _06537_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13796_ _07081_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15535_ clknet_leaf_149_clk _01120_ VGND VGND VPWR VPWR cpuregs\[24\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12747_ cpuregs\[12\]\[31\] cpuregs\[13\]\[31\] cpuregs\[14\]\[31\] cpuregs\[15\]\[31\]
+ _03133_ _03134_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15466_ clknet_leaf_150_clk _01056_ VGND VGND VPWR VPWR cpuregs\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_12678_ cpuregs\[0\]\[28\] cpuregs\[1\]\[28\] cpuregs\[2\]\[28\] cpuregs\[3\]\[28\]
+ _03091_ _05829_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11629_ _05237_ _05240_ _05494_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__o21a_1
X_14417_ clknet_leaf_62_clk _00075_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_42_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15397_ clknet_leaf_82_clk _00987_ VGND VGND VPWR VPWR decoded_imm\[11\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14348_ _01801_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__clkbuf_1
Xhold606 cpuregs\[22\]\[8\] VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 cpuregs\[21\]\[0\] VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 cpuregs\[10\]\[10\] VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ net654 VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__clkbuf_1
Xhold639 cpuregs\[24\]\[10\] VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_760 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08840_ reg_pc\[22\] _03319_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_146_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ reg_out\[13\] alu_out_q\[13\] _03174_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__mux2_1
X_07722_ _02343_ net488 VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07653_ _02071_ _02276_ _02279_ _02282_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_0_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07584_ reg_pc\[18\] decoded_imm\[18\] VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09323_ _03434_ _03785_ _03787_ _03789_ _03431_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09254_ cpuregs\[12\]\[6\] cpuregs\[13\]\[6\] cpuregs\[14\]\[6\] cpuregs\[15\]\[6\]
+ _03587_ _03442_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08205_ _02237_ _02793_ _02804_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09185_ _03613_ _03612_ _03654_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__or3b_1
XFILLER_0_141_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_16_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08136_ _02468_ _02581_ _02740_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_389 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08067_ _02585_ _02674_ _02677_ VGND VGND VPWR VPWR alu_out\[9\] sky130_fd_sc_hd__a21o_1
XFILLER_0_12_793 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08969_ cpuregs\[16\]\[0\] cpuregs\[17\]\[0\] cpuregs\[18\]\[0\] cpuregs\[19\]\[0\]
+ _03440_ _03443_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__mux4_1
X_11980_ _05776_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__clkbuf_1
X_10931_ net1118 _04850_ _04970_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13650_ _07004_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__clkbuf_1
X_10862_ _04939_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_78_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12601_ net219 _06346_ _06282_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__mux2_1
X_13581_ net1217 _06960_ _06946_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__mux2_1
X_10793_ net970 _04848_ _04898_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_819 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_692 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15320_ clknet_leaf_130_clk _00910_ VGND VGND VPWR VPWR cpuregs\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12532_ _06132_ _06271_ _06280_ _06153_ decoded_imm\[21\] VGND VGND VPWR VPWR _06281_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_152_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12463_ cpuregs\[28\]\[18\] cpuregs\[29\]\[18\] _03085_ VGND VGND VPWR VPWR _06215_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15251_ clknet_leaf_80_clk _00844_ VGND VGND VPWR VPWR instr_srl sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14202_ cpuregs\[8\]\[14\] _06954_ _01721_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__mux2_1
X_11414_ _05273_ _05297_ _05199_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__o21bai_1
X_15182_ clknet_leaf_81_clk _00807_ VGND VGND VPWR VPWR latched_stalu sky130_fd_sc_hd__dfxtp_2
X_12394_ cpuregs\[24\]\[15\] cpuregs\[25\]\[15\] cpuregs\[26\]\[15\] cpuregs\[27\]\[15\]
+ _06074_ _05932_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__mux4_1
X_14133_ _01689_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11345_ _05194_ net795 _05239_ _05250_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__o211a_1
X_14064_ net1333 _06952_ _01649_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__mux2_1
X_11276_ _05188_ reg_pc\[6\] VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__or2_1
X_13015_ _06644_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__clkbuf_1
X_10227_ net1150 _03314_ _04586_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10158_ _04549_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10089_ _04511_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__clkbuf_1
X_14966_ clknet_leaf_87_clk _00624_ VGND VGND VPWR VPWR reg_pc\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_546 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13917_ net1090 _06941_ _01566_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14897_ clknet_leaf_112_clk _00555_ VGND VGND VPWR VPWR count_instr\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13848_ net965 _06941_ _07100_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13779_ _07072_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15518_ clknet_leaf_29_clk _01103_ VGND VGND VPWR VPWR cpuregs\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15449_ clknet_leaf_29_clk _01039_ VGND VGND VPWR VPWR cpuregs\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_682 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold403 cpuregs\[17\]\[21\] VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold414 cpuregs\[27\]\[25\] VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold425 reg_next_pc\[18\] VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 reg_pc\[26\] VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold447 cpuregs\[13\]\[18\] VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 cpuregs\[3\]\[30\] VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 cpuregs\[22\]\[28\] VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _01870_ _04387_ _04388_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09872_ _03446_ _04321_ _03417_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_55_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ reg_pc\[19\] _03299_ reg_pc\[20\] VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08754_ _03250_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__clkbuf_1
X_07705_ net189 VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__buf_4
X_08685_ _03190_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_92_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_2
X_07636_ _02065_ _02265_ _02184_ _02266_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07567_ net8 _02202_ _02180_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_24_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09306_ _02139_ _03481_ _03669_ _03075_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07498_ _02134_ _02136_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_744 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09237_ _03652_ _03655_ _03705_ _03697_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09168_ _03500_ _03638_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08119_ _02154_ _02471_ _02724_ _02725_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_75_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09099_ _03397_ _03542_ _03543_ _03571_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__a31o_1
XFILLER_0_160_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11130_ _05095_ _05098_ _05099_ _05052_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__a211oi_1
Xhold970 reg_next_pc\[2\] VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 cpuregs\[18\]\[25\] VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ count_instr\[3\] count_instr\[2\] _05037_ _05050_ VGND VGND VPWR VPWR _05051_
+ sky130_fd_sc_hd__and4_1
Xhold992 cpuregs\[29\]\[31\] VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10012_ _04425_ _04455_ _04454_ _04453_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__o211ai_2
X_14820_ clknet_leaf_149_clk _00478_ VGND VGND VPWR VPWR cpuregs\[25\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_844 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14751_ clknet_leaf_125_clk _00409_ VGND VGND VPWR VPWR cpuregs\[26\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_123_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_2
X_13702_ net1261 _06931_ _07028_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__mux2_1
X_10914_ net1392 _04833_ _04959_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__mux2_1
X_14682_ clknet_leaf_155_clk _00340_ VGND VGND VPWR VPWR cpuregs\[27\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11894_ net1399 _05706_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__nand2_1
X_10845_ _04930_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__clkbuf_1
X_13633_ _06995_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13564_ _06949_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10776_ net1297 _04831_ _04887_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__mux2_1
X_15303_ clknet_leaf_34_clk _00893_ VGND VGND VPWR VPWR cpuregs\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12515_ cpuregs\[4\]\[21\] cpuregs\[5\]\[21\] cpuregs\[6\]\[21\] cpuregs\[7\]\[21\]
+ _06011_ _06156_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__mux4_1
X_13495_ net971 _04854_ _06899_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12446_ net211 _06198_ _06052_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__mux2_1
X_15234_ clknet_leaf_77_clk _00827_ VGND VGND VPWR VPWR instr_sb sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_507 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_23_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12377_ _05900_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__clkbuf_4
X_15165_ clknet_leaf_51_clk _00790_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_140_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11328_ _05227_ _05237_ _05238_ _05224_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__o211a_1
X_14116_ _01680_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__clkbuf_1
X_15096_ clknet_leaf_104_clk _07119_ VGND VGND VPWR VPWR reg_out\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11259_ _05186_ _05187_ _05189_ _01885_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14047_ cpuregs\[6\]\[5\] _06935_ _01638_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14949_ clknet_leaf_118_clk _00607_ VGND VGND VPWR VPWR count_instr\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_2
X_08470_ _03006_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_1
XFILLER_0_148_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07421_ net200 VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07352_ reg_pc\[3\] decoded_imm\[3\] VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_662 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07283_ net171 mem_wordsize\[1\] VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__and2_2
XFILLER_0_5_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09022_ _03408_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold200 count_instr\[24\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold211 count_cycle\[13\] VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold222 cpuregs\[0\]\[22\] VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold233 cpuregs\[0\]\[21\] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 cpuregs\[14\]\[12\] VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 cpuregs\[0\]\[16\] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 cpuregs\[30\]\[1\] VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 cpuregs\[7\]\[5\] VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 is_sb_sh_sw VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__buf_1
Xhold299 cpuregs\[24\]\[16\] VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ cpuregs\[16\]\[27\] cpuregs\[17\]\[27\] cpuregs\[18\]\[27\] cpuregs\[19\]\[27\]
+ _03598_ _03460_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ decoded_imm\[25\] net188 VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__or2_2
X_08806_ cpuregs\[11\]\[17\] _03295_ _03249_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09786_ _04215_ _04216_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_29_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ net880 _03235_ _03185_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_106 decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
*XANTENNA_117 reg_pc\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_128 net187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_139 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08668_ _03174_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07619_ _01932_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__buf_4
X_08599_ _03104_ _03111_ _03116_ net244 VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_936 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10630_ net683 _03295_ _04793_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10561_ _04764_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12300_ _03153_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13280_ _06793_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_101_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10492_ _04727_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12231_ cpuregs\[0\]\[9\] cpuregs\[1\]\[9\] cpuregs\[2\]\[9\] cpuregs\[3\]\[9\] _05908_
+ _05909_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__mux4_1
X_12162_ cpuregs\[16\]\[6\] cpuregs\[17\]\[6\] cpuregs\[18\]\[6\] cpuregs\[19\]\[6\]
+ _03133_ _05925_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__mux4_1
X_11113_ net516 _05085_ _05044_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__o21ai_1
X_12093_ _01839_ _01840_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__and2_2
X_11044_ _05036_ _05037_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__nor2_1
X_15921_ clknet_leaf_9_clk _01493_ VGND VGND VPWR VPWR cpuregs\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_110_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15852_ clknet_leaf_8_clk _01424_ VGND VGND VPWR VPWR cpuregs\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14803_ clknet_leaf_29_clk _00461_ VGND VGND VPWR VPWR cpuregs\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15783_ clknet_leaf_55_clk _01358_ VGND VGND VPWR VPWR cpuregs\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_56_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_2
X_12995_ is_sll_srl_sra _06541_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14734_ clknet_leaf_45_clk _00392_ VGND VGND VPWR VPWR cpuregs\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11946_ _02340_ _02380_ _03073_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ clknet_leaf_21_clk _00323_ VGND VGND VPWR VPWR cpuregs\[14\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_11877_ net479 _05695_ _01905_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13616_ _06984_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__clkbuf_1
X_10828_ net890 _04883_ _04886_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__mux2_1
X_14596_ clknet_leaf_145_clk _00254_ VGND VGND VPWR VPWR cpuregs\[28\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13547_ net1099 _06937_ _06925_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_928 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10759_ net856 _04883_ _04818_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13478_ net835 _04837_ _06888_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_513 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15217_ clknet_leaf_73_clk alu_out\[30\] VGND VGND VPWR VPWR alu_out_q\[30\] sky130_fd_sc_hd__dfxtp_1
X_12429_ _03054_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__buf_4
XFILLER_0_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_557 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15148_ clknet_leaf_82_clk _00000_ VGND VGND VPWR VPWR decoder_trigger sky130_fd_sc_hd__dfxtp_4
XFILLER_0_77_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07970_ net193 _02587_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__nand2_1
X_15079_ clknet_leaf_117_clk _00737_ VGND VGND VPWR VPWR count_cycle\[62\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09640_ _04095_ _04096_ _03579_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09571_ _03953_ _04029_ _03483_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_47_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_2
X_08522_ _00009_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_195 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08453_ _02994_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_1
X_07404_ count_instr\[38\] _02013_ count_cycle\[6\] _01951_ _02049_ VGND VGND VPWR
+ VPWR _02050_ sky130_fd_sc_hd__a221o_2
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08384_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__buf_2
XFILLER_0_135_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07335_ _01977_ _01978_ _01981_ _01928_ _01984_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07266_ _01905_ _01851_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__nand2_1
X_09005_ _03479_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__buf_2
XFILLER_0_131_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07197_ mem_do_prefetch _01861_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__nand2_2
XFILLER_0_130_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_111_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09907_ cpuregs\[0\]\[26\] cpuregs\[1\]\[26\] cpuregs\[2\]\[26\] cpuregs\[3\]\[26\]
+ _03457_ _03595_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__mux4_1
X_09838_ cpuregs\[4\]\[24\] cpuregs\[5\]\[24\] cpuregs\[6\]\[24\] cpuregs\[7\]\[24\]
+ _03641_ _03642_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__mux4_1
X_09769_ cpuregs\[24\]\[22\] cpuregs\[25\]\[22\] cpuregs\[26\]\[22\] cpuregs\[27\]\[22\]
+ _03640_ _03492_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_38_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_103_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ count_cycle\[22\] count_cycle\[23\] _05640_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12780_ _06512_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__buf_2
XFILLER_0_139_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11731_ count_cycle\[0\] count_cycle\[1\] count_cycle\[2\] VGND VGND VPWR VPWR _05598_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_83_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ clknet_leaf_57_clk _00108_ VGND VGND VPWR VPWR cpuregs\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11662_ _05032_ _05524_ _05246_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13401_ _06857_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__clkbuf_1
X_10613_ net858 _03241_ _04782_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__mux2_1
X_11593_ decoded_imm_j\[20\] _05235_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__or2_1
X_14381_ clknet_leaf_35_clk _00044_ VGND VGND VPWR VPWR cpuregs\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10544_ _04755_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13332_ net767 _04827_ _06816_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13263_ _06784_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__clkbuf_1
X_10475_ _04718_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15002_ clknet_leaf_107_clk _00660_ VGND VGND VPWR VPWR reg_next_pc\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12214_ cpuregs\[28\]\[8\] cpuregs\[29\]\[8\] _03085_ VGND VGND VPWR VPWR _05976_
+ sky130_fd_sc_hd__mux2_1
X_13194_ decoded_imm\[27\] _06740_ _06737_ _06745_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_131_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12145_ _03047_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_131_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12076_ _03050_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__buf_4
X_11027_ _05026_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__clkbuf_1
X_15904_ clknet_leaf_21_clk _01476_ VGND VGND VPWR VPWR cpuregs\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15835_ clknet_leaf_132_clk _01407_ VGND VGND VPWR VPWR cpuregs\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_29_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_2
X_15766_ clknet_leaf_135_clk _01341_ VGND VGND VPWR VPWR cpuregs\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12978_ decoded_imm_j\[2\] _01084_ _03021_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__mux2_1
X_14717_ clknet_leaf_13_clk _00375_ VGND VGND VPWR VPWR cpuregs\[15\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11929_ cpuregs\[0\]\[31\] cpuregs\[1\]\[31\] cpuregs\[2\]\[31\] cpuregs\[3\]\[31\]
+ _03404_ _03576_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__mux4_1
X_15697_ clknet_leaf_16_clk _01272_ VGND VGND VPWR VPWR cpuregs\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_880 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14648_ clknet_leaf_17_clk _00306_ VGND VGND VPWR VPWR cpuregs\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_17 _03085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
*XANTENNA_28 _03151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_649 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_39 _03262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14579_ clknet_leaf_30_clk _00237_ VGND VGND VPWR VPWR cpuregs\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput102 net102 VGND VGND VPWR VPWR mem_la_wdata[14] sky130_fd_sc_hd__buf_2
Xoutput113 net113 VGND VGND VPWR VPWR mem_la_wdata[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput124 net124 VGND VGND VPWR VPWR mem_la_wdata[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput135 net135 VGND VGND VPWR VPWR mem_wdata[0] sky130_fd_sc_hd__buf_2
XFILLER_0_88_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput146 net146 VGND VGND VPWR VPWR mem_wdata[1] sky130_fd_sc_hd__clkbuf_4
Xoutput157 net157 VGND VGND VPWR VPWR mem_wdata[2] sky130_fd_sc_hd__clkbuf_4
Xoutput168 net168 VGND VGND VPWR VPWR mem_wstrb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput179 net179 VGND VGND VPWR VPWR pcpi_rs1[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07953_ instr_sub VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07884_ net182 _02503_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__or2_1
X_09623_ _01977_ _04078_ _04080_ _03486_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__a31o_1
X_09554_ _03962_ _03967_ _04012_ _01869_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__a31o_1
X_08505_ decoded_imm_j\[18\] _01080_ _03022_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09485_ cpuregs\[24\]\[13\] cpuregs\[25\]\[13\] cpuregs\[26\]\[13\] cpuregs\[27\]\[13\]
+ _03438_ _03812_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_839 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08436_ _02982_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_1
XFILLER_0_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_850 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08367_ net250 net215 _02251_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07318_ _01964_ _01967_ _01968_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08298_ net222 _02881_ _02757_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07249_ instr_rdcycle is_slli_srli_srai _01825_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_780 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10260_ _04604_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10191_ net1001 _03202_ _04564_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13950_ _01592_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__clkbuf_1
X_12901_ mem_rdata_q\[2\] VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__inv_2
X_13881_ _01555_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15620_ clknet_leaf_38_clk _01195_ VGND VGND VPWR VPWR cpuregs\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12832_ mem_rdata_q\[12\] net4 _03017_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_633 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ clknet_leaf_52_clk _01126_ VGND VGND VPWR VPWR cpuregs\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12763_ _06501_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14502_ clknet_leaf_129_clk _00160_ VGND VGND VPWR VPWR cpuregs\[30\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11714_ _05259_ _05569_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15482_ clknet_leaf_83_clk _01067_ VGND VGND VPWR VPWR mem_rdata_q\[5\] sky130_fd_sc_hd__dfxtp_1
X_12694_ _05900_ _06426_ _06435_ _01918_ decoded_imm\[28\] VGND VGND VPWR VPWR _06436_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14433_ clknet_leaf_96_clk _00091_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_127_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11645_ _05503_ _05242_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_154_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14364_ _01809_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__clkbuf_1
Xinput15 net425 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
X_11576_ _05289_ _05456_ _05458_ _05368_ _05184_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__a221o_1
Xinput26 net1373 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XFILLER_0_13_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13315_ _06811_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10527_ net1387 _03179_ _04746_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__mux2_1
X_14295_ net540 VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__clkbuf_1
X_13246_ _06763_ decoded_imm_j\[3\] _06732_ mem_rdata_q\[10\] _06540_ VGND VGND VPWR
+ VPWR _06774_ sky130_fd_sc_hd__a221o_1
X_10458_ net1383 _03179_ _04709_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10389_ _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__clkbuf_8
X_13177_ _06627_ _06732_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__or2_2
X_12128_ _05889_ _05891_ _05892_ _03090_ _05879_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__o221a_1
X_12059_ _03047_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__clkbuf_8
X_15818_ clknet_leaf_55_clk _01390_ VGND VGND VPWR VPWR cpuregs\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15749_ clknet_leaf_35_clk _01324_ VGND VGND VPWR VPWR cpuregs\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09270_ _03737_ _03706_ _03703_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_118_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08221_ _02818_ _02819_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_820 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08152_ _02752_ _02754_ _02755_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__or3_2
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08083_ _02573_ net248 _02678_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_9_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_641 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08985_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__buf_6
XFILLER_0_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07936_ instr_bge _02555_ instr_bgeu VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__o21bai_1
X_07867_ _02483_ _02486_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__nand2_1
X_09606_ _03647_ _04063_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_79_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07798_ net179 net211 VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__or2_1
X_09537_ cpuregs\[20\]\[15\] cpuregs\[21\]\[15\] cpuregs\[22\]\[15\] cpuregs\[23\]\[15\]
+ _03594_ _03595_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_78_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09468_ _03928_ _03929_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_716 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_19_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08419_ _01816_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_628 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09399_ decoded_imm\[11\] net173 VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11430_ _05313_ _05316_ _05314_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11361_ _05231_ reg_pc\[31\] VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10312_ _04631_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13100_ _06692_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__clkbuf_1
X_14080_ _01661_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__clkbuf_1
X_11292_ _01871_ _05212_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_95_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13031_ cpuregs\[1\]\[15\] _04850_ _06647_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__mux2_1
X_10243_ net1162 _03367_ _04586_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__mux2_1
X_10174_ _04557_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__clkbuf_1
X_14982_ clknet_leaf_103_clk _00640_ VGND VGND VPWR VPWR reg_pc\[28\] sky130_fd_sc_hd__dfxtp_2
X_13933_ _01583_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_161_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13864_ _01546_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15603_ clknet_leaf_145_clk _01178_ VGND VGND VPWR VPWR cpuregs\[31\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12815_ _06536_ _06533_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__nand2_1
X_13795_ net645 _06956_ _07075_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ clknet_leaf_124_clk _01119_ VGND VGND VPWR VPWR cpuregs\[24\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12746_ _06483_ _06484_ _03082_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15465_ clknet_leaf_125_clk _01055_ VGND VGND VPWR VPWR cpuregs\[19\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12677_ cpuregs\[4\]\[28\] cpuregs\[5\]\[28\] cpuregs\[6\]\[28\] cpuregs\[7\]\[28\]
+ _05908_ _06156_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14416_ clknet_leaf_62_clk _00074_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_142_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11628_ _05418_ net600 _05343_ _05506_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15396_ clknet_leaf_94_clk _00986_ VGND VGND VPWR VPWR decoded_imm\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14347_ net693 _03313_ _01800_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11559_ _05393_ _05410_ _05421_ _05434_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__and4_1
Xhold607 cpuregs\[25\]\[17\] VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 cpuregs\[28\]\[20\] VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold629 cpuregs\[18\]\[26\] VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ _01764_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_571 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_122_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_772 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13229_ decoded_imm\[11\] _06752_ _06762_ _06764_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _03264_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_146_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07721_ net487 _02051_ _02345_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__a21oi_1
X_07652_ count_cycle\[22\] _02051_ _02281_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07583_ reg_pc\[18\] decoded_imm\[18\] VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09322_ _03403_ _03788_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09253_ _03575_ _03715_ _03718_ _03721_ _03430_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08204_ net181 _02793_ _02784_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09184_ _03609_ _03610_ _03611_ _03654_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_105_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08135_ _02177_ net209 _02598_ _02641_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__a31o_1
XFILLER_0_161_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08066_ _02099_ _02482_ _02675_ _02676_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_413 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ _03442_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__buf_8
X_07919_ _02200_ net247 VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__nand2_1
X_08899_ reg_pc\[30\] _03371_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__or2_1
X_10930_ _04975_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10861_ cpuregs\[25\]\[14\] _04848_ _04934_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_625 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12600_ _06132_ _06336_ _06345_ _06153_ decoded_imm\[24\] VGND VGND VPWR VPWR _06346_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13580_ _03294_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10792_ _04902_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__clkbuf_1
X_12531_ _06273_ _06275_ _06277_ _06279_ _06151_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15250_ clknet_leaf_76_clk _00843_ VGND VGND VPWR VPWR instr_xor sky130_fd_sc_hd__dfxtp_1
X_12462_ _05974_ cpuregs\[30\]\[18\] _05896_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14201_ _01725_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11413_ _01889_ _05306_ _05308_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15181_ clknet_leaf_81_clk _00806_ VGND VGND VPWR VPWR latched_store sky130_fd_sc_hd__dfxtp_2
XFILLER_0_152_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12393_ _06026_ _06147_ _03081_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_823 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14132_ cpuregs\[7\]\[13\] _06952_ _01685_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__mux2_1
X_11344_ _05031_ _05249_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_878 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14063_ _01652_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__clkbuf_1
X_11275_ reg_next_pc\[6\] _03217_ _02946_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__mux2_2
X_13014_ cpuregs\[1\]\[7\] _04833_ _06636_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10226_ _04563_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__buf_4
X_10157_ net789 _03314_ _04548_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10088_ net1232 _03322_ _04509_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__mux2_1
X_14965_ clknet_leaf_87_clk _00623_ VGND VGND VPWR VPWR reg_pc\[11\] sky130_fd_sc_hd__dfxtp_2
X_13916_ _01574_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__clkbuf_1
X_14896_ clknet_leaf_112_clk net463 VGND VGND VPWR VPWR count_instr\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13847_ _07108_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_84_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13778_ cpuregs\[3\]\[7\] _06939_ _07064_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15517_ clknet_leaf_55_clk _01102_ VGND VGND VPWR VPWR cpuregs\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12729_ _05969_ _06468_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15448_ clknet_leaf_55_clk _01038_ VGND VGND VPWR VPWR cpuregs\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_213 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15379_ clknet_leaf_89_clk _00969_ VGND VGND VPWR VPWR decoded_imm\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_694 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold404 cpuregs\[3\]\[1\] VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold415 cpuregs\[15\]\[18\] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold426 cpuregs\[30\]\[30\] VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold437 net170 VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 cpuregs\[1\]\[4\] VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ _04384_ _04385_ _04386_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__a21oi_1
Xhold459 cpuregs\[12\]\[8\] VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09871_ cpuregs\[28\]\[25\] cpuregs\[29\]\[25\] cpuregs\[30\]\[25\] cpuregs\[31\]\[25\]
+ _03586_ _03449_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_799 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ reg_out\[20\] alu_out_q\[20\] _03175_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__mux2_1
X_08753_ net790 _03248_ _03249_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07704_ _02327_ _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__xor2_1
X_08684_ net975 _03189_ _03185_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__mux2_1
X_07635_ net14 _02202_ _02179_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_156_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07566_ _01932_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09305_ _02099_ _03770_ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_24_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07497_ _02134_ _02136_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09236_ decoded_imm\[5\] net198 VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_376 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_145_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_398 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_17_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_50_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09167_ cpuregs\[24\]\[4\] cpuregs\[25\]\[4\] cpuregs\[26\]\[4\] cpuregs\[27\]\[4\]
+ _03636_ _03637_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_834 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08118_ _02154_ _02471_ _02561_ _02563_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09098_ _01953_ _03545_ _03546_ _03476_ _03570_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08049_ net201 _02659_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__or2_1
Xhold960 cpuregs\[19\]\[12\] VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 cpuregs\[27\]\[18\] VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_777 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold982 cpuregs\[28\]\[11\] VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ count_instr\[5\] count_instr\[4\] VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__and2_1
Xhold993 cpuregs\[11\]\[21\] VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__dlygate4sd3_1
X_10011_ _04453_ _04454_ _04455_ _04425_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14750_ clknet_leaf_149_clk _00408_ VGND VGND VPWR VPWR cpuregs\[26\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__clkbuf_4
X_13701_ _07031_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_123_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ _04966_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__clkbuf_1
X_14681_ clknet_leaf_160_clk _00339_ VGND VGND VPWR VPWR cpuregs\[27\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11893_ count_cycle\[53\] _05706_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__or2_1
X_13632_ net643 _06929_ _06992_ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__mux2_1
X_10844_ net909 _04831_ _04923_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13563_ net900 _06948_ _06946_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10775_ _04893_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15302_ clknet_leaf_34_clk _00892_ VGND VGND VPWR VPWR cpuregs\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12514_ _06263_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13494_ _06906_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15233_ clknet_leaf_80_clk _00826_ VGND VGND VPWR VPWR instr_lhu sky130_fd_sc_hd__dfxtp_1
X_12445_ _06132_ _06186_ _06197_ _06153_ decoded_imm\[17\] VGND VGND VPWR VPWR _06198_
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_35_694 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_519 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15164_ clknet_leaf_51_clk _00789_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dfxtp_4
X_12376_ _06131_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14115_ net636 _06935_ _01674_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11327_ _05231_ reg_pc\[21\] VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__or2_1
X_15095_ clknet_leaf_99_clk _07118_ VGND VGND VPWR VPWR reg_out\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14046_ _01643_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11258_ _05188_ reg_pc\[1\] VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10209_ _04577_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__clkbuf_1
X_11189_ net380 _05140_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__nor2_1
X_14948_ clknet_leaf_117_clk _00606_ VGND VGND VPWR VPWR count_instr\[57\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14879_ clknet_leaf_124_clk _00537_ VGND VGND VPWR VPWR cpuregs\[17\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07420_ _01958_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07351_ _01970_ _01990_ _01991_ _01999_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_425 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07282_ _01934_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_4
XFILLER_0_155_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09021_ cpuregs\[22\]\[1\] cpuregs\[23\]\[1\] _03494_ VGND VGND VPWR VPWR _03495_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_26_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold201 cpuregs\[0\]\[30\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 reg_next_pc\[5\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 cpuregs\[11\]\[15\] VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 cpuregs\[22\]\[21\] VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 count_instr\[29\] VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 instr_xor VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold267 cpuregs\[4\]\[5\] VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 count_cycle\[15\] VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _03593_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold289 _00828_ VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ decoded_imm\[25\] net188 VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__nand2_1
X_08805_ _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__clkbuf_4
X_09785_ _02277_ _03624_ _04237_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08736_ _03234_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__buf_2
*XANTENNA_107 decoded_imm\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_118 reg_pc\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_129 net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08667_ latched_stalu VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ net183 VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__buf_4
XFILLER_0_139_939 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ decoded_imm_j\[3\] decoded_imm_j\[2\] decoded_imm_j\[1\] _03057_ VGND VGND
+ VPWR VPWR _03117_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_101_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ _02007_ _02177_ _01955_ _02185_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_285 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10560_ net649 _03287_ _04757_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__mux2_1
X_09219_ _03455_ _03688_ _03420_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10491_ cpuregs\[14\]\[16\] _03287_ _04720_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12230_ cpuregs\[4\]\[9\] cpuregs\[5\]\[9\] cpuregs\[6\]\[9\] cpuregs\[7\]\[9\] _05834_
+ _03097_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12161_ _03063_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_541 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11112_ count_instr\[20\] net478 count_instr\[18\] _05082_ VGND VGND VPWR VPWR _05087_
+ sky130_fd_sc_hd__and4_1
X_12092_ decoded_imm\[1\] _05860_ _01906_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__mux2_1
Xhold790 cpuregs\[20\]\[6\] VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__dlygate4sd3_1
X_15920_ clknet_leaf_142_clk _01492_ VGND VGND VPWR VPWR cpuregs\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11043_ cpu_state\[1\] count_instr\[1\] count_instr\[0\] decoder_trigger VGND VGND
+ VPWR VPWR _05037_ sky130_fd_sc_hd__and4_1
X_15851_ clknet_leaf_32_clk _01423_ VGND VGND VPWR VPWR cpuregs\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_14802_ clknet_leaf_54_clk _00460_ VGND VGND VPWR VPWR cpuregs\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15782_ clknet_leaf_34_clk _01357_ VGND VGND VPWR VPWR cpuregs\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12994_ _01067_ _06629_ _06630_ _06513_ net647 VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14733_ clknet_leaf_37_clk _00391_ VGND VGND VPWR VPWR cpuregs\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11945_ _03473_ _05740_ _05749_ _03526_ reg_pc\[31\] VGND VGND VPWR VPWR _05750_
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_158_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ clknet_leaf_59_clk _00322_ VGND VGND VPWR VPWR cpuregs\[14\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11876_ _05697_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__clkbuf_1
X_13615_ net735 _06983_ _06967_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10827_ _04920_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__clkbuf_1
X_14595_ clknet_leaf_131_clk _00253_ VGND VGND VPWR VPWR cpuregs\[28\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_414 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_520 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13546_ _03220_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__clkbuf_4
X_10758_ _03385_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__buf_2
XFILLER_0_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13477_ _06897_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_136_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10689_ _04836_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15216_ clknet_leaf_72_clk alu_out\[29\] VGND VGND VPWR VPWR alu_out_q\[29\] sky130_fd_sc_hd__dfxtp_1
X_12428_ cpuregs\[12\]\[17\] cpuregs\[13\]\[17\] cpuregs\[14\]\[17\] cpuregs\[15\]\[17\]
+ _05913_ _05994_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15147_ clknet_leaf_73_clk _00773_ VGND VGND VPWR VPWR mem_do_wdata sky130_fd_sc_hd__dfxtp_2
XFILLER_0_140_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_569 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12359_ _05845_ _06112_ _06114_ _03139_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15078_ clknet_leaf_117_clk _00736_ VGND VGND VPWR VPWR count_cycle\[61\] sky130_fd_sc_hd__dfxtp_1
X_14029_ cpuregs\[5\]\[29\] _06985_ _01624_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ _02250_ _03660_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08521_ _03037_ _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__or2_1
X_08452_ _02265_ _02992_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07403_ count_instr\[6\] _01965_ count_cycle\[38\] _02014_ VGND VGND VPWR VPWR _02049_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08383_ latched_branch latched_store VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07334_ _01982_ _01983_ _01955_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__o21a_2
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07265_ is_slli_srli_srai _01920_ _01840_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09004_ _03391_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07196_ net34 _01859_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09906_ cpuregs\[4\]\[26\] cpuregs\[5\]\[26\] cpuregs\[6\]\[26\] cpuregs\[7\]\[26\]
+ _03457_ _03595_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09837_ _03403_ _04287_ _03420_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__o21a_1
X_09768_ _04219_ _04220_ _03413_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _03173_ _03217_ _03218_ _03219_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__a22o_2
X_09699_ decoded_imm\[20\] net183 VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__or2_1
X_11730_ net431 net435 _05597_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__a21oi_1
X_11661_ _01890_ _05528_ _05536_ _05368_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13400_ cpuregs\[24\]\[4\] _04827_ _06852_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__mux2_1
X_10612_ _04791_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14380_ clknet_leaf_33_clk _00043_ VGND VGND VPWR VPWR cpuregs\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11592_ decoded_imm_j\[20\] _05235_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13331_ _06820_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10543_ net1209 _03235_ _04746_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13262_ cpuregs\[18\]\[3\] _04825_ _06780_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__mux2_1
X_10474_ net1037 _03235_ _04709_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_20_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15001_ clknet_leaf_106_clk _00659_ VGND VGND VPWR VPWR reg_next_pc\[16\] sky130_fd_sc_hd__dfxtp_1
X_12213_ _05974_ cpuregs\[30\]\[8\] _05896_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__o21a_1
X_13193_ mem_rdata_q\[27\] _06742_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_121_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12144_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_131_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12075_ _03061_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__nor2_1
X_11026_ net1038 _04877_ _05017_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__mux2_1
X_15903_ clknet_leaf_101_clk _01475_ VGND VGND VPWR VPWR cpuregs\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15834_ clknet_leaf_135_clk _01406_ VGND VGND VPWR VPWR cpuregs\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15765_ clknet_leaf_141_clk _01340_ VGND VGND VPWR VPWR cpuregs\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_12977_ _06623_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_634 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_151_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14716_ clknet_leaf_14_clk _00374_ VGND VGND VPWR VPWR cpuregs\[15\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11928_ cpuregs\[4\]\[31\] cpuregs\[5\]\[31\] cpuregs\[6\]\[31\] cpuregs\[7\]\[31\]
+ _03439_ _03576_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_522 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15696_ clknet_leaf_6_clk _01271_ VGND VGND VPWR VPWR cpuregs\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14647_ clknet_leaf_13_clk _00305_ VGND VGND VPWR VPWR cpuregs\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11859_ count_cycle\[40\] count_cycle\[41\] count_cycle\[42\] _05680_ VGND VGND VPWR
+ VPWR _05686_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
*XANTENNA_18 _03095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_29 _03170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ clknet_leaf_55_clk _00236_ VGND VGND VPWR VPWR cpuregs\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13529_ net1358 _06923_ _06925_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_923 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_794 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput103 net103 VGND VGND VPWR VPWR mem_la_wdata[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput114 net114 VGND VGND VPWR VPWR mem_la_wdata[25] sky130_fd_sc_hd__clkbuf_4
Xoutput125 net125 VGND VGND VPWR VPWR mem_la_wdata[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput136 net136 VGND VGND VPWR VPWR mem_wdata[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput147 net147 VGND VGND VPWR VPWR mem_wdata[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput158 net158 VGND VGND VPWR VPWR mem_wdata[30] sky130_fd_sc_hd__clkbuf_4
Xoutput169 net169 VGND VGND VPWR VPWR mem_wstrb[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07952_ net448 _02558_ _02565_ _02571_ VGND VGND VPWR VPWR alu_out\[0\] sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_149_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07883_ net108 VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__clkbuf_4
X_09622_ _03959_ _04079_ _03670_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__o21ai_1
X_09553_ _03962_ _03967_ _04012_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__a21oi_1
X_08504_ _03028_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_19_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09484_ _03446_ _03945_ _03417_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08435_ _02200_ _02981_ _02971_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08366_ _02939_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_1
XFILLER_0_74_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07317_ _01954_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08297_ _02433_ _02880_ _02889_ VGND VGND VPWR VPWR alu_out\[27\] sky130_fd_sc_hd__a21o_1
XFILLER_0_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07248_ is_jalr_addi_slti_sltiu_xori_ori_andi is_lui_auipc_jal VGND VGND VPWR VPWR
+ _01906_ sky130_fd_sc_hd__nor2_4
XFILLER_0_21_409 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07179_ _01844_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__clkbuf_4
X_10190_ _04567_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12900_ _02054_ _06553_ net1415 net239 VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__a22o_1
X_13880_ net898 _06973_ _01551_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12831_ _06546_ _06542_ _06548_ _06530_ net469 VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15550_ clknet_leaf_81_clk _00023_ VGND VGND VPWR VPWR cpu_state\[6\] sky130_fd_sc_hd__dfxtp_4
X_12762_ net227 _06500_ _05862_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ clknet_leaf_144_clk _00159_ VGND VGND VPWR VPWR cpuregs\[30\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11713_ _05259_ _05569_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15481_ clknet_leaf_83_clk _01066_ VGND VGND VPWR VPWR mem_rdata_q\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12693_ _06428_ _06430_ _06432_ _06434_ _06151_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__a221o_2
XFILLER_0_37_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14432_ clknet_leaf_96_clk _00090_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dfxtp_4
X_11644_ _05517_ _05511_ _05519_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14363_ net878 _03366_ _01800_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__mux2_1
Xinput16 mem_rdata[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_4
X_11575_ _05032_ _05457_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__nand2_1
Xinput27 mem_rdata[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_133_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13314_ net1369 _04877_ _06802_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10526_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__clkbuf_8
X_14294_ _01772_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13245_ mem_rdata_q\[23\] _06627_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10457_ _04708_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__buf_6
XFILLER_0_110_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13176_ is_beq_bne_blt_bge_bltu_bgeu is_sb_sh_sw VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__or2_2
X_10388_ _04562_ _04671_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__nor2_4
X_12127_ cpuregs\[0\]\[5\] cpuregs\[1\]\[5\] cpuregs\[2\]\[5\] cpuregs\[3\]\[5\] _03096_
+ _03098_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__mux4_1
X_12058_ _03061_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__or2_1
X_11009_ _04994_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15817_ clknet_leaf_34_clk _01389_ VGND VGND VPWR VPWR cpuregs\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ clknet_leaf_41_clk _01323_ VGND VGND VPWR VPWR cpuregs\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15679_ clknet_leaf_48_clk _01254_ VGND VGND VPWR VPWR cpuregs\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08220_ _02801_ _02808_ _02799_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08151_ _02710_ _02753_ _02750_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_60_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_180 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08082_ _02484_ _02581_ _02690_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_628 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08984_ _03407_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07935_ instr_bne is_slti_blt_slt is_sltiu_bltu_sltu net238 VGND VGND VPWR VPWR _02555_
+ sky130_fd_sc_hd__or4b_1
X_07866_ _02484_ _02485_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__nand2_1
X_09605_ cpuregs\[12\]\[17\] cpuregs\[13\]\[17\] cpuregs\[14\]\[17\] cpuregs\[15\]\[17\]
+ _03516_ _03409_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07797_ net179 net211 VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09536_ _03575_ _03991_ _03993_ _03995_ _03591_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__a221o_2
XFILLER_0_78_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09467_ decoded_imm\[13\] net175 VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_503 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08418_ reg_next_pc\[11\] reg_out\[11\] _02969_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__mux2_2
XFILLER_0_53_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09398_ _03862_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08349_ _01880_ net251 net205 _01913_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_394 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11360_ reg_next_pc\[31\] _03383_ _02948_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__mux2_2
X_10311_ net660 _03367_ _04622_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11291_ reg_next_pc\[11\] _03251_ _02946_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_95_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13030_ _06652_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10242_ _04594_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_784 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10173_ net751 _03367_ _04548_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14981_ clknet_leaf_103_clk _00639_ VGND VGND VPWR VPWR reg_pc\[27\] sky130_fd_sc_hd__dfxtp_2
X_13932_ cpuregs\[4\]\[15\] _06956_ _01577_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13863_ cpuregs\[22\]\[15\] _06956_ _07111_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15602_ clknet_leaf_3_clk _01177_ VGND VGND VPWR VPWR cpuregs\[31\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12814_ mem_rdata_q\[13\] VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13794_ _07080_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_913 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_96_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15533_ clknet_leaf_126_clk _01118_ VGND VGND VPWR VPWR cpuregs\[24\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12745_ cpuregs\[0\]\[31\] cpuregs\[1\]\[31\] cpuregs\[2\]\[31\] cpuregs\[3\]\[31\]
+ _03091_ _05829_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15464_ clknet_leaf_126_clk _01054_ VGND VGND VPWR VPWR cpuregs\[19\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12676_ _06418_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_65_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14415_ clknet_leaf_62_clk _00073_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11627_ _05285_ _05241_ _05505_ _05300_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15395_ clknet_leaf_94_clk _00985_ VGND VGND VPWR VPWR decoded_imm\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_108_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_439 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14346_ _01777_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__buf_4
XFILLER_0_142_539 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11558_ _05435_ _05423_ _05432_ _05433_ _05441_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__o311a_1
XFILLER_0_13_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold608 cpuregs\[27\]\[11\] VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10509_ _04736_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14277_ net700 VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__clkbuf_1
Xhold619 cpuregs\[13\]\[10\] VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11489_ _05378_ _05307_ _05206_ _05201_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_150_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13228_ is_beq_bne_blt_bge_bltu_bgeu net445 decoded_imm_j\[11\] _06763_ _06541_ VGND
+ VGND VPWR VPWR _06764_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13159_ net133 _05764_ _06721_ _06673_ net796 VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07720_ count_instr\[59\] _02013_ _02017_ _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_69_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07651_ count_instr\[54\] _02013_ _02017_ _02280_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07582_ _02019_ _02207_ _02216_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09321_ cpuregs\[28\]\[8\] cpuregs\[29\]\[8\] cpuregs\[30\]\[8\] cpuregs\[31\]\[8\]
+ _03641_ _03497_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09252_ _03447_ _03720_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08203_ _02764_ _02774_ _02802_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__nor3_1
X_09183_ _03652_ _03653_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_78_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08134_ _02608_ _02735_ _02736_ _02739_ VGND VGND VPWR VPWR alu_out\[14\] sky130_fd_sc_hd__a31o_1
XFILLER_0_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_695 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_241 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08065_ _02099_ _02482_ _02561_ _02595_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpicorv32_350 VGND VGND VPWR VPWR picorv32_350/HI trace_data[27] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_73_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_90_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07918_ _02200_ net247 VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__or2_1
X_08898_ _03375_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07849_ _02177_ net209 VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10860_ _04938_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09519_ cpuregs\[8\]\[14\] cpuregs\[9\]\[14\] cpuregs\[10\]\[14\] cpuregs\[11\]\[14\]
+ _03601_ _03583_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10791_ net1036 _04846_ _04898_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _06073_ _06278_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_938 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_136_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12461_ cpuregs\[31\]\[18\] _03092_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__or2b_1
XFILLER_0_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14200_ net757 _06952_ _01721_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11412_ _01889_ _05307_ _05273_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__a21oi_1
X_15180_ clknet_leaf_67_clk _00805_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dfxtp_2
X_12392_ cpuregs\[28\]\[15\] cpuregs\[29\]\[15\] cpuregs\[30\]\[15\] cpuregs\[31\]\[15\]
+ _05895_ _05929_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__mux4_1
X_14131_ _01688_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__clkbuf_1
X_11343_ reg_next_pc\[26\] _02999_ _05248_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14062_ net942 _06950_ _01649_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__mux2_1
X_11274_ _05186_ _05199_ _05200_ _01885_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13013_ _06643_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__clkbuf_1
X_10225_ _04585_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ _04525_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_7_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10087_ _04510_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__clkbuf_1
X_14964_ clknet_leaf_88_clk _00622_ VGND VGND VPWR VPWR reg_pc\[10\] sky130_fd_sc_hd__dfxtp_2
X_13915_ cpuregs\[4\]\[7\] _06939_ _01566_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__mux2_1
X_14895_ clknet_leaf_112_clk _00553_ VGND VGND VPWR VPWR count_instr\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13846_ cpuregs\[22\]\[7\] _06939_ _07100_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_581 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13777_ _07071_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__clkbuf_1
X_10989_ cpuregs\[17\]\[10\] _04839_ _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15516_ clknet_leaf_37_clk _01101_ VGND VGND VPWR VPWR cpuregs\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12728_ cpuregs\[24\]\[30\] cpuregs\[25\]\[30\] cpuregs\[26\]\[30\] cpuregs\[27\]\[30\]
+ _03107_ _03108_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12659_ _03124_ _06399_ _06401_ _03139_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__o211a_1
X_15447_ clknet_leaf_37_clk _01037_ VGND VGND VPWR VPWR cpuregs\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15378_ clknet_leaf_89_clk _00968_ VGND VGND VPWR VPWR decoded_imm\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14329_ _01791_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__clkbuf_1
Xhold405 cpuregs\[12\]\[23\] VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 cpuregs\[16\]\[18\] VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold427 cpuregs\[15\]\[30\] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 count_cycle\[24\] VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold449 cpuregs\[14\]\[18\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlygate4sd3_1
X_09870_ _03435_ _04319_ _03425_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _03308_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08752_ _03184_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__buf_4
X_07703_ _02304_ _02328_ _02310_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__o21a_1
X_08683_ _03188_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__buf_2
XFILLER_0_136_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07634_ net184 VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07565_ _02184_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09304_ _02066_ _03619_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_24_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07496_ _02105_ _02111_ _02120_ _02135_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09235_ _03702_ _03703_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_506 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09166_ _03583_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__buf_8
XFILLER_0_32_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08117_ _02154_ _02471_ _02593_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09097_ _03473_ _03560_ _03569_ _03526_ _01971_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08048_ net201 _02659_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold950 cpuregs\[28\]\[7\] VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 cpuregs\[6\]\[8\] VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 cpuregs\[9\]\[7\] VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 cpuregs\[23\]\[13\] VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 cpuregs\[28\]\[10\] VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ _04424_ _04426_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__nor2_1
X_09999_ _04438_ _04440_ _04442_ _04444_ _03429_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11961_ _05763_ _05764_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10912_ net1149 _04831_ _04959_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__mux2_1
X_13700_ net704 _06929_ _07028_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ clknet_leaf_153_clk _00338_ VGND VGND VPWR VPWR cpuregs\[27\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11892_ _05708_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__clkbuf_1
X_13631_ _06994_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__clkbuf_1
X_10843_ _04929_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__clkbuf_1
X_13562_ _03254_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10774_ net868 _04829_ _04887_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12513_ net215 _06262_ _06052_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__mux2_1
X_15301_ clknet_leaf_41_clk _00891_ VGND VGND VPWR VPWR cpuregs\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13493_ net1176 _04852_ _06899_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_160_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_160_clk sky130_fd_sc_hd__clkbuf_2
X_12444_ _06188_ _06190_ _06194_ _06196_ _06151_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__a221o_2
X_15232_ clknet_leaf_76_clk _00825_ VGND VGND VPWR VPWR instr_lbu sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15163_ clknet_leaf_50_clk _00788_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dfxtp_2
X_12375_ _02466_ _06130_ _06052_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14114_ _01679_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__clkbuf_1
X_11326_ reg_next_pc\[21\] _03317_ _02947_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__mux2_2
X_15094_ clknet_leaf_89_clk _07117_ VGND VGND VPWR VPWR reg_out\[12\] sky130_fd_sc_hd__dfxtp_1
X_14045_ net576 _06933_ _01638_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__mux2_1
X_11257_ _01891_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__buf_2
XFILLER_0_66_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10208_ net718 _03255_ _04575_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__mux2_1
X_11188_ net572 _05137_ _05133_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__o21ai_1
X_10139_ _04539_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14947_ clknet_leaf_119_clk _00605_ VGND VGND VPWR VPWR count_instr\[56\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14878_ clknet_leaf_148_clk _00536_ VGND VGND VPWR VPWR cpuregs\[17\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_13829_ _07098_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07350_ _01977_ _01992_ _01995_ _01928_ _01998_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07281_ _01930_ _01931_ _01933_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_151_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_151_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09020_ _03405_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__buf_6
XFILLER_0_143_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold202 count_cycle\[16\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 count_instr\[43\] VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold224 cpuregs\[1\]\[0\] VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 cpuregs\[0\]\[13\] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 cpuregs\[0\]\[4\] VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 cpuregs\[0\]\[7\] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 cpuregs\[29\]\[7\] VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ cpuregs\[20\]\[27\] cpuregs\[21\]\[27\] cpuregs\[22\]\[27\] cpuregs\[23\]\[27\]
+ _03594_ _03442_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__mux4_1
Xhold279 cpuregs\[8\]\[26\] VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09853_ _02306_ _03624_ _04303_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_70_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _03289_ _03292_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__mux2_4
X_09784_ _03672_ _04218_ _04236_ _03665_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__o211a_1
X_08735_ _03173_ _03230_ _03231_ _03233_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__a22o_2
*XANTENNA_108 decoded_imm\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08666_ _03172_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__clkbuf_4
*XANTENNA_119 reg_pc\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07617_ _02247_ _02248_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _03090_ _03112_ _03115_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07548_ _02180_ _02181_ _02184_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_101_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_142_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_142_clk sky130_fd_sc_hd__clkbuf_2
X_07479_ reg_pc\[11\] decoded_imm\[11\] VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09218_ cpuregs\[28\]\[5\] cpuregs\[29\]\[5\] cpuregs\[30\]\[5\] cpuregs\[31\]\[5\]
+ _03641_ _03642_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10490_ _04726_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09149_ _03616_ _03618_ _03620_ _01942_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12160_ _03143_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_15_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_553 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11111_ _05085_ _05086_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__nor2_1
X_12091_ _03080_ _05850_ _05859_ net244 VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold780 cpuregs\[25\]\[7\] VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold791 cpuregs\[13\]\[20\] VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__dlygate4sd3_1
X_11042_ _01820_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__clkbuf_8
X_15850_ clknet_leaf_58_clk _01422_ VGND VGND VPWR VPWR cpuregs\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14801_ clknet_leaf_37_clk _00459_ VGND VGND VPWR VPWR cpuregs\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15781_ clknet_leaf_34_clk _01356_ VGND VGND VPWR VPWR cpuregs\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12993_ is_jalr_addi_slti_sltiu_xori_ori_andi _06626_ _06633_ VGND VGND VPWR VPWR
+ _00882_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_28_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ clknet_leaf_27_clk _00390_ VGND VGND VPWR VPWR cpuregs\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_24_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11944_ _05742_ _05744_ _05746_ _05748_ _03430_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11875_ _05695_ _01842_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__and3b_1
X_14663_ clknet_leaf_136_clk _00321_ VGND VGND VPWR VPWR cpuregs\[14\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13614_ _03366_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__buf_2
X_10826_ net1293 _04881_ _04886_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_940 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14594_ clknet_leaf_130_clk _00252_ VGND VGND VPWR VPWR cpuregs\[28\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10757_ _04882_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__clkbuf_1
X_13545_ _06936_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_133_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_133_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13476_ net843 _04835_ _06888_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__mux2_1
X_10688_ cpuregs\[26\]\[8\] _04835_ _04819_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12427_ _06178_ _06179_ _06014_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__mux2_1
X_15215_ clknet_leaf_71_clk alu_out\[28\] VGND VGND VPWR VPWR alu_out_q\[28\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_33_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12358_ _03042_ _06113_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__or2_1
X_15146_ clknet_leaf_73_clk _00772_ VGND VGND VPWR VPWR mem_do_rdata sky130_fd_sc_hd__dfxtp_2
XFILLER_0_23_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11309_ reg_next_pc\[16\] _03284_ _02947_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__mux2_2
X_15077_ clknet_leaf_117_clk _00735_ VGND VGND VPWR VPWR count_cycle\[60\] sky130_fd_sc_hd__dfxtp_1
X_12289_ cpuregs\[24\]\[11\] cpuregs\[25\]\[11\] cpuregs\[26\]\[11\] cpuregs\[27\]\[11\]
+ _03095_ _05932_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14028_ _01633_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08520_ cpuregs\[20\]\[2\] cpuregs\[21\]\[2\] cpuregs\[22\]\[2\] cpuregs\[23\]\[2\]
+ _03038_ _03039_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08451_ _01816_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07402_ _02007_ _02044_ _02047_ _01927_ _01968_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__a221o_1
X_08382_ net227 _02252_ _02935_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__a21o_2
XFILLER_0_42_50 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07333_ count_instr\[2\] instr_rdinstr count_cycle\[2\] _01950_ VGND VGND VPWR VPWR
+ _01983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_124_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_124_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_144_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07264_ is_sll_srl_sra _01916_ _01919_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09003_ _03397_ _03398_ _03399_ _03477_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07195_ _01820_ _01859_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3 _06564_ VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__buf_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09905_ _03746_ _04353_ _03467_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09836_ cpuregs\[12\]\[24\] cpuregs\[13\]\[24\] cpuregs\[14\]\[24\] cpuregs\[15\]\[24\]
+ _03494_ _03497_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__mux4_1
X_09767_ cpuregs\[20\]\[22\] cpuregs\[21\]\[22\] cpuregs\[22\]\[22\] cpuregs\[23\]\[22\]
+ _03719_ _03450_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ reg_pc\[6\] _03211_ _03172_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__a21oi_1
X_09698_ decoded_imm\[20\] net183 VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__nand2_1
X_08649_ decoded_imm_j\[1\] _01083_ _03022_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11660_ _05534_ _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__nor2_1
X_10611_ net916 _03235_ _04782_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_115_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_115_clk sky130_fd_sc_hd__clkbuf_2
X_11591_ _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13330_ net1356 _04825_ _06816_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10542_ _04754_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_930 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _06783_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__clkbuf_1
X_10473_ _04717_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__clkbuf_1
X_12212_ _05816_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__buf_4
X_15000_ clknet_leaf_107_clk _00658_ VGND VGND VPWR VPWR reg_next_pc\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13192_ decoded_imm\[28\] _06740_ _06737_ _06744_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12143_ _00007_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12074_ cpuregs\[8\]\[1\] cpuregs\[9\]\[1\] cpuregs\[10\]\[1\] cpuregs\[11\]\[1\]
+ _05819_ _03086_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__mux4_1
X_11025_ _05025_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__clkbuf_1
X_15902_ clknet_leaf_135_clk _01474_ VGND VGND VPWR VPWR cpuregs\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15833_ clknet_leaf_140_clk _01405_ VGND VGND VPWR VPWR cpuregs\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15764_ clknet_leaf_102_clk _01339_ VGND VGND VPWR VPWR cpuregs\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12976_ decoded_imm_j\[1\] _01083_ _03021_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__mux2_1
X_14715_ clknet_leaf_9_clk _00373_ VGND VGND VPWR VPWR cpuregs\[15\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11927_ net459 _05730_ _05732_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15695_ clknet_leaf_6_clk _01270_ VGND VGND VPWR VPWR cpuregs\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14646_ clknet_leaf_12_clk _00304_ VGND VGND VPWR VPWR cpuregs\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11858_ _05685_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_329 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10809_ _04911_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_106_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_106_clk sky130_fd_sc_hd__clkbuf_2
*XANTENNA_19 _03106_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_768 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11789_ count_cycle\[19\] _05634_ count_cycle\[20\] VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__a21o_1
X_14577_ clknet_leaf_36_clk _00235_ VGND VGND VPWR VPWR cpuregs\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13528_ _06924_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13459_ _06887_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_935 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput104 net104 VGND VGND VPWR VPWR mem_la_wdata[16] sky130_fd_sc_hd__buf_2
XFILLER_0_11_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput115 net115 VGND VGND VPWR VPWR mem_la_wdata[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput126 net126 VGND VGND VPWR VPWR mem_la_wdata[7] sky130_fd_sc_hd__clkbuf_4
Xoutput137 net137 VGND VGND VPWR VPWR mem_wdata[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput148 net148 VGND VGND VPWR VPWR mem_wdata[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_389 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15129_ clknet_leaf_71_clk _00755_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfxtp_1
Xoutput159 net159 VGND VGND VPWR VPWR mem_wdata[31] sky130_fd_sc_hd__clkbuf_4
X_07951_ _02508_ _02566_ _02569_ net1416 VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_149_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_50_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07882_ net251 VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__inv_2
X_09621_ _02265_ _03770_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09552_ _04010_ _04011_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__nand2_1
X_08503_ mem_rdata_q\[18\] net10 _03018_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__mux2_1
X_09483_ cpuregs\[28\]\[13\] cpuregs\[29\]\[13\] cpuregs\[30\]\[13\] cpuregs\[31\]\[13\]
+ _03586_ _03441_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08434_ reg_next_pc\[16\] reg_out\[16\] _02969_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_82_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_770 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08365_ net251 net213 _02251_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07316_ count_instr\[1\] _01965_ count_cycle\[1\] _01951_ _01966_ VGND VGND VPWR
+ VPWR _01967_ sky130_fd_sc_hd__a221o_2
XFILLER_0_74_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08296_ _02885_ _02886_ _02887_ _02888_ _02584_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__o311a_1
XFILLER_0_46_598 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_132_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07247_ _01839_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_456 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07178_ net182 VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_113_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09819_ _02316_ _03619_ _04269_ _03616_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__a211o_1
X_12830_ _06532_ mem_rdata_q\[13\] _06533_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12761_ _05900_ _06490_ _06499_ _01918_ decoded_imm\[31\] VGND VGND VPWR VPWR _06500_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_139_512 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ clknet_leaf_144_clk _00158_ VGND VGND VPWR VPWR cpuregs\[30\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11712_ _05579_ _05582_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__xor2_1
X_12692_ _03106_ _06433_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__or2_1
X_15480_ clknet_leaf_83_clk _01065_ VGND VGND VPWR VPWR mem_rdata_q\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11643_ _05517_ _05511_ _05519_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__nand3_1
XFILLER_0_65_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14431_ clknet_leaf_97_clk _00089_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_543 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14362_ _01808_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__clkbuf_1
X_11574_ _05230_ _05448_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__and2_1
Xinput17 mem_rdata[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_4
Xinput28 mem_rdata[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_133_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _06810_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__clkbuf_1
X_10525_ _03183_ _04744_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_133_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14293_ net668 VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13244_ decoded_imm\[4\] _06531_ _06771_ _06772_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__o22a_1
X_10456_ _04481_ _04524_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13175_ _01944_ _06730_ _06731_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__o21a_1
X_10387_ latched_rd\[3\] latched_rd\[4\] latched_rd\[2\] VGND VGND VPWR VPWR _04671_
+ sky130_fd_sc_hd__nand3b_4
X_12126_ _03098_ _05890_ _03083_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__a21o_1
X_12057_ cpuregs\[16\]\[0\] cpuregs\[17\]\[0\] cpuregs\[18\]\[0\] cpuregs\[19\]\[0\]
+ _05819_ _03086_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__mux4_1
X_11008_ _05016_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
X_15816_ clknet_leaf_34_clk _01388_ VGND VGND VPWR VPWR cpuregs\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15747_ clknet_leaf_46_clk _01322_ VGND VGND VPWR VPWR cpuregs\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12959_ _06614_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_47_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15678_ clknet_leaf_17_clk _01253_ VGND VGND VPWR VPWR cpuregs\[29\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14629_ clknet_leaf_153_clk _00287_ VGND VGND VPWR VPWR cpuregs\[21\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08150_ _02709_ _02753_ _02750_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_513 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_56_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08081_ _02125_ net205 _02598_ _02563_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08983_ _03457_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__buf_6
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07934_ _02544_ _02549_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__nor2_1
X_07865_ _02125_ net205 VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ _03437_ _04061_ _03419_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07796_ net211 VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__inv_2
X_09535_ _03447_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_318 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09466_ decoded_imm\[13\] net175 VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_35_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08417_ _02948_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09397_ _02112_ _03861_ _03395_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__mux2_1
X_08348_ net248 _02927_ _02930_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__a21o_1
XFILLER_0_62_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08279_ _02316_ _02863_ _02872_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__o21ai_1
X_10310_ _04630_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11290_ _05186_ _05210_ _05211_ _01885_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_95_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10241_ net1216 _03360_ _04586_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__mux2_1
X_10172_ _04556_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14980_ clknet_leaf_109_clk _00638_ VGND VGND VPWR VPWR reg_pc\[26\] sky130_fd_sc_hd__dfxtp_2
X_13931_ _01582_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_161_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13862_ _01545_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15601_ clknet_leaf_154_clk _01176_ VGND VGND VPWR VPWR cpuregs\[31\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12813_ net470 _06530_ _06535_ _05804_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13793_ net1282 _06954_ _07075_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ clknet_leaf_148_clk _01117_ VGND VGND VPWR VPWR cpuregs\[24\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12744_ cpuregs\[4\]\[31\] cpuregs\[5\]\[31\] cpuregs\[6\]\[31\] cpuregs\[7\]\[31\]
+ _05908_ _05909_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15463_ clknet_leaf_148_clk _01053_ VGND VGND VPWR VPWR cpuregs\[19\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12675_ net222 _06417_ _06282_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_800 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14414_ clknet_4_12_0_clk _00072_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_154_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11626_ _05500_ _05501_ _05504_ _01889_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__a22o_1
X_15394_ clknet_leaf_94_clk _00984_ VGND VGND VPWR VPWR decoded_imm\[14\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_42_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_389 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_343 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14345_ _01799_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11557_ _05420_ _05432_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__or2_1
X_10508_ cpuregs\[14\]\[24\] _03341_ _04731_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__mux2_1
Xhold609 cpuregs\[17\]\[0\] VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__dlygate4sd3_1
X_14276_ _01763_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11488_ reg_next_pc\[7\] _02999_ _05203_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10439_ _04699_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__clkbuf_1
X_13227_ _05367_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13158_ net449 _05767_ _06722_ _05763_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__o22a_1
X_12109_ cpuregs\[20\]\[5\] cpuregs\[21\]\[5\] _03096_ VGND VGND VPWR VPWR _05874_
+ sky130_fd_sc_hd__mux2_1
X_13089_ net740 _02503_ _06685_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07650_ count_instr\[22\] _01949_ count_cycle\[54\] _01947_ VGND VGND VPWR VPWR _02280_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07581_ _02058_ _02212_ _02215_ _02071_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09320_ _03415_ _03786_ _03420_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09251_ cpuregs\[28\]\[6\] cpuregs\[29\]\[6\] cpuregs\[30\]\[6\] cpuregs\[31\]\[6\]
+ _03719_ _03450_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08202_ _02784_ _02785_ _02794_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09182_ decoded_imm\[4\] net197 VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_490 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08133_ _02165_ _02466_ _02737_ _02738_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_570 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08064_ _02099_ _02482_ _02593_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_340 VGND VGND VPWR VPWR picorv32_340/HI trace_data[17] sky130_fd_sc_hd__conb_1
Xpicorv32_351 VGND VGND VPWR VPWR picorv32_351/HI trace_data[28] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_90_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ _03407_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_90_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07917_ _02177_ _02462_ _02474_ _02531_ _02536_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__o221a_1
X_08897_ net894 _03374_ _03315_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_95_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_2
X_07848_ _02177_ net209 VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07779_ net216 VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09518_ _03454_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10790_ _04901_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09449_ cpuregs\[24\]\[12\] cpuregs\[25\]\[12\] cpuregs\[26\]\[12\] cpuregs\[27\]\[12\]
+ _03640_ _03496_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12460_ _05969_ _06211_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11411_ _05191_ _05195_ _05197_ _05199_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__nand4_1
X_12391_ _06023_ _06145_ _05927_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_151_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_592 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14130_ net926 _06950_ _01685_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__mux2_1
X_11342_ _02948_ _03350_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14061_ _01651_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__clkbuf_1
X_11273_ _05188_ reg_pc\[5\] VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10224_ net928 _03307_ _04575_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__mux2_1
X_13012_ cpuregs\[1\]\[6\] _04831_ _06636_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__mux2_1
X_10155_ _04547_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10086_ cpuregs\[12\]\[20\] _03314_ _04509_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__mux2_1
X_14963_ clknet_leaf_88_clk _00621_ VGND VGND VPWR VPWR reg_pc\[9\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_86_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_2
X_13914_ _01573_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__clkbuf_1
X_14894_ clknet_leaf_112_clk _00552_ VGND VGND VPWR VPWR count_instr\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13845_ _07107_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_593 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13776_ net1102 _06937_ _07064_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__mux2_1
X_10988_ _04994_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_44_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15515_ clknet_leaf_27_clk _01100_ VGND VGND VPWR VPWR cpuregs\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12727_ _03142_ _06462_ _06466_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_26_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15446_ clknet_leaf_27_clk _01036_ VGND VGND VPWR VPWR cpuregs\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12658_ _03042_ _06400_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11609_ _05487_ _05488_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__or2_1
X_15377_ clknet_leaf_88_clk _00967_ VGND VGND VPWR VPWR decoded_imm\[31\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12589_ _06138_ _06334_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14328_ cpuregs\[10\]\[11\] _03254_ _01789_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__mux2_1
Xhold406 count_instr\[7\] VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold417 cpuregs\[3\]\[13\] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 cpuregs\[12\]\[16\] VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 cpuregs\[31\]\[16\] VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14259_ net568 VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_110_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ net905 _03307_ _03249_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _03247_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_77_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_2
X_07702_ _02302_ _02311_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__or2b_1
XFILLER_0_136_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08682_ reg_pc\[1\] _03187_ _03172_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__mux2_2
XFILLER_0_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07633_ _02262_ _02263_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_914 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07564_ net178 VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09303_ net243 VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_608 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_76_777 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07495_ reg_pc\[11\] decoded_imm\[11\] VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09234_ decoded_imm\[6\] net199 VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_693 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_145_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_518 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09165_ _03582_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__buf_8
XFILLER_0_32_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_674 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_90_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08116_ _02720_ _02721_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09096_ _03562_ _03564_ _03566_ _03568_ _03430_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08047_ _02476_ _02658_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_793 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold940 cpuregs\[14\]\[21\] VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold951 cpuregs\[15\]\[20\] VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_880 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold962 cpuregs\[3\]\[22\] VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 cpuregs\[11\]\[4\] VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 cpuregs\[31\]\[8\] VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 cpuregs\[8\]\[21\] VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__dlygate4sd3_1
X_09998_ _03435_ _04443_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ cpuregs\[0\]\[0\] cpuregs\[1\]\[0\] cpuregs\[2\]\[0\] cpuregs\[3\]\[0\] _03406_
+ _03410_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_68_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11960_ net96 net129 VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_123_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _04965_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_123_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _05706_ _01842_ _05707_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__and3b_1
X_13630_ net641 _06927_ _06992_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10842_ net869 _04829_ _04923_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_744 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13561_ _06947_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__clkbuf_1
X_10773_ _04892_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__clkbuf_1
X_15300_ clknet_leaf_42_clk _00890_ VGND VGND VPWR VPWR cpuregs\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12512_ _06132_ _06252_ _06261_ _06153_ decoded_imm\[20\] VGND VGND VPWR VPWR _06262_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13492_ _06905_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15231_ clknet_leaf_77_clk _00824_ VGND VGND VPWR VPWR instr_lw sky130_fd_sc_hd__dfxtp_1
X_12443_ _06073_ _06195_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_600 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15162_ clknet_leaf_50_clk _00787_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dfxtp_2
X_12374_ _05901_ _06116_ _06129_ _05904_ decoded_imm\[14\] VGND VGND VPWR VPWR _06130_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14113_ net591 _06933_ _01674_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__mux2_1
X_11325_ _05227_ _05235_ _05236_ _05224_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__o211a_1
X_15093_ clknet_leaf_89_clk _07116_ VGND VGND VPWR VPWR reg_out\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_97_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11256_ reg_next_pc\[1\] _03187_ _02946_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__mux2_2
X_14044_ _01642_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_120_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10207_ _04576_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__clkbuf_1
X_11187_ count_instr\[43\] count_instr\[42\] count_instr\[41\] _05132_ VGND VGND VPWR
+ VPWR _05139_ sky130_fd_sc_hd__and4_1
X_10138_ cpuregs\[30\]\[11\] _03255_ _04537_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_59_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_2
X_14946_ clknet_leaf_120_clk _00604_ VGND VGND VPWR VPWR count_instr\[55\] sky130_fd_sc_hd__dfxtp_1
X_10069_ net1306 _03263_ _04498_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14877_ clknet_leaf_157_clk _00535_ VGND VGND VPWR VPWR cpuregs\[17\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13828_ net1160 _06989_ _07063_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_307 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13759_ _07061_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_632 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_45_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07280_ _01930_ mem_wordsize\[2\] _01932_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__a21o_4
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_490 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_128_687 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15429_ clknet_leaf_125_clk _01019_ VGND VGND VPWR VPWR cpuregs\[18\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold203 count_cycle\[55\] VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold214 cpuregs\[6\]\[3\] VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 cpuregs\[2\]\[15\] VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 count_instr\[34\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold247 cpuregs\[0\]\[1\] VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 cpuregs\[11\]\[20\] VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 cpuregs\[10\]\[23\] VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _03575_ _04364_ _04366_ _04368_ _03489_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09852_ _03672_ _04284_ _04302_ _03665_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_70_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _03199_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__buf_4
X_09783_ reg_pc\[22\] _03528_ _04235_ _03626_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__a211o_1
X_08734_ _03172_ _03232_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__nor2_1
*XANTENNA_109 decoded_imm\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08665_ _03171_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _02246_ _02242_ _02245_ _01893_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_70 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08596_ _03113_ _03114_ _03054_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07547_ _02183_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07478_ reg_pc\[11\] decoded_imm\[11\] VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_91_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09217_ _03455_ _03686_ _03575_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_348 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09148_ _02066_ _03619_ _03074_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09079_ _03400_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__buf_6
XFILLER_0_20_828 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11110_ net478 _05083_ _05044_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12090_ _05852_ _05854_ _05856_ _05858_ _00011_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__o221a_1
Xhold770 cpuregs\[8\]\[12\] VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 cpuregs\[27\]\[4\] VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 cpuregs\[19\]\[18\] VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _05035_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__clkbuf_1
X_14800_ clknet_leaf_29_clk _00458_ VGND VGND VPWR VPWR cpuregs\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15780_ clknet_leaf_38_clk _01355_ VGND VGND VPWR VPWR cpuregs\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12992_ is_alu_reg_imm _06537_ _06553_ instr_jalr VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_28_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ clknet_leaf_45_clk _00389_ VGND VGND VPWR VPWR cpuregs\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11943_ _03436_ _05747_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14662_ clknet_leaf_137_clk _00320_ VGND VGND VPWR VPWR cpuregs\[14\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11874_ count_cycle\[46\] _05692_ count_cycle\[47\] VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_158_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13613_ _06982_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__clkbuf_1
X_10825_ _04919_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14593_ clknet_leaf_145_clk _00251_ VGND VGND VPWR VPWR cpuregs\[28\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_138_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13544_ cpuregs\[31\]\[5\] _06935_ _06925_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__mux2_1
X_10756_ cpuregs\[26\]\[30\] _04881_ _04818_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_70_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13475_ _06896_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__clkbuf_1
X_10687_ _03234_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_136_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15214_ clknet_leaf_101_clk alu_out\[27\] VGND VGND VPWR VPWR alu_out_q\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12426_ cpuregs\[0\]\[17\] cpuregs\[1\]\[17\] cpuregs\[2\]\[17\] cpuregs\[3\]\[17\]
+ _06055_ _05909_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15145_ clknet_leaf_80_clk _00771_ VGND VGND VPWR VPWR mem_do_rinst sky130_fd_sc_hd__dfxtp_2
X_12357_ cpuregs\[8\]\[14\] cpuregs\[9\]\[14\] cpuregs\[10\]\[14\] cpuregs\[11\]\[14\]
+ _05907_ _03047_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11308_ _05186_ _05222_ _05223_ _05224_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15076_ clknet_leaf_118_clk _00734_ VGND VGND VPWR VPWR count_cycle\[59\] sky130_fd_sc_hd__dfxtp_1
X_12288_ _06026_ _06046_ _03081_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__o21a_1
X_14027_ net1159 _06983_ _01624_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__mux2_1
X_11239_ count_instr\[59\] count_instr\[58\] count_instr\[57\] _05168_ VGND VGND VPWR
+ VPWR _05175_ sky130_fd_sc_hd__and4_4
XTAP_TAPCELL_ROW_52_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14929_ clknet_leaf_114_clk _00587_ VGND VGND VPWR VPWR count_instr\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08450_ reg_next_pc\[21\] reg_out\[21\] _02991_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__mux2_1
X_07401_ net29 net130 _02046_ _01940_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08381_ net226 _02252_ _02934_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__a21o_1
XFILLER_0_86_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07332_ count_instr\[34\] _01946_ _01947_ count_cycle\[34\] VGND VGND VPWR VPWR _01982_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_46_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07263_ _01918_ _01908_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09002_ _03432_ _03470_ _03474_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__and4b_1
XFILLER_0_26_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07194_ mem_do_rinst _01855_ _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_476 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_131_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09904_ cpuregs\[8\]\[26\] cpuregs\[9\]\[26\] cpuregs\[10\]\[26\] cpuregs\[11\]\[26\]
+ _03601_ _03583_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09835_ _03415_ _04285_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__or2_1
X_09766_ cpuregs\[16\]\[22\] cpuregs\[17\]\[22\] cpuregs\[18\]\[22\] cpuregs\[19\]\[22\]
+ _03587_ _03588_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08717_ reg_pc\[6\] _03211_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__or2_1
X_09697_ _04149_ _04151_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__and2_1
Xrebuffer40 net400 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08648_ _03162_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__buf_1
XFILLER_0_138_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08579_ _03097_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10610_ _04790_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__clkbuf_1
X_11590_ _05233_ _05235_ _05457_ instr_jal VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_566 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10541_ net1365 _03228_ _04746_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13260_ net1296 _04823_ _06780_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__mux2_1
X_10472_ cpuregs\[14\]\[7\] _03228_ _04709_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12211_ cpuregs\[31\]\[8\] _03092_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13191_ net1210 _06742_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__and2_1
X_12142_ cpuregs\[4\]\[6\] cpuregs\[5\]\[6\] cpuregs\[6\]\[6\] cpuregs\[7\]\[6\] _05834_
+ _03097_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_131_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12073_ _03082_ _05841_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__nor2_1
X_11024_ net925 _04875_ _05017_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__mux2_1
X_15901_ clknet_leaf_20_clk _01473_ VGND VGND VPWR VPWR cpuregs\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_15832_ clknet_leaf_142_clk _01404_ VGND VGND VPWR VPWR cpuregs\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15763_ clknet_leaf_140_clk _01338_ VGND VGND VPWR VPWR cpuregs\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12975_ _06622_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
X_14714_ clknet_leaf_10_clk _00372_ VGND VGND VPWR VPWR cpuregs\[15\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11926_ net459 _05730_ _05036_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__a21oi_1
X_15694_ clknet_leaf_9_clk _01269_ VGND VGND VPWR VPWR cpuregs\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14645_ clknet_leaf_10_clk _00303_ VGND VGND VPWR VPWR cpuregs\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11857_ _05683_ _01842_ _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__and3b_1
XFILLER_0_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10808_ net772 _04863_ _04909_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_12 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14576_ clknet_leaf_33_clk _00234_ VGND VGND VPWR VPWR cpuregs\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11788_ count_cycle\[19\] count_cycle\[20\] _05634_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__and3_1
X_13527_ _03183_ _04522_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__nor2_4
XFILLER_0_126_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10739_ _04870_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13458_ _03180_ _04562_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__nor2_2
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12409_ _06138_ _06162_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__or2_1
Xoutput105 net105 VGND VGND VPWR VPWR mem_la_wdata[17] sky130_fd_sc_hd__clkbuf_4
X_13389_ _06850_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__clkbuf_1
Xoutput116 net116 VGND VGND VPWR VPWR mem_la_wdata[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_625 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput127 net127 VGND VGND VPWR VPWR mem_la_wdata[8] sky130_fd_sc_hd__clkbuf_4
Xoutput138 net138 VGND VGND VPWR VPWR mem_wdata[12] sky130_fd_sc_hd__clkbuf_4
X_15128_ clknet_leaf_72_clk _00754_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
Xoutput149 net149 VGND VGND VPWR VPWR mem_wdata[22] sky130_fd_sc_hd__buf_2
XFILLER_0_11_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15059_ clknet_leaf_113_clk _00717_ VGND VGND VPWR VPWR count_cycle\[42\] sky130_fd_sc_hd__dfxtp_1
X_07950_ is_compare _02562_ _02560_ _02568_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__nor4_1
X_07881_ _02491_ _02495_ _02500_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09620_ _02222_ _03481_ _04077_ _03483_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__a211o_1
X_09551_ decoded_imm\[15\] net177 VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08502_ _03027_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09482_ _03557_ _03943_ _03425_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_19_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08433_ _02980_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_65_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_714 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_736 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_58_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08364_ _02938_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07315_ count_instr\[33\] _01946_ _01947_ count_cycle\[33\] VGND VGND VPWR VPWR _01966_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08295_ _02885_ _02886_ _02887_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07246_ _01904_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07177_ _01842_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09818_ _02290_ _03660_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09749_ _02250_ _03479_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__nor2_1
X_12760_ _06492_ _06494_ _06496_ _06498_ _05978_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11711_ _05580_ _05581_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12691_ cpuregs\[24\]\[28\] cpuregs\[25\]\[28\] cpuregs\[26\]\[28\] cpuregs\[27\]\[28\]
+ _03150_ _03151_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14430_ clknet_leaf_59_clk _00088_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dfxtp_4
X_11642_ _05518_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14361_ net1192 _03359_ _01800_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11573_ _05454_ _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__xor2_1
Xinput18 net415 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
X_13312_ net950 _04875_ _06802_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__mux2_1
Xinput29 mem_rdata[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
X_10524_ latched_rd\[2\] latched_rd\[4\] latched_rd\[3\] VGND VGND VPWR VPWR _04744_
+ sky130_fd_sc_hd__nand3b_4
XFILLER_0_107_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14292_ _01771_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_878 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13243_ _06763_ decoded_imm_j\[4\] _06732_ mem_rdata_q\[11\] _06541_ VGND VGND VPWR
+ VPWR _06772_ sky130_fd_sc_hd__a221o_1
X_10455_ _04707_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13174_ net544 _06726_ _01915_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10386_ _04670_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12125_ cpuregs\[6\]\[5\] cpuregs\[7\]\[5\] _03085_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12056_ _05815_ _05818_ _05821_ _05823_ _05825_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__a32o_1
X_11007_ cpuregs\[17\]\[19\] _04858_ _05006_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15815_ clknet_leaf_39_clk _01387_ VGND VGND VPWR VPWR cpuregs\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15746_ clknet_leaf_40_clk _01321_ VGND VGND VPWR VPWR cpuregs\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12958_ mem_rdata_q\[10\] net2 _03018_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11909_ count_cycle\[55\] count_cycle\[56\] count_cycle\[57\] count_cycle\[58\] VGND
+ VGND VPWR VPWR _05720_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_16_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15677_ clknet_leaf_25_clk _01252_ VGND VGND VPWR VPWR cpuregs\[29\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12889_ _06572_ _06573_ _06574_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__or3_2
XFILLER_0_23_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14628_ clknet_leaf_150_clk _00286_ VGND VGND VPWR VPWR cpuregs\[21\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_56_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_427 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_23_86 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14559_ clknet_leaf_133_clk _00217_ VGND VGND VPWR VPWR cpuregs\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_525 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08080_ _02584_ _02686_ _02687_ _02689_ _02479_ VGND VGND VPWR VPWR alu_out\[10\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08982_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07933_ instr_bne _02552_ net238 VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_48_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07864_ _02125_ net205 VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__nand2_1
X_09603_ cpuregs\[8\]\[17\] cpuregs\[9\]\[17\] cpuregs\[10\]\[17\] cpuregs\[11\]\[17\]
+ _03440_ _03451_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07795_ _02413_ _02414_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__and2_1
X_09534_ cpuregs\[12\]\[15\] cpuregs\[13\]\[15\] cpuregs\[14\]\[15\] cpuregs\[15\]\[15\]
+ _03587_ _03588_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09465_ _02139_ _03624_ _03927_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_35_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08416_ _02968_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
XFILLER_0_148_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09396_ _03488_ _03842_ _03860_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08347_ _01880_ _02509_ net248 _01913_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_558 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08278_ _02306_ _02852_ _02863_ _02316_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07229_ instr_jal VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_15_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10240_ _04593_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_1
X_10171_ cpuregs\[30\]\[27\] _03360_ _04548_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13930_ cpuregs\[4\]\[14\] _06954_ _01577_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__mux2_1
X_13861_ cpuregs\[22\]\[14\] _06954_ _07111_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_161_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15600_ clknet_leaf_2_clk _01175_ VGND VGND VPWR VPWR cpuregs\[31\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_126_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12812_ _06531_ _06534_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13792_ _07079_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__clkbuf_1
X_15531_ clknet_leaf_149_clk _01116_ VGND VGND VPWR VPWR cpuregs\[24\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_12743_ _06482_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15462_ clknet_leaf_149_clk _01052_ VGND VGND VPWR VPWR cpuregs\[19\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12674_ _05900_ _06403_ _06416_ _01918_ decoded_imm\[27\] VGND VGND VPWR VPWR _06417_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_127_538 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14413_ clknet_leaf_64_clk _00071_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_53_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11625_ _05502_ _05503_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15393_ clknet_leaf_99_clk _00983_ VGND VGND VPWR VPWR decoded_imm\[15\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_108_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_519 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14344_ net791 _03306_ _01789_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__mux2_1
X_11556_ _05418_ net543 _05343_ _05440_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_582 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10507_ _04735_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__clkbuf_1
X_14275_ net537 VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__clkbuf_1
X_11487_ _05212_ _05365_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13226_ net1406 _06627_ net446 VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10438_ cpuregs\[21\]\[23\] _03334_ _04695_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13157_ _01822_ net132 _01818_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__o21ba_1
X_10369_ cpuregs\[28\]\[23\] _03334_ _04658_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12108_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__buf_4
X_13088_ _06686_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_146_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12039_ _01860_ _05811_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07580_ _02065_ _02213_ _02201_ _02214_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_904 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15729_ clknet_leaf_154_clk _01304_ VGND VGND VPWR VPWR cpuregs\[22\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09250_ _03548_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__buf_8
XFILLER_0_8_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08201_ _02799_ _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__or2_2
XFILLER_0_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09181_ decoded_imm\[4\] net197 VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08132_ _02165_ _02466_ _02598_ _02563_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_117_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08063_ _02672_ _02673_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_330 VGND VGND VPWR VPWR picorv32_330/HI trace_data[7] sky130_fd_sc_hd__conb_1
Xpicorv32_341 VGND VGND VPWR VPWR picorv32_341/HI trace_data[18] sky130_fd_sc_hd__conb_1
XFILLER_0_3_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_352 VGND VGND VPWR VPWR picorv32_352/HI trace_data[29] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_110_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08965_ _03439_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_90_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07916_ _02532_ _02535_ _02470_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_126_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08896_ _03373_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__clkbuf_4
X_07847_ net176 _02466_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_108_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07778_ _02396_ _02397_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__and2_1
X_09517_ cpuregs\[12\]\[14\] cpuregs\[13\]\[14\] cpuregs\[14\]\[14\] cpuregs\[15\]\[14\]
+ _03582_ _03716_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_94_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09448_ _03909_ _03910_ _03436_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09379_ cpuregs\[16\]\[10\] cpuregs\[17\]\[10\] cpuregs\[18\]\[10\] cpuregs\[19\]\[10\]
+ _03586_ _03449_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_135_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11410_ _05304_ _05305_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12390_ cpuregs\[16\]\[15\] cpuregs\[17\]\[15\] cpuregs\[18\]\[15\] cpuregs\[19\]\[15\]
+ _05948_ _06068_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11341_ _05227_ _05246_ _05247_ _05224_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14060_ net1237 _06948_ _01649_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__mux2_1
X_11272_ reg_next_pc\[5\] _03213_ _02945_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__mux2_2
XFILLER_0_132_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13011_ _06642_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__clkbuf_1
X_10223_ _04584_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__clkbuf_1
X_10154_ cpuregs\[30\]\[19\] _03307_ _04537_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ clknet_leaf_85_clk _00620_ VGND VGND VPWR VPWR reg_pc\[8\] sky130_fd_sc_hd__dfxtp_2
X_10085_ _04486_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__buf_4
X_13913_ net696 _06937_ _01566_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__mux2_1
X_14893_ clknet_leaf_112_clk _00551_ VGND VGND VPWR VPWR count_instr\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13844_ net1174 _06937_ _07100_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13775_ _07070_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__clkbuf_1
X_10987_ _05005_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_44_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12726_ _03124_ _06463_ _06465_ _03139_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15514_ clknet_leaf_43_clk _01099_ VGND VGND VPWR VPWR cpuregs\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15445_ clknet_leaf_42_clk _01035_ VGND VGND VPWR VPWR cpuregs\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12657_ cpuregs\[8\]\[27\] cpuregs\[9\]\[27\] cpuregs\[10\]\[27\] cpuregs\[11\]\[27\]
+ _05907_ _03039_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_288 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_127_357 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11608_ _05486_ _05481_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__and2b_1
XFILLER_0_154_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15376_ clknet_leaf_64_clk _00966_ VGND VGND VPWR VPWR reg_sh\[1\] sky130_fd_sc_hd__dfxtp_1
X_12588_ cpuregs\[8\]\[24\] cpuregs\[9\]\[24\] cpuregs\[10\]\[24\] cpuregs\[11\]\[24\]
+ _06061_ _03137_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14327_ _01790_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__clkbuf_1
X_11539_ _05421_ _05424_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold407 cpuregs\[31\]\[2\] VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold418 cpuregs\[12\]\[31\] VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 cpuregs\[20\]\[21\] VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ _01754_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13209_ decoded_imm\[20\] _06752_ _06736_ _06753_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14189_ net940 _06941_ _01710_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _03173_ _03243_ _03244_ _03246_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__a22o_4
X_07701_ _02325_ _02326_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__nor2_1
X_08681_ reg_out\[1\] alu_out_q\[1\] _03174_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07632_ reg_pc\[20\] decoded_imm\[20\] _02247_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_926 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07563_ _02195_ _02197_ _01893_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09302_ _03765_ _03766_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07494_ _02132_ _02133_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09233_ decoded_imm\[6\] net199 VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09164_ _03434_ _03628_ _03630_ _03634_ _03490_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__a311o_1
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08115_ _02720_ _02721_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_390 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_483 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09095_ _03557_ _03567_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_714 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08046_ _02656_ _02657_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_92_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold930 cpuregs\[28\]\[4\] VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold941 cpuregs\[13\]\[14\] VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 cpuregs\[22\]\[12\] VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold963 cpuregs\[12\]\[5\] VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 cpuregs\[6\]\[13\] VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 cpuregs\[21\]\[17\] VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 cpuregs\[10\]\[9\] VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09997_ cpuregs\[24\]\[29\] cpuregs\[25\]\[29\] cpuregs\[26\]\[29\] cpuregs\[27\]\[29\]
+ _03808_ _03812_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_4_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _03403_ _03422_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08879_ _03357_ _03358_ _03293_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__mux2_2
X_10910_ cpuregs\[20\]\[5\] _04829_ _04959_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ count_cycle\[50\] net447 net379 count_cycle\[52\] VGND VGND VPWR VPWR _05707_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_123_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10841_ _04928_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13560_ net997 _06945_ _06946_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_756 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_143_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10772_ net780 _04827_ _04887_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12511_ _06254_ _06256_ _06258_ _06260_ _06151_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13491_ net754 _04850_ _06899_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_631 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15230_ clknet_leaf_77_clk _00823_ VGND VGND VPWR VPWR instr_lh sky130_fd_sc_hd__dfxtp_1
X_12442_ cpuregs\[24\]\[17\] cpuregs\[25\]\[17\] cpuregs\[26\]\[17\] cpuregs\[27\]\[17\]
+ _06074_ _05932_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_152_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15161_ clknet_leaf_50_clk _00786_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dfxtp_2
X_12373_ _05886_ _06118_ _06122_ _05978_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__a311o_2
XFILLER_0_23_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_325 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_50_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14112_ _01678_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__clkbuf_1
X_11324_ _05231_ reg_pc\[20\] VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__or2_1
X_15092_ clknet_leaf_90_clk _07115_ VGND VGND VPWR VPWR reg_out\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14043_ net573 _06931_ _01638_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__mux2_1
X_11255_ _05185_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_152_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10206_ net978 _03248_ _04575_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11186_ _05137_ _05138_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__nor2_1
X_10137_ _04538_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__clkbuf_1
X_14945_ clknet_leaf_120_clk _00603_ VGND VGND VPWR VPWR count_instr\[54\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10068_ _04500_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14876_ clknet_leaf_151_clk _00534_ VGND VGND VPWR VPWR cpuregs\[17\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_161_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13827_ _07097_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13758_ net725 _06987_ _07027_ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_789 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12709_ cpuregs\[28\]\[29\] cpuregs\[29\]\[29\] cpuregs\[30\]\[29\] cpuregs\[31\]\[29\]
+ _06191_ _05914_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13689_ _07024_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15428_ clknet_leaf_148_clk _01018_ VGND VGND VPWR VPWR cpuregs\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15359_ clknet_leaf_68_clk _00949_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold204 cpuregs\[0\]\[9\] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold215 mem_rdata_q\[24\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 cpuregs\[0\]\[26\] VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 cpuregs\[2\]\[5\] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 cpuregs\[11\]\[23\] VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _03447_ _04367_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__or2_1
Xhold259 count_instr\[15\] VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09851_ _03474_ _04292_ _04300_ _04301_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_70_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _03290_ _03291_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09782_ _03574_ _04226_ _04234_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08733_ reg_pc\[8\] _03223_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08664_ latched_branch latched_store VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_105_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_870 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07615_ _02242_ _02245_ _02246_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08595_ cpuregs\[28\]\[3\] cpuregs\[29\]\[3\] cpuregs\[30\]\[3\] cpuregs\[31\]\[3\]
+ _03107_ _03108_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ _02179_ _02182_ cpu_state\[6\] VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_64_704 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_119_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07477_ _01893_ _02110_ _02111_ _02118_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__o31ai_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09216_ cpuregs\[20\]\[5\] cpuregs\[21\]\[5\] cpuregs\[22\]\[5\] cpuregs\[23\]\[5\]
+ _03636_ _03637_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09147_ _03479_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_161_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09078_ cpuregs\[0\]\[2\] cpuregs\[1\]\[2\] cpuregs\[2\]\[2\] cpuregs\[3\]\[2\] _03438_
+ _03549_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_9_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08029_ _02494_ _02569_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold760 cpuregs\[25\]\[8\] VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 cpuregs\[18\]\[18\] VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 net158 VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _05033_ _01884_ _05034_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__and3b_1
Xhold793 cpuregs\[13\]\[8\] VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__dlygate4sd3_1
X_12991_ is_slli_srli_srai _06553_ _06559_ _06632_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__a22o_1
X_11942_ cpuregs\[24\]\[31\] cpuregs\[25\]\[31\] cpuregs\[26\]\[31\] cpuregs\[27\]\[31\]
+ _03594_ _03442_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__mux4_1
X_14730_ clknet_leaf_44_clk _00388_ VGND VGND VPWR VPWR cpuregs\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14661_ clknet_leaf_21_clk _00319_ VGND VGND VPWR VPWR cpuregs\[14\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_706 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11873_ count_cycle\[46\] count_cycle\[47\] _05692_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_158_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ net695 _06981_ _06967_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__mux2_1
X_10824_ net1337 _04879_ _04909_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__mux2_1
X_14592_ clknet_leaf_144_clk _00250_ VGND VGND VPWR VPWR cpuregs\[28\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13543_ _03214_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__buf_2
XFILLER_0_54_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10755_ _03380_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__buf_2
X_13474_ net1331 _04833_ _06888_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__mux2_1
X_10686_ _04834_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15213_ clknet_leaf_101_clk alu_out\[26\] VGND VGND VPWR VPWR alu_out_q\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12425_ cpuregs\[4\]\[17\] cpuregs\[5\]\[17\] cpuregs\[6\]\[17\] cpuregs\[7\]\[17\]
+ _06011_ _06156_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_932 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15144_ clknet_leaf_80_clk _00770_ VGND VGND VPWR VPWR mem_do_prefetch sky130_fd_sc_hd__dfxtp_1
X_12356_ cpuregs\[12\]\[14\] cpuregs\[13\]\[14\] cpuregs\[14\]\[14\] cpuregs\[15\]\[14\]
+ _03107_ _03129_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_39_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11307_ _01884_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__buf_2
X_15075_ clknet_leaf_118_clk _00733_ VGND VGND VPWR VPWR count_cycle\[58\] sky130_fd_sc_hd__dfxtp_1
X_12287_ cpuregs\[28\]\[11\] cpuregs\[29\]\[11\] cpuregs\[30\]\[11\] cpuregs\[31\]\[11\]
+ _05895_ _05929_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14026_ _01632_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11238_ _05174_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ count_instr\[35\] count_instr\[34\] _05116_ _05126_ VGND VGND VPWR VPWR _05127_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14928_ clknet_leaf_116_clk _00586_ VGND VGND VPWR VPWR count_instr\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14859_ clknet_leaf_47_clk _00517_ VGND VGND VPWR VPWR cpuregs\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_07400_ net15 _01937_ _02045_ _01935_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__a22o_1
X_08380_ net224 _02252_ _02933_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_67_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07331_ net23 net130 _01980_ _01940_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07262_ _01917_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09001_ _03475_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__buf_4
XFILLER_0_155_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07193_ mem_do_wdata mem_do_rdata mem_do_rinst _01856_ _01857_ VGND VGND VPWR VPWR
+ _01858_ sky130_fd_sc_hd__o311a_1
XFILLER_0_14_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_13_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09903_ _03454_ _04351_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09834_ cpuregs\[8\]\[24\] cpuregs\[9\]\[24\] cpuregs\[10\]\[24\] cpuregs\[11\]\[24\]
+ _03494_ _03497_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__mux4_1
X_09765_ _01958_ _04210_ _04212_ _03397_ _04217_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_87_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08716_ reg_out\[6\] alu_out_q\[6\] _03174_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ _04084_ _04114_ _04115_ _04150_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__o211a_1
Xrebuffer30 net390 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_1
Xrebuffer41 net401 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08647_ mem_rdata_q\[21\] net14 _03018_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08578_ _03047_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__buf_6
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07529_ _02083_ _02166_ _02085_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10540_ _04753_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10471_ _04716_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _05969_ _05971_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13190_ decoded_imm\[29\] _06740_ _06737_ _06743_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__o22a_1
XFILLER_0_161_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12141_ net249 _05863_ _05903_ _05905_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_131_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12072_ cpuregs\[12\]\[1\] cpuregs\[13\]\[1\] cpuregs\[14\]\[1\] cpuregs\[15\]\[1\]
+ _05816_ _03086_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__mux4_1
Xhold590 cpuregs\[29\]\[16\] VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ _05024_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__clkbuf_1
X_15900_ clknet_leaf_139_clk _01472_ VGND VGND VPWR VPWR cpuregs\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15831_ clknet_leaf_133_clk _01403_ VGND VGND VPWR VPWR cpuregs\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15762_ clknet_leaf_15_clk _01337_ VGND VGND VPWR VPWR cpuregs\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12974_ decoded_imm_j\[11\] _01082_ _03021_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__mux2_1
X_14713_ clknet_leaf_10_clk _00371_ VGND VGND VPWR VPWR cpuregs\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11925_ _05730_ _05731_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__nor2_1
X_15693_ clknet_leaf_142_clk _01268_ VGND VGND VPWR VPWR cpuregs\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11856_ count_cycle\[40\] _05680_ count_cycle\[41\] VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__a21o_1
X_14644_ clknet_leaf_10_clk _00302_ VGND VGND VPWR VPWR cpuregs\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10807_ _04910_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__clkbuf_1
X_14575_ clknet_leaf_43_clk _00233_ VGND VGND VPWR VPWR cpuregs\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11787_ net550 _05634_ _05636_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_119 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_83_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10738_ net833 _04869_ _04861_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13526_ _03178_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_422 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13457_ _06886_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__clkbuf_1
X_10669_ _03193_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_151_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12408_ cpuregs\[8\]\[16\] cpuregs\[9\]\[16\] cpuregs\[10\]\[16\] cpuregs\[11\]\[16\]
+ _06061_ _05917_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13388_ net974 _04883_ _06815_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__mux2_1
Xoutput106 net106 VGND VGND VPWR VPWR mem_la_wdata[18] sky130_fd_sc_hd__clkbuf_4
Xoutput117 net117 VGND VGND VPWR VPWR mem_la_wdata[28] sky130_fd_sc_hd__buf_2
Xoutput128 net128 VGND VGND VPWR VPWR mem_la_wdata[9] sky130_fd_sc_hd__clkbuf_4
X_12339_ _06093_ _06094_ _06095_ _05873_ _03113_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_637 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15127_ clknet_leaf_71_clk _00753_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_1
Xoutput139 net139 VGND VGND VPWR VPWR mem_wdata[13] sky130_fd_sc_hd__buf_2
XFILLER_0_121_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15058_ clknet_leaf_114_clk _00716_ VGND VGND VPWR VPWR count_cycle\[41\] sky130_fd_sc_hd__dfxtp_1
X_14009_ _01623_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__clkbuf_1
X_07880_ _02496_ _02497_ _02498_ _02499_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09550_ decoded_imm\[15\] net177 VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08501_ decoded_imm_j\[17\] _01079_ _03022_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__mux2_1
X_09481_ cpuregs\[16\]\[13\] cpuregs\[17\]\[13\] cpuregs\[18\]\[13\] cpuregs\[19\]\[13\]
+ _03548_ _03549_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_78_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08432_ _02177_ _02979_ _02971_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_144_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_547 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_92_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08363_ _02509_ net212 _02251_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07314_ instr_rdinstr VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__buf_4
X_08294_ _02869_ _02876_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_15_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07245_ _01851_ _01878_ _01903_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07176_ _01839_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09817_ _04244_ _04263_ _04268_ _03396_ _02290_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__o32a_1
X_09748_ _03475_ _04201_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__and2_1
X_09679_ _04128_ _04130_ _04132_ _04134_ _03430_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__a221o_2
XFILLER_0_97_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11710_ _05495_ _05259_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_38_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _05912_ _06431_ _06193_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11641_ _05494_ _05244_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14360_ _01807_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__clkbuf_1
X_11572_ decoded_imm_j\[17\] _05228_ _05446_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13311_ _06809_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__clkbuf_1
X_10523_ _04743_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__clkbuf_1
Xinput19 net418 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
X_14291_ net585 VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_122_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13242_ mem_rdata_q\[24\] _06627_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__and2_1
X_10454_ net729 _03386_ _04672_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13173_ _05860_ decoded_imm_j\[1\] is_slli_srli_srai VGND VGND VPWR VPWR _06730_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10385_ cpuregs\[28\]\[31\] _03386_ _04635_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__mux2_1
X_12124_ _05873_ _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__and2_1
X_12055_ _03113_ _05824_ _03139_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__o21a_1
X_11006_ _05015_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15814_ clknet_leaf_47_clk _01386_ VGND VGND VPWR VPWR cpuregs\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15745_ clknet_leaf_26_clk _01320_ VGND VGND VPWR VPWR cpuregs\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12957_ _06613_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11908_ net476 _05716_ _05719_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_16_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ clknet_leaf_132_clk _01251_ VGND VGND VPWR VPWR cpuregs\[29\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12888_ mem_rdata_q\[23\] mem_rdata_q\[22\] mem_rdata_q\[2\] mem_rdata_q\[3\] VGND
+ VGND VPWR VPWR _06574_ sky130_fd_sc_hd__or4_1
XFILLER_0_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14627_ clknet_leaf_122_clk _00285_ VGND VGND VPWR VPWR cpuregs\[21\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11839_ _05672_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_651 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_138_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14558_ clknet_leaf_145_clk _00216_ VGND VGND VPWR VPWR cpuregs\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_537 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13509_ _06914_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__clkbuf_1
X_14489_ clknet_leaf_2_clk _00147_ VGND VGND VPWR VPWR cpuregs\[30\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_121_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08981_ _00012_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__buf_8
XFILLER_0_139_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07932_ _02544_ _02549_ is_sltiu_bltu_sltu VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__o21a_1
X_07863_ net202 _02482_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09602_ _04058_ _04059_ _03402_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__mux2_1
X_07794_ _02222_ net212 VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09533_ _03581_ _03992_ _03467_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__o21a_1
X_09464_ _03903_ _03908_ _03926_ _03665_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_35_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08415_ _02112_ _02967_ _02951_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__mux2_1
X_09395_ reg_pc\[10\] _03527_ _03859_ _03625_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_539 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08346_ _02482_ _02927_ _02929_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__a21o_1
XFILLER_0_62_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08277_ _02869_ _02870_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07228_ instr_rdcycle _01825_ _01840_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_907 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07159_ instr_rdinstrh instr_rdcycleh instr_rdinstr VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_95_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10170_ _04555_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13860_ _01544_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_161_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12811_ _06532_ mem_rdata_q\[13\] _06533_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_126_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ net776 _06952_ _07075_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15530_ clknet_leaf_124_clk _01115_ VGND VGND VPWR VPWR cpuregs\[24\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12742_ net226 _06481_ _06282_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12673_ _05886_ _06405_ _06409_ _05978_ _06415_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__a311o_4
X_15461_ clknet_leaf_125_clk _01051_ VGND VGND VPWR VPWR cpuregs\[19\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11624_ _05240_ _05490_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__nand2_1
X_14412_ clknet_leaf_63_clk _00070_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15392_ clknet_leaf_94_clk _00982_ VGND VGND VPWR VPWR decoded_imm\[16\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14343_ _01798_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__clkbuf_1
X_11555_ _05285_ _05226_ _05439_ _05300_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_786 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10506_ net1200 _03334_ _04731_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14274_ _01762_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11486_ _05373_ _05374_ _05269_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13225_ decoded_imm\[12\] _06752_ _06735_ _06761_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__o22a_1
X_10437_ _04698_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_789 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_21_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13156_ net131 _05764_ _06721_ _06673_ net712 VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__a32o_1
X_10368_ _04661_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__clkbuf_1
X_12107_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_12 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13087_ net135 _02507_ _06685_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__mux2_1
X_10299_ net1263 _03329_ _04622_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12038_ _05807_ _05809_ mem_do_rinst _05810_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_109_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13989_ _01601_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_38_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15728_ clknet_leaf_0_clk _01303_ VGND VGND VPWR VPWR cpuregs\[22\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15659_ clknet_leaf_3_clk _01234_ VGND VGND VPWR VPWR cpuregs\[29\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_320 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08200_ _02250_ _02798_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_21 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09180_ _01854_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08131_ _02165_ _02466_ _02593_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08062_ _02662_ _02666_ _02660_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpicorv32_320 VGND VGND VPWR VPWR picorv32_320/HI pcpi_insn[30] sky130_fd_sc_hd__conb_1
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_331 VGND VGND VPWR VPWR picorv32_331/HI trace_data[8] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_342 VGND VGND VPWR VPWR picorv32_342/HI trace_data[19] sky130_fd_sc_hd__conb_1
Xpicorv32_353 VGND VGND VPWR VPWR picorv32_353/HI trace_data[30] sky130_fd_sc_hd__conb_1
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08964_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_90_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07915_ _02533_ _02534_ _02467_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__a21o_1
X_08895_ _03261_ _03369_ _03372_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__o21a_1
X_07846_ net208 VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_518 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_79_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07777_ _02277_ net217 VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__nand2_1
X_09516_ _03433_ _03972_ _03974_ _03976_ _03760_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_631 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09447_ cpuregs\[20\]\[12\] cpuregs\[21\]\[12\] cpuregs\[22\]\[12\] cpuregs\[23\]\[12\]
+ _03719_ _03588_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09378_ cpuregs\[20\]\[10\] cpuregs\[21\]\[10\] cpuregs\[22\]\[10\] cpuregs\[23\]\[10\]
+ _03456_ _03441_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_46_172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08329_ _02757_ net226 _02908_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11340_ _05231_ reg_pc\[25\] VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11271_ _05194_ reg_pc\[4\] _01843_ _05198_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13010_ net612 _04829_ _06636_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__mux2_1
X_10222_ net806 _03302_ _04575_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__mux2_1
X_10153_ _04546_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10084_ _04508_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__clkbuf_1
X_14961_ clknet_leaf_82_clk _00619_ VGND VGND VPWR VPWR reg_pc\[7\] sky130_fd_sc_hd__dfxtp_2
X_13912_ _01572_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__clkbuf_1
X_14892_ clknet_leaf_112_clk net495 VGND VGND VPWR VPWR count_instr\[1\] sky130_fd_sc_hd__dfxtp_1
X_13843_ _07106_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10986_ net948 _04837_ _04995_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__mux2_1
X_13774_ net644 _06935_ _07064_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15513_ clknet_leaf_45_clk _01098_ VGND VGND VPWR VPWR cpuregs\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12725_ _03042_ _06464_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15444_ clknet_leaf_42_clk _01034_ VGND VGND VPWR VPWR cpuregs\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12656_ cpuregs\[12\]\[27\] cpuregs\[13\]\[27\] cpuregs\[14\]\[27\] cpuregs\[15\]\[27\]
+ _05834_ _03129_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11607_ _05481_ _05486_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12587_ _06058_ _06332_ _06182_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__o21a_1
X_15375_ clknet_leaf_63_clk _00965_ VGND VGND VPWR VPWR reg_sh\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_25_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14326_ net987 _03247_ _01789_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11538_ _05401_ _05409_ _05423_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold408 cpuregs\[19\]\[4\] VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 cpuregs\[24\]\[31\] VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__dlygate4sd3_1
X_14257_ net563 VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__clkbuf_1
X_11469_ decoded_imm_j\[10\] _05210_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13208_ mem_rdata_q\[20\] _06742_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14188_ _01718_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13139_ net152 net114 _06707_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ reg_pc\[26\] decoded_imm\[26\] VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__and2_1
X_08680_ _03186_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__clkbuf_1
X_07631_ _02260_ _02261_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07562_ _02195_ _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_938 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09301_ _01870_ _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_595 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_154_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_154_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07493_ reg_pc\[12\] decoded_imm\[12\] VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_64_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09232_ _02030_ _03396_ _03694_ _03701_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_90_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09163_ _03455_ _03631_ _03633_ _03468_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08114_ _02706_ _02711_ _02704_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__o21a_1
X_09094_ cpuregs\[24\]\[2\] cpuregs\[25\]\[2\] cpuregs\[26\]\[2\] cpuregs\[27\]\[2\]
+ _03456_ _03441_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08045_ net126 net125 _02609_ _02630_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__or4_4
XFILLER_0_114_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold920 cpuregs\[24\]\[0\] VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 cpuregs\[18\]\[15\] VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold942 cpuregs\[26\]\[17\] VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold953 cpuregs\[1\]\[12\] VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 cpuregs\[9\]\[19\] VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold975 cpuregs\[16\]\[8\] VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 cpuregs\[7\]\[7\] VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 cpuregs\[19\]\[3\] VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ _03446_ _04441_ _03417_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ cpuregs\[4\]\[0\] cpuregs\[5\]\[0\] cpuregs\[6\]\[0\] cpuregs\[7\]\[0\] _03406_
+ _03410_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_4_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ reg_pc\[27\] _03352_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__xor2_1
X_07829_ _02369_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10840_ net1128 _04827_ _04923_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__mux2_1
X_10771_ _04891_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_145_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_145_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12510_ _06073_ _06259_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13490_ _06904_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_807 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12441_ _06026_ _06192_ _06193_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12372_ _06124_ _06126_ _06127_ _03132_ _05815_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15160_ clknet_leaf_50_clk _00785_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11323_ reg_next_pc\[20\] _03309_ _02947_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__mux2_2
X_14111_ net770 _06931_ _01674_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_15091_ clknet_leaf_89_clk _07145_ VGND VGND VPWR VPWR reg_out\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_105_586 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11254_ _05184_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__buf_4
X_14042_ _01641_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10205_ _04563_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11185_ net703 _05135_ _05133_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__o21ai_1
X_10136_ cpuregs\[30\]\[10\] _03248_ _04537_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14944_ clknet_leaf_120_clk _00602_ VGND VGND VPWR VPWR count_instr\[53\] sky130_fd_sc_hd__dfxtp_1
X_10067_ net1225 _03255_ _04498_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14875_ clknet_leaf_158_clk _00533_ VGND VGND VPWR VPWR cpuregs\[17\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13826_ net817 _06987_ _07063_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13757_ _07060_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_136_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_136_clk sky130_fd_sc_hd__clkbuf_2
X_10969_ _04996_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__clkbuf_1
X_12708_ _03132_ _06448_ _05840_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__o21a_1
X_13688_ cpuregs\[23\]\[29\] _06985_ _07014_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15427_ clknet_leaf_157_clk _01017_ VGND VGND VPWR VPWR cpuregs\[18\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12639_ _06380_ _06381_ _06382_ _05873_ _05845_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15358_ clknet_leaf_68_clk _00948_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_124_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold205 mem_rdata_q\[26\] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__buf_1
X_14309_ cpuregs\[10\]\[2\] _03193_ _01778_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold216 count_instr\[22\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ clknet_leaf_78_clk _00881_ VGND VGND VPWR VPWR is_slli_srli_srai sky130_fd_sc_hd__dfxtp_4
Xhold227 cpuregs\[29\]\[25\] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold238 instr_sltu VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 count_instr\[3\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09850_ reg_pc\[24\] _03527_ _03625_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__a21o_1
X_08801_ reg_pc\[17\] reg_pc\[16\] _03279_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09781_ _04228_ _04230_ _04233_ _03575_ _03591_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__a221o_1
X_08732_ reg_pc\[8\] _03223_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__or2_1
X_08663_ _03170_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_105_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07614_ reg_pc\[20\] decoded_imm\[20\] VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08594_ _03050_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07545_ latched_is_lh _02181_ _02085_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_127_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_127_clk sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_119_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_716 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_76_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07476_ _01944_ _02112_ _02114_ _01928_ _02117_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_9_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_689 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09215_ _03500_ _03684_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_579 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09146_ _01978_ _02008_ _03617_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09077_ cpuregs\[4\]\[2\] cpuregs\[5\]\[2\] cpuregs\[6\]\[2\] cpuregs\[7\]\[2\] _03548_
+ _03549_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08028_ _02044_ _02492_ _02618_ _02641_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__a31o_1
Xhold750 cpuregs\[27\]\[17\] VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 cpuregs\[3\]\[25\] VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 cpuregs\[7\]\[31\] VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold783 cpuregs\[26\]\[5\] VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 cpuregs\[3\]\[23\] VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__dlygate4sd3_1
X_09979_ decoded_imm\[29\] _02369_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12990_ _06536_ _06533_ net242 _06566_ _06544_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__a32o_1
X_11941_ _03402_ _05745_ _03603_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ clknet_leaf_138_clk _00318_ VGND VGND VPWR VPWR cpuregs\[14\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11872_ net545 _05692_ _05694_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_158_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13611_ _03359_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10823_ _04918_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__clkbuf_1
X_14591_ clknet_leaf_131_clk _00249_ VGND VGND VPWR VPWR cpuregs\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_118_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_118_clk sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13542_ _06934_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__clkbuf_1
X_10754_ _04880_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_401 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13473_ _06895_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__clkbuf_1
X_10685_ cpuregs\[26\]\[7\] _04833_ _04819_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__mux2_1
X_15212_ clknet_leaf_101_clk alu_out\[25\] VGND VGND VPWR VPWR alu_out_q\[25\] sky130_fd_sc_hd__dfxtp_1
X_12424_ _05927_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_136_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15143_ clknet_leaf_105_clk _00769_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12355_ _06107_ _06109_ _06110_ _03128_ _03035_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11306_ _05188_ reg_pc\[15\] VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__or2_1
X_12286_ _06023_ _06044_ _05927_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__o21a_1
X_15074_ clknet_leaf_118_clk _00732_ VGND VGND VPWR VPWR count_cycle\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11237_ _05172_ _05113_ _05173_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__and3b_1
X_14025_ net1267 _06981_ _01624_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ count_instr\[37\] count_instr\[36\] VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__and2_1
X_10119_ net1155 _03194_ _04526_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__mux2_1
X_11099_ net1398 _05075_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14927_ clknet_leaf_111_clk _00585_ VGND VGND VPWR VPWR count_instr\[36\] sky130_fd_sc_hd__dfxtp_1
X_14858_ clknet_leaf_46_clk _00516_ VGND VGND VPWR VPWR cpuregs\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_11_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13809_ _07088_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_206 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_109_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_109_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_67_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14789_ clknet_leaf_151_clk _00447_ VGND VGND VPWR VPWR cpuregs\[16\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07330_ net10 _01937_ _01979_ _01935_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07261_ is_jalr_addi_slti_sltiu_xori_ori_andi is_lui_auipc_jal VGND VGND VPWR VPWR
+ _01917_ sky130_fd_sc_hd__or2_2
XFILLER_0_155_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_115_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09000_ cpu_state\[4\] _01854_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_14_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_602 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07192_ net33 net134 VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__and2_2
XFILLER_0_5_356 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_54_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_41_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09902_ cpuregs\[12\]\[26\] cpuregs\[13\]\[26\] cpuregs\[14\]\[26\] cpuregs\[15\]\[26\]
+ _03598_ _03716_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09833_ _01958_ _04270_ _04272_ _03651_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__a32o_1
X_09764_ _04215_ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_87_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08715_ _03216_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09695_ _04082_ _04147_ _04087_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__or3b_1
Xrebuffer20 _05700_ VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer31 net391 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer42 net402 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08646_ _03161_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _03095_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07528_ _01846_ _01848_ net24 _01933_ net6 VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07459_ _02065_ _02099_ _02101_ _01927_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10470_ net1245 _03221_ _04709_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_106_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09129_ _03554_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__buf_6
XFILLER_0_150_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12140_ decoded_imm\[5\] _05904_ _01841_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12071_ _03034_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold580 cpuregs\[9\]\[2\] VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 cpuregs\[18\]\[27\] VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ net822 _04873_ _05017_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__mux2_1
X_15830_ clknet_leaf_140_clk _01402_ VGND VGND VPWR VPWR cpuregs\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15761_ clknet_leaf_16_clk _01336_ VGND VGND VPWR VPWR cpuregs\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12973_ _06621_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14712_ clknet_leaf_17_clk _00370_ VGND VGND VPWR VPWR cpuregs\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11924_ net567 _05728_ _05141_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__o21ai_1
X_15692_ clknet_leaf_14_clk _01267_ VGND VGND VPWR VPWR cpuregs\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14643_ clknet_leaf_31_clk _00301_ VGND VGND VPWR VPWR cpuregs\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11855_ count_cycle\[40\] count_cycle\[41\] _05680_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10806_ cpuregs\[16\]\[20\] _04860_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__mux2_1
X_14574_ clknet_leaf_45_clk _00232_ VGND VGND VPWR VPWR cpuregs\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11786_ count_cycle\[19\] _05634_ _05622_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_693 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_138_773 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13525_ _06922_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_36 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10737_ _03340_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_11_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13456_ net778 _04883_ _06851_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10668_ _04822_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12407_ _06058_ _06160_ _03123_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13387_ _06849_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__clkbuf_1
X_10599_ net687 _03194_ _04782_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__mux2_1
Xoutput107 net107 VGND VGND VPWR VPWR mem_la_wdata[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput118 net118 VGND VGND VPWR VPWR mem_la_wdata[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15126_ clknet_leaf_72_clk _00752_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_4
Xoutput129 net129 VGND VGND VPWR VPWR mem_la_write sky130_fd_sc_hd__buf_2
X_12338_ cpuregs\[28\]\[13\] cpuregs\[29\]\[13\] _03085_ VGND VGND VPWR VPWR _06095_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_649 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15057_ clknet_leaf_114_clk _00715_ VGND VGND VPWR VPWR count_cycle\[40\] sky130_fd_sc_hd__dfxtp_1
X_12269_ cpuregs\[24\]\[10\] cpuregs\[25\]\[10\] cpuregs\[26\]\[10\] cpuregs\[27\]\[10\]
+ _03095_ _05932_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__mux4_1
X_14008_ cpuregs\[5\]\[19\] _06964_ _01613_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__mux2_1
X_15959_ clknet_leaf_133_clk _01531_ VGND VGND VPWR VPWR cpuregs\[10\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08500_ _03026_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__buf_1
X_09480_ _03807_ _03941_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08431_ reg_next_pc\[15\] reg_out\[15\] _02969_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__mux2_2
XFILLER_0_148_515 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_74 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_59_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08362_ _02937_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07313_ _01846_ _01958_ _01961_ _01927_ _01963_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_610 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08293_ _02340_ _02883_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_899 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07244_ _01902_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_15_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07175_ _01839_ _01840_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__nand2_2
XFILLER_0_30_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_100_824 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09816_ _01977_ _04265_ _04267_ _03485_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__a31o_1
X_09747_ _03472_ _04191_ _04200_ _03525_ reg_pc\[21\] VGND VGND VPWR VPWR _04201_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09678_ _03435_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _03045_ _03146_ _03034_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11640_ _05508_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_25_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11571_ _05452_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13310_ net988 _04873_ _06802_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_294 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10522_ net1223 _03386_ _04708_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__mux2_1
X_14290_ _01770_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_133_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10453_ _04706_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__clkbuf_1
X_13241_ decoded_imm\[5\] _06626_ _06770_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__o21a_1
X_10384_ _04669_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__clkbuf_1
X_13172_ _01944_ net434 _03670_ _06729_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__a31o_1
X_12123_ cpuregs\[4\]\[5\] cpuregs\[5\]\[5\] _03085_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__mux2_1
X_12054_ cpuregs\[12\]\[0\] cpuregs\[13\]\[0\] cpuregs\[14\]\[0\] cpuregs\[15\]\[0\]
+ _03150_ _03151_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__mux4_1
X_11005_ net1182 _04856_ _05006_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15813_ clknet_leaf_40_clk _01385_ VGND VGND VPWR VPWR cpuregs\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15744_ clknet_leaf_50_clk _01319_ VGND VGND VPWR VPWR cpuregs\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12956_ net427 _01071_ _06587_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11907_ net476 _05716_ _01905_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__o21ai_1
X_15675_ clknet_leaf_129_clk _01250_ VGND VGND VPWR VPWR cpuregs\[29\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ mem_rdata_q\[4\] mem_rdata_q\[5\] mem_rdata_q\[6\] VGND VGND VPWR VPWR _06573_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_142_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_68_671 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14626_ clknet_leaf_127_clk _00284_ VGND VGND VPWR VPWR cpuregs\[21\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11838_ _05670_ _05625_ _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__and3b_1
XFILLER_0_28_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14557_ clknet_leaf_3_clk _00215_ VGND VGND VPWR VPWR cpuregs\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11769_ count_cycle\[13\] count_cycle\[14\] _05620_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_40_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13508_ net1157 _04867_ _06910_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14488_ clknet_leaf_154_clk _00146_ VGND VGND VPWR VPWR cpuregs\[30\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13439_ _06877_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_379 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_125_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15109_ clknet_leaf_103_clk _07133_ VGND VGND VPWR VPWR reg_out\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_21 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08980_ _03454_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__buf_8
X_07931_ is_slti_blt_slt instr_bge _02550_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__mux2_1
X_07862_ net234 VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__clkbuf_4
X_09601_ cpuregs\[0\]\[17\] cpuregs\[1\]\[17\] cpuregs\[2\]\[17\] cpuregs\[3\]\[17\]
+ _03405_ _03496_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07793_ net180 net212 VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__or2_1
X_09532_ cpuregs\[8\]\[15\] cpuregs\[9\]\[15\] cpuregs\[10\]\[15\] cpuregs\[11\]\[15\]
+ _03582_ _03583_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__mux4_1
X_09463_ reg_pc\[12\] _03528_ _03925_ _03626_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_35_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08414_ reg_next_pc\[10\] reg_out\[10\] _02949_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__mux2_1
X_09394_ _03473_ _03850_ _03858_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__and3_2
XFILLER_0_19_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08345_ _01880_ _02503_ _02482_ _01913_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_31_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08276_ _02331_ _02868_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_916 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07227_ _01820_ _01870_ _01887_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__nor3_1
XFILLER_0_116_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07158_ _01824_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_95_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_161_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12810_ mem_rdata_q\[12\] VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13790_ _07078_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_126_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12741_ _05900_ _06467_ _06480_ _01918_ decoded_imm\[30\] VGND VGND VPWR VPWR _06481_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15460_ clknet_leaf_148_clk _01050_ VGND VGND VPWR VPWR cpuregs\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12672_ _06411_ _06413_ _06414_ _03149_ _05815_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__o221a_1
X_14411_ clknet_leaf_63_clk _00069_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11623_ _05240_ _05490_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__nor2_1
X_15391_ clknet_leaf_94_clk _00981_ VGND VGND VPWR VPWR decoded_imm\[17\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_25_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_22_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_527 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ net960 _03301_ _01789_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11554_ _05430_ _05431_ _05437_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_108_798 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10505_ _04734_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14273_ net674 VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11485_ _05373_ _05374_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13224_ _06525_ decoded_imm_j\[12\] _06738_ _06533_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__a22o_1
X_10436_ cpuregs\[21\]\[22\] _03329_ _04695_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13155_ _01818_ _05763_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__nor2_1
X_10367_ net1213 _03329_ _04658_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12106_ _00008_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__inv_2
X_13086_ _06684_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__buf_4
X_10298_ _04624_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_89_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12037_ _01891_ _03389_ _05809_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_109_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13988_ _01612_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15727_ clknet_leaf_0_clk _01302_ VGND VGND VPWR VPWR cpuregs\[22\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12939_ _06604_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15658_ clknet_leaf_1_clk _01233_ VGND VGND VPWR VPWR cpuregs\[29\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14609_ clknet_leaf_36_clk _00267_ VGND VGND VPWR VPWR cpuregs\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15589_ clknet_leaf_33_clk _01164_ VGND VGND VPWR VPWR cpuregs\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_33 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_2
X_08130_ _02732_ _02734_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__nand2_1
X_08061_ _02670_ _02671_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_310 VGND VGND VPWR VPWR picorv32_310/HI pcpi_insn[20] sky130_fd_sc_hd__conb_1
Xpicorv32_321 VGND VGND VPWR VPWR picorv32_321/HI pcpi_insn[31] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_332 VGND VGND VPWR VPWR picorv32_332/HI trace_data[9] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_343 VGND VGND VPWR VPWR picorv32_343/HI trace_data[20] sky130_fd_sc_hd__conb_1
XFILLER_0_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpicorv32_354 VGND VGND VPWR VPWR picorv32_354/HI trace_data[31] sky130_fd_sc_hd__conb_1
XFILLER_0_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08963_ _00012_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__buf_8
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07914_ _02139_ _02472_ _02463_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__or3b_1
X_08894_ _03370_ _03371_ _03261_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07845_ _02139_ _02463_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_3_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07776_ _02277_ net217 VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__or2_1
X_09515_ _03593_ _03975_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_906 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09446_ cpuregs\[16\]\[12\] cpuregs\[17\]\[12\] cpuregs\[18\]\[12\] cpuregs\[19\]\[12\]
+ _03587_ _03588_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_137_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09377_ _01854_ _03835_ _03836_ _03841_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08328_ _02584_ _02914_ _02915_ _02917_ net450 VGND VGND VPWR VPWR alu_out\[30\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08259_ _02853_ _02854_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11270_ _01872_ _05197_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10221_ _04583_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_563 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10152_ cpuregs\[30\]\[18\] _03302_ _04537_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ cpuregs\[12\]\[19\] _03307_ _04498_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__mux2_1
X_14960_ clknet_leaf_82_clk _00618_ VGND VGND VPWR VPWR reg_pc\[6\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_128_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13911_ net626 _06935_ _01566_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__mux2_1
X_14891_ clknet_leaf_111_clk _00549_ VGND VGND VPWR VPWR count_instr\[0\] sky130_fd_sc_hd__dfxtp_1
X_13842_ net1313 _06935_ _07100_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_69_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13773_ _07069_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__clkbuf_1
X_10985_ _05004_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__clkbuf_1
X_15512_ clknet_leaf_37_clk _01097_ VGND VGND VPWR VPWR cpuregs\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12724_ cpuregs\[8\]\[30\] cpuregs\[9\]\[30\] cpuregs\[10\]\[30\] cpuregs\[11\]\[30\]
+ _03038_ _03039_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15443_ clknet_leaf_26_clk _01033_ VGND VGND VPWR VPWR cpuregs\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12655_ _06394_ _06396_ _06397_ _03061_ _03035_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11606_ _05446_ _05454_ _05482_ _05485_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__a31oi_2
X_15374_ clknet_leaf_93_clk _00964_ VGND VGND VPWR VPWR latched_rd\[4\] sky130_fd_sc_hd__dfxtp_4
X_12586_ cpuregs\[12\]\[24\] cpuregs\[13\]\[24\] cpuregs\[14\]\[24\] cpuregs\[15\]\[24\]
+ _03133_ _03134_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14325_ _01777_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__buf_4
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11537_ _05422_ _05413_ _05409_ _05407_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__o31a_1
XFILLER_0_151_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold409 cpuregs\[5\]\[11\] VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ _01753_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__clkbuf_1
X_11468_ decoded_imm_j\[10\] _05210_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_59_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13207_ _06531_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__clkbuf_4
X_10419_ cpuregs\[21\]\[14\] _03275_ _04684_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__mux2_1
X_14187_ net1115 _06939_ _01710_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__mux2_1
X_11399_ _05191_ _05195_ _05197_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__and3_1
X_13138_ _06712_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ instr_sltu _06671_ _06530_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07630_ reg_pc\[21\] decoded_imm\[21\] VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__nand2_1
X_07561_ _02196_ _02174_ _02172_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__o21ai_1
X_09300_ _03765_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07492_ reg_pc\[12\] decoded_imm\[12\] VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09231_ _03699_ _03700_ _03486_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_326 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_119_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09162_ _03436_ _03632_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08113_ _02718_ _02719_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__nand2_1
X_09093_ _03401_ _03565_ _03418_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08044_ _02573_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold910 cpuregs\[16\]\[27\] VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 cpuregs\[28\]\[3\] VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold932 cpuregs\[24\]\[2\] VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 cpuregs\[27\]\[5\] VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 cpuregs\[22\]\[5\] VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 cpuregs\[11\]\[30\] VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 cpuregs\[11\]\[13\] VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 cpuregs\[22\]\[0\] VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 cpuregs\[23\]\[15\] VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ cpuregs\[28\]\[29\] cpuregs\[29\]\[29\] cpuregs\[30\]\[29\] cpuregs\[31\]\[29\]
+ _03586_ _03449_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08946_ _03415_ _03416_ _03420_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_4_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ reg_out\[27\] alu_out_q\[27\] _03176_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__mux2_1
X_07828_ _02447_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07759_ net24 _02202_ _02180_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_714 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10770_ cpuregs\[16\]\[3\] _04825_ _04887_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09429_ _03868_ _03887_ _03892_ _03396_ _02125_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__o32a_1
XFILLER_0_94_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12440_ _03054_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12371_ cpuregs\[16\]\[14\] cpuregs\[17\]\[14\] cpuregs\[18\]\[14\] cpuregs\[19\]\[14\]
+ _05984_ _05985_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14110_ _01677_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__clkbuf_1
X_11322_ _05227_ _05233_ _05234_ _05224_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__o211a_1
X_15090_ clknet_leaf_90_clk _07144_ VGND VGND VPWR VPWR reg_out\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_105_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14041_ cpuregs\[6\]\[2\] _06929_ _01638_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__mux2_1
X_11253_ _01872_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__clkbuf_4
X_10204_ _04574_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__clkbuf_1
X_11184_ count_instr\[42\] count_instr\[41\] net1418 VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__and3_1
X_10135_ _04525_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_66_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14943_ clknet_leaf_119_clk _00601_ VGND VGND VPWR VPWR count_instr\[52\] sky130_fd_sc_hd__dfxtp_1
X_10066_ _04499_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__clkbuf_1
X_14874_ clknet_leaf_158_clk _00532_ VGND VGND VPWR VPWR cpuregs\[17\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13825_ _07096_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_97_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13756_ cpuregs\[29\]\[29\] _06985_ _07050_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10968_ net968 _04817_ _04995_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12707_ cpuregs\[16\]\[29\] cpuregs\[17\]\[29\] cpuregs\[18\]\[29\] cpuregs\[19\]\[29\]
+ _05984_ _05985_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13687_ _07023_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_75_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10899_ _04958_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15426_ clknet_leaf_157_clk _01016_ VGND VGND VPWR VPWR cpuregs\[18\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12638_ cpuregs\[28\]\[26\] cpuregs\[29\]\[26\] _03085_ VGND VGND VPWR VPWR _06382_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_649 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15357_ clknet_leaf_49_clk _00947_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dfxtp_1
X_12569_ _06138_ _06315_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14308_ _01780_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__clkbuf_1
Xhold206 count_cycle\[43\] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ clknet_leaf_77_clk _00880_ VGND VGND VPWR VPWR is_lb_lh_lw_lbu_lhu sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_57_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold217 cpuregs\[6\]\[4\] VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold228 cpuregs\[0\]\[8\] VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold239 cpuregs\[28\]\[29\] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ net524 VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08800_ reg_pc\[16\] _03279_ reg_pc\[17\] VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__a21oi_1
X_09780_ _04231_ _04232_ _03579_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08731_ reg_out\[8\] alu_out_q\[8\] _03174_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__mux2_1
X_08662_ decoded_imm_j\[4\] _01086_ _03169_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__mux2_2
XFILLER_0_89_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07613_ _02218_ _02232_ _02233_ _02244_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08593_ cpuregs\[24\]\[3\] cpuregs\[25\]\[3\] cpuregs\[26\]\[3\] cpuregs\[27\]\[3\]
+ _03092_ _03087_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__mux4_1
X_07544_ _01844_ _01848_ net25 net7 _01933_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07475_ _02115_ _02116_ _01955_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_107_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09214_ cpuregs\[16\]\[5\] cpuregs\[17\]\[5\] cpuregs\[18\]\[5\] cpuregs\[19\]\[5\]
+ _03458_ _03461_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_430 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_627 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09145_ _03479_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09076_ _00013_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__buf_8
XFILLER_0_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_513 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08027_ _02562_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__clkbuf_4
Xhold740 cpuregs\[31\]\[6\] VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 cpuregs\[24\]\[11\] VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 cpuregs\[1\]\[29\] VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 cpuregs\[8\]\[30\] VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 cpuregs\[20\]\[17\] VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 net142 VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ decoded_imm\[29\] _02369_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__nor2_1
X_08929_ _00012_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__buf_6
X_11940_ cpuregs\[28\]\[31\] cpuregs\[29\]\[31\] cpuregs\[30\]\[31\] cpuregs\[31\]\[31\]
+ _03601_ _03583_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_28_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ count_cycle\[46\] _05692_ _05622_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__o21ai_1
X_13610_ _06980_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_158_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ net1271 _04877_ _04909_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__mux2_1
X_14590_ clknet_leaf_146_clk _00248_ VGND VGND VPWR VPWR cpuregs\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13541_ net910 _06933_ _06925_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__mux2_1
X_10753_ net1091 _04879_ _04861_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13472_ cpuregs\[9\]\[6\] _04831_ _06888_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__mux2_1
X_10684_ _03227_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_178 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15211_ clknet_leaf_102_clk alu_out\[24\] VGND VGND VPWR VPWR alu_out_q\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12423_ _06176_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_136_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15142_ clknet_leaf_104_clk _00768_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_1
X_12354_ cpuregs\[0\]\[14\] cpuregs\[1\]\[14\] cpuregs\[2\]\[14\] cpuregs\[3\]\[14\]
+ _05819_ _03125_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_885 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ _05221_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15073_ clknet_leaf_119_clk _00731_ VGND VGND VPWR VPWR count_cycle\[56\] sky130_fd_sc_hd__dfxtp_1
X_12285_ cpuregs\[16\]\[11\] cpuregs\[17\]\[11\] cpuregs\[18\]\[11\] cpuregs\[19\]\[11\]
+ _05948_ _05925_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14024_ _01631_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11236_ count_instr\[57\] net385 count_instr\[58\] VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ net442 VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10118_ _04528_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__clkbuf_1
X_11098_ count_instr\[16\] _05075_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14926_ clknet_leaf_116_clk _00584_ VGND VGND VPWR VPWR count_instr\[35\] sky130_fd_sc_hd__dfxtp_1
X_10049_ _04490_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_1
X_14857_ clknet_leaf_19_clk _00515_ VGND VGND VPWR VPWR cpuregs\[20\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_13808_ cpuregs\[3\]\[21\] _06969_ _07086_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__mux2_1
X_14788_ clknet_leaf_148_clk _00446_ VGND VGND VPWR VPWR cpuregs\[16\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13739_ _07051_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07260_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_61_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15409_ clknet_leaf_46_clk _00999_ VGND VGND VPWR VPWR cpuregs\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_07191_ mem_state\[1\] mem_state\[0\] VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_14_614 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_143_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_14_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_13_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_541 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09901_ _03433_ _04345_ _04347_ _04349_ _03760_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_585 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09832_ _04281_ _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09763_ _04177_ _04181_ _04178_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__a21oi_1
X_08714_ net1252 _03215_ _03185_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _04026_ _04148_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__nand2_1
Xrebuffer10 net385 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_87_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer21 _05139_ VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_1
Xrebuffer32 net392 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_1
X_08645_ decoded_imm_j\[11\] _01082_ _03022_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__mux2_1
Xrebuffer43 net403 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08576_ _03046_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__buf_8
XFILLER_0_77_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_577 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07527_ net176 VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_641 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07458_ _02083_ _02100_ _02085_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07389_ _01970_ _02028_ _02029_ _02035_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_118_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09128_ _03581_ _03599_ _03547_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_693 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09059_ net171 _01978_ _03479_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_630 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12070_ _02507_ _01841_ _05814_ _05839_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__a22o_1
Xhold570 cpuregs\[1\]\[9\] VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_376 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold581 cpuregs\[8\]\[8\] VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 cpuregs\[2\]\[30\] VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _05023_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__clkbuf_1
X_15760_ clknet_leaf_6_clk _01335_ VGND VGND VPWR VPWR cpuregs\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12972_ decoded_imm_j\[18\] _01080_ _03021_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11923_ count_cycle\[60\] count_cycle\[61\] count_cycle\[62\] _05724_ VGND VGND VPWR
+ VPWR _05730_ sky130_fd_sc_hd__and4_1
X_14711_ clknet_leaf_13_clk _00369_ VGND VGND VPWR VPWR cpuregs\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_15691_ clknet_leaf_8_clk _01266_ VGND VGND VPWR VPWR cpuregs\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14642_ clknet_leaf_56_clk _00300_ VGND VGND VPWR VPWR cpuregs\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11854_ net506 net370 _05682_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10805_ _04886_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__buf_4
XFILLER_0_83_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14573_ clknet_leaf_44_clk _00231_ VGND VGND VPWR VPWR cpuregs\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11785_ _05634_ _05635_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13524_ net871 _04883_ _06887_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__mux2_1
X_10736_ _04868_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13455_ _06885_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_149_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10667_ net1268 _04821_ _04819_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12406_ cpuregs\[12\]\[16\] cpuregs\[13\]\[16\] cpuregs\[14\]\[16\] cpuregs\[15\]\[16\]
+ _05913_ _05994_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13386_ net947 _04881_ _06815_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10598_ _04784_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__clkbuf_1
X_15125_ clknet_leaf_72_clk _00751_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_1
Xoutput108 net108 VGND VGND VPWR VPWR mem_la_wdata[1] sky130_fd_sc_hd__clkbuf_4
X_12337_ _05974_ cpuregs\[30\]\[13\] _05896_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput119 net119 VGND VGND VPWR VPWR mem_la_wdata[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15056_ clknet_leaf_114_clk _00714_ VGND VGND VPWR VPWR count_cycle\[39\] sky130_fd_sc_hd__dfxtp_1
X_12268_ _06026_ _06027_ _03081_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__o21a_1
X_14007_ _01622_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_184 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11219_ _05160_ _05161_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__nor2_1
X_12199_ _03134_ _05960_ _03050_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__a21o_1
Xoutput90 net90 VGND VGND VPWR VPWR mem_la_addr[4] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_158_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15958_ clknet_leaf_139_clk _01530_ VGND VGND VPWR VPWR cpuregs\[10\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14909_ clknet_leaf_119_clk _00567_ VGND VGND VPWR VPWR count_instr\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15889_ clknet_leaf_14_clk _01461_ VGND VGND VPWR VPWR cpuregs\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ _02978_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_19_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_86 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08361_ _02503_ net211 _02251_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07312_ reg_pc\[1\] decoded_imm\[1\] _01962_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08292_ _02884_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_622 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07243_ instr_jal _01901_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__nor2_2
XFILLER_0_61_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07174_ cpu_state\[2\] VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_836 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09815_ _04145_ _04266_ _03670_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__o21ai_1
X_09746_ _04193_ _04195_ _04197_ _04199_ _03429_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__a221o_1
X_09677_ cpuregs\[24\]\[19\] cpuregs\[25\]\[19\] cpuregs\[26\]\[19\] cpuregs\[27\]\[19\]
+ _03548_ _03549_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__mux4_1
X_08628_ cpuregs\[16\]\[4\] cpuregs\[17\]\[4\] cpuregs\[18\]\[4\] cpuregs\[19\]\[4\]
+ _03062_ _03063_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_38_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ reg_sh\[3\] reg_sh\[2\] net521 VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__or3b_1
X_11570_ decoded_imm_j\[18\] _05230_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10521_ _04742_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13240_ _06763_ net719 _06733_ mem_rdata_q\[25\] _06541_ VGND VGND VPWR VPWR _06770_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_133_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10452_ net1388 _03381_ _04672_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13171_ _01944_ _06726_ _06727_ _06728_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__o2bb2a_1
X_10383_ net756 _03381_ _04635_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__mux2_1
X_12122_ _03090_ _05881_ _05885_ _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__o211a_1
X_12053_ _03128_ _05822_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__or2_1
X_11004_ _05014_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15812_ clknet_leaf_26_clk _01384_ VGND VGND VPWR VPWR cpuregs\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12955_ _06612_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__clkbuf_1
X_15743_ clknet_leaf_49_clk _01318_ VGND VGND VPWR VPWR cpuregs\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11906_ _05718_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_240 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15674_ clknet_leaf_142_clk _01249_ VGND VGND VPWR VPWR cpuregs\[29\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12886_ mem_rdata_q\[25\] mem_rdata_q\[24\] _06540_ _06571_ VGND VGND VPWR VPWR _06572_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_16_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_650 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11837_ count_cycle\[34\] _05667_ count_cycle\[35\] VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__a21o_1
X_14625_ clknet_leaf_147_clk _00283_ VGND VGND VPWR VPWR cpuregs\[21\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14556_ clknet_leaf_3_clk _00214_ VGND VGND VPWR VPWR cpuregs\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11768_ net570 _05620_ _05623_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_722 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10719_ net1087 _04856_ _04840_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__mux2_1
X_13507_ _06913_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14487_ clknet_leaf_3_clk _00145_ VGND VGND VPWR VPWR cpuregs\[30\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11699_ _05551_ _05554_ _05563_ _05570_ _05553_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_99_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13438_ net1173 _04865_ _06874_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_799 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xrebuffer1 _05686_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__buf_1
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13369_ _06840_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15108_ clknet_leaf_103_clk _07132_ VGND VGND VPWR VPWR reg_out\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_33 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15039_ clknet_leaf_122_clk _00697_ VGND VGND VPWR VPWR count_cycle\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07930_ _02545_ net238 _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__or3_1
X_07861_ _02479_ _02480_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__and2_1
X_09600_ cpuregs\[4\]\[17\] cpuregs\[5\]\[17\] cpuregs\[6\]\[17\] cpuregs\[7\]\[17\]
+ _03405_ _03496_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07792_ _02222_ net212 VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__or2b_1
XFILLER_0_155_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09531_ _03989_ _03990_ _03579_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09462_ _03574_ _03916_ _03924_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__and3_2
XFILLER_0_78_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08413_ _02966_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_1
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09393_ _03852_ _03854_ _03857_ _03426_ _03489_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__a221o_1
X_08344_ _02476_ _02927_ _02928_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__a21o_1
XFILLER_0_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_686 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08275_ _02331_ _02868_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_196 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_105_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07226_ mem_do_prefetch _01886_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_358 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_15_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_15_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07157_ instr_jal _01823_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_95_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09729_ _04180_ _04181_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_126_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ _05886_ _06469_ _06473_ _05978_ _06479_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__a311o_1
XFILLER_0_96_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12671_ cpuregs\[16\]\[27\] cpuregs\[17\]\[27\] cpuregs\[18\]\[27\] cpuregs\[19\]\[27\]
+ _05921_ _05985_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14410_ clknet_leaf_57_clk _00031_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__dfxtp_4
X_11622_ _05496_ _05499_ _05367_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__o21a_1
X_15390_ clknet_leaf_94_clk _00980_ VGND VGND VPWR VPWR decoded_imm\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_355 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14341_ _01797_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_42_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11553_ _05434_ _05436_ _05367_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_135_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10504_ net721 _03329_ _04731_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14272_ _01761_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__clkbuf_1
X_11484_ _05360_ _05363_ _05359_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13223_ decoded_imm\[13\] _06752_ _06735_ _06760_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__o22a_1
XFILLER_0_150_544 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10435_ _04697_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13154_ net477 _05767_ _06720_ _05763_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__o22a_1
X_10366_ _04660_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__clkbuf_1
X_12105_ _05870_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_1
X_13085_ _01821_ _05763_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__nor2_2
X_10297_ cpuregs\[2\]\[21\] _03322_ _04622_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__mux2_1
X_12036_ _01840_ _05808_ _01915_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_109_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_18_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13987_ net1004 _06943_ _01602_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15726_ clknet_leaf_1_clk _01301_ VGND VGND VPWR VPWR cpuregs\[22\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12938_ decoded_imm_j\[14\] _01076_ _03169_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15657_ clknet_leaf_1_clk _01232_ VGND VGND VPWR VPWR cpuregs\[29\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_119 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_666 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12869_ _06546_ net242 _06565_ _06562_ net429 VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14608_ clknet_leaf_30_clk _00266_ VGND VGND VPWR VPWR cpuregs\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_99_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15588_ clknet_leaf_43_clk _01163_ VGND VGND VPWR VPWR cpuregs\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14539_ clknet_leaf_50_clk _00197_ VGND VGND VPWR VPWR cpuregs\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08060_ net202 _02669_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_300 VGND VGND VPWR VPWR picorv32_300/HI pcpi_insn[10] sky130_fd_sc_hd__conb_1
XFILLER_0_114_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpicorv32_311 VGND VGND VPWR VPWR picorv32_311/HI pcpi_insn[21] sky130_fd_sc_hd__conb_1
Xpicorv32_322 VGND VGND VPWR VPWR picorv32_322/HI pcpi_valid sky130_fd_sc_hd__conb_1
XFILLER_0_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_333 VGND VGND VPWR VPWR picorv32_333/HI trace_data[10] sky130_fd_sc_hd__conb_1
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_344 VGND VGND VPWR VPWR picorv32_344/HI trace_data[21] sky130_fd_sc_hd__conb_1
Xpicorv32_355 VGND VGND VPWR VPWR picorv32_355/HI trace_data[32] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_110_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08962_ _03436_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__buf_6
X_07913_ _02154_ _02471_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_90_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ reg_pc\[29\] _03364_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07844_ _02139_ _02463_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__or2_1
X_07775_ net186 net218 VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_108_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09514_ cpuregs\[28\]\[14\] cpuregs\[29\]\[14\] cpuregs\[30\]\[14\] cpuregs\[31\]\[14\]
+ _03598_ _03460_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09445_ _02065_ _03905_ _03907_ _03488_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_149_655 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_115_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09376_ _03074_ _03838_ _03840_ _01953_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08327_ _02595_ _02916_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_105_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08258_ net187 _02852_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__or2_1
X_07209_ mem_do_wdata net34 cpu_state\[5\] _01862_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_104_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08189_ _02410_ _02581_ _02789_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__a21o_1
X_10220_ net953 _03295_ _04575_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_575 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10151_ _04545_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ _04507_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ _01571_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__clkbuf_1
X_14890_ clknet_leaf_73_clk _00548_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dfxtp_4
XPHY_EDGE_ROW_113_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13841_ _07105_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_141_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13772_ net810 _06933_ _07064_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__mux2_1
X_10984_ net620 _04835_ _04995_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15511_ clknet_leaf_27_clk _01096_ VGND VGND VPWR VPWR cpuregs\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12723_ cpuregs\[12\]\[30\] cpuregs\[13\]\[30\] cpuregs\[14\]\[30\] cpuregs\[15\]\[30\]
+ _05834_ _03129_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ cpuregs\[0\]\[27\] cpuregs\[1\]\[27\] cpuregs\[2\]\[27\] cpuregs\[3\]\[27\]
+ _05819_ _03086_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__mux4_1
X_15442_ clknet_leaf_29_clk _01032_ VGND VGND VPWR VPWR cpuregs\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_686 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11605_ decoded_imm_j\[20\] _05235_ _05482_ _05483_ _05484_ VGND VGND VPWR VPWR _05485_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12585_ _06329_ _06330_ _03082_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__mux2_1
X_15373_ clknet_leaf_93_clk _00963_ VGND VGND VPWR VPWR latched_rd\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_108_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11536_ decoded_imm_j\[13\] VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__inv_2
X_14324_ _01788_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_122_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14255_ net587 VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__clkbuf_1
X_11467_ _05040_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_59_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13206_ decoded_imm\[21\] _06740_ _06736_ _06751_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__o22a_1
XFILLER_0_151_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10418_ _04688_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__clkbuf_1
X_14186_ _01717_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__clkbuf_1
X_11398_ _05292_ _05294_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__or2_1
X_13137_ net151 net113 _06707_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10349_ _04651_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ is_beq_bne_blt_bge_bltu_bgeu instr_slt instr_sltiu instr_slti VGND VGND VPWR
+ VPWR _06671_ sky130_fd_sc_hd__or4_1
X_12019_ _05796_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_131_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07560_ reg_pc\[15\] decoded_imm\[15\] VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__and2_1
X_15709_ clknet_leaf_58_clk _01284_ VGND VGND VPWR VPWR cpuregs\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_07491_ _02071_ _02124_ _02128_ _02131_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_817 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09230_ _03695_ _03698_ _03397_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_338 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09161_ cpuregs\[8\]\[4\] cpuregs\[9\]\[4\] cpuregs\[10\]\[4\] cpuregs\[11\]\[4\]
+ _03463_ _03464_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__mux4_1
XFILLER_0_134_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08112_ net175 _02717_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09092_ cpuregs\[28\]\[2\] cpuregs\[29\]\[2\] cpuregs\[30\]\[2\] cpuregs\[31\]\[2\]
+ _03404_ _03408_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08043_ _02478_ _02581_ _02654_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__a21o_1
Xhold900 cpuregs\[23\]\[20\] VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 cpuregs\[14\]\[14\] VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 cpuregs\[17\]\[29\] VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold933 net55 VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 cpuregs\[19\]\[8\] VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 cpuregs\[24\]\[14\] VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 cpuregs\[17\]\[17\] VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold977 cpuregs\[6\]\[21\] VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _03435_ _04439_ _03425_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__o21a_1
Xhold988 cpuregs\[2\]\[24\] VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 cpuregs\[31\]\[0\] VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08945_ _03419_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_4_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ _03356_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07827_ _02437_ _02443_ _02446_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07758_ net194 VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07689_ net188 VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__buf_4
XFILLER_0_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09428_ _01977_ _03889_ _03891_ _03486_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09359_ _02112_ _03770_ _03824_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_47_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12370_ _03087_ _06125_ _03153_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11321_ _05231_ reg_pc\[19\] VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14040_ _01640_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11252_ net466 _05181_ _05183_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10203_ net826 _03241_ _04564_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__mux2_1
X_11183_ _05135_ _05136_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10134_ _04536_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__clkbuf_1
X_14942_ clknet_leaf_119_clk _00600_ VGND VGND VPWR VPWR count_instr\[51\] sky130_fd_sc_hd__dfxtp_1
X_10065_ net1117 _03248_ _04498_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__mux2_1
X_14873_ clknet_leaf_158_clk _00531_ VGND VGND VPWR VPWR cpuregs\[17\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13824_ cpuregs\[3\]\[29\] _06985_ _07086_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_249 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13755_ _07059_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__clkbuf_1
X_10967_ _04994_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12706_ _03113_ _06446_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13686_ net805 _06983_ _07014_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__mux2_1
X_10898_ _04485_ _04671_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__nor2_2
X_15425_ clknet_leaf_159_clk _01015_ VGND VGND VPWR VPWR cpuregs\[18\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12637_ _05974_ cpuregs\[30\]\[26\] _05896_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12568_ cpuregs\[8\]\[23\] cpuregs\[9\]\[23\] cpuregs\[10\]\[23\] cpuregs\[11\]\[23\]
+ _06061_ _03137_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__mux4_1
X_15356_ clknet_leaf_49_clk _00946_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11519_ _05185_ _05405_ _05406_ _05257_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__o211a_1
X_14307_ net864 _03188_ _01778_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12499_ _06058_ _06248_ _06182_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15287_ clknet_leaf_78_clk _00001_ VGND VGND VPWR VPWR is_lui_auipc_jal sky130_fd_sc_hd__dfxtp_2
Xhold207 cpuregs\[4\]\[3\] VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 cpuregs\[0\]\[31\] VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold229 cpuregs\[22\]\[1\] VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14238_ _01744_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_350 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14169_ net1131 _06989_ _01673_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08730_ _03229_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08661_ _03021_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__buf_4
X_07612_ _02194_ _02208_ _02243_ _02241_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_105_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08592_ _03083_ _03105_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07543_ _02179_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07474_ count_instr\[10\] _01949_ count_cycle\[10\] _01951_ VGND VGND VPWR VPWR _02116_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09213_ _03434_ _03677_ _03679_ _03682_ _03490_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__a221o_2
XFILLER_0_45_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_119_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_483 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_17_634 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_442 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09144_ _03482_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09075_ _00012_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__buf_8
XFILLER_0_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08026_ _02635_ _02638_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold730 cpuregs\[26\]\[2\] VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 cpuregs\[14\]\[4\] VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold752 cpuregs\[22\]\[30\] VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 cpuregs\[13\]\[29\] VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 is_alu_reg_reg VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 cpuregs\[24\]\[25\] VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 cpuregs\[30\]\[2\] VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__dlygate4sd3_1
X_09977_ net253 _03396_ _04404_ _04423_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__o22a_1
X_08928_ _03402_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__buf_4
X_08859_ net955 _03341_ _03315_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ net1396 _05689_ _05693_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__o21a_1
X_10821_ _04917_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_258 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10752_ _03373_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__clkbuf_4
X_13540_ _03208_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13471_ _06894_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__clkbuf_1
X_10683_ _04832_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15210_ clknet_leaf_102_clk alu_out\[23\] VGND VGND VPWR VPWR alu_out_q\[23\] sky130_fd_sc_hd__dfxtp_1
X_12422_ net247 _06175_ _06052_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12353_ _03134_ _06108_ _03050_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__a21o_1
X_15141_ clknet_leaf_104_clk _00767_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_294 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11304_ reg_next_pc\[15\] _03277_ _02946_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15072_ clknet_leaf_119_clk _00730_ VGND VGND VPWR VPWR count_cycle\[55\] sky130_fd_sc_hd__dfxtp_1
X_12284_ _03143_ _06042_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14023_ net1134 _06979_ _01624_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11235_ count_instr\[58\] count_instr\[57\] _05168_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__and3_1
X_11166_ _05124_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsplit2 decoder_trigger VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_2
X_10117_ net625 _03189_ _04526_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__mux2_1
X_11097_ _05075_ _05076_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__nor2_1
X_14925_ clknet_leaf_116_clk _00583_ VGND VGND VPWR VPWR count_instr\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10048_ net922 _03194_ _04487_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold90 net169 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
X_14856_ clknet_leaf_22_clk _00514_ VGND VGND VPWR VPWR cpuregs\[20\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13807_ _07087_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__clkbuf_1
X_14787_ clknet_leaf_124_clk _00445_ VGND VGND VPWR VPWR cpuregs\[16\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11999_ _05786_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13738_ net930 _06966_ _07050_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_58_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13669_ _06991_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15408_ clknet_leaf_46_clk _00998_ VGND VGND VPWR VPWR cpuregs\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07190_ mem_state\[1\] mem_state\[0\] VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_626 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_115_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15339_ clknet_leaf_69_clk _00929_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09900_ _03593_ _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_597 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09831_ _04273_ _04274_ _04280_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_96 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09762_ _04213_ _04214_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__nand2_1
X_08713_ _03214_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__buf_2
X_09693_ _04054_ _04147_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xrebuffer11 _05680_ VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_87_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer22 _05139_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_1
X_08644_ _03160_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__buf_1
Xrebuffer33 net393 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_1
Xrebuffer44 net404 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08575_ _03090_ _03093_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07526_ _02161_ _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07457_ _01845_ _01848_ net18 net32 _01933_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__a32o_1
XFILLER_0_107_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07388_ _01954_ _02034_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09127_ cpuregs\[16\]\[3\] cpuregs\[17\]\[3\] cpuregs\[18\]\[3\] cpuregs\[19\]\[3\]
+ _03598_ _03460_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09058_ _03529_ _03530_ _03398_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08009_ net198 _02623_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold560 net62 VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 cpuregs\[29\]\[20\] VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ cpuregs\[17\]\[25\] _04871_ _05017_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold582 cpuregs\[17\]\[4\] VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 cpuregs\[31\]\[23\] VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__dlygate4sd3_1
X_12971_ _06620_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
X_14710_ clknet_leaf_12_clk _00368_ VGND VGND VPWR VPWR cpuregs\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11922_ _05728_ _05729_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__nor2_1
X_15690_ clknet_leaf_7_clk _01265_ VGND VGND VPWR VPWR cpuregs\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_14641_ clknet_leaf_34_clk _00299_ VGND VGND VPWR VPWR cpuregs\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11853_ net1407 net370 _05622_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10804_ _04908_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ net1258 _05631_ _05169_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__o21ai_1
X_14572_ clknet_leaf_26_clk _00230_ VGND VGND VPWR VPWR cpuregs\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13523_ _06921_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__clkbuf_1
X_10735_ net1253 _04867_ _04861_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13454_ net1348 _04881_ _06851_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__mux2_1
X_10666_ _03188_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_11_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_153_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12405_ _06157_ _06158_ _06014_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__mux2_1
X_13385_ _06848_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10597_ net1136 _03189_ _04782_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_277 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_51_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15124_ clknet_leaf_72_clk _00750_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
Xoutput109 net109 VGND VGND VPWR VPWR mem_la_wdata[20] sky130_fd_sc_hd__buf_2
X_12336_ cpuregs\[31\]\[13\] _03092_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__or2b_1
X_12267_ cpuregs\[28\]\[10\] cpuregs\[29\]\[10\] cpuregs\[30\]\[10\] cpuregs\[31\]\[10\]
+ _05895_ _05929_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__mux4_1
X_15055_ clknet_leaf_113_clk _00713_ VGND VGND VPWR VPWR count_cycle\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11218_ net549 _05158_ _05133_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__o21ai_1
X_14006_ net1284 _06962_ _01613_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__mux2_1
X_12198_ cpuregs\[6\]\[8\] cpuregs\[7\]\[8\] _03084_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__mux2_1
Xoutput80 net80 VGND VGND VPWR VPWR mem_la_addr[24] sky130_fd_sc_hd__buf_2
Xoutput91 net91 VGND VGND VPWR VPWR mem_la_addr[5] sky130_fd_sc_hd__clkbuf_4
X_11149_ count_instr\[32\] count_instr\[31\] _05109_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15957_ clknet_leaf_14_clk _01529_ VGND VGND VPWR VPWR cpuregs\[10\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14908_ clknet_leaf_121_clk _00566_ VGND VGND VPWR VPWR count_instr\[17\] sky130_fd_sc_hd__dfxtp_1
X_15888_ clknet_leaf_17_clk _01460_ VGND VGND VPWR VPWR cpuregs\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14839_ clknet_leaf_153_clk _00497_ VGND VGND VPWR VPWR cpuregs\[20\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08360_ _02936_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_1
XFILLER_0_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07311_ reg_pc\[1\] decoded_imm\[1\] cpu_state\[3\] VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__o21ai_1
X_08291_ _02340_ _02883_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_128_274 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07242_ decoder_trigger VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07173_ net34 VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_100_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09814_ _02340_ _03770_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__nor2_1
X_09745_ _03435_ _04198_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__or2_1
X_09676_ _03401_ _04131_ _03418_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__o21a_1
X_08627_ cpuregs\[20\]\[4\] cpuregs\[21\]\[4\] cpuregs\[22\]\[4\] cpuregs\[23\]\[4\]
+ _03095_ _03144_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_38_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08558_ _03077_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07509_ count_cycle\[13\] _02051_ _02146_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08489_ _03019_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__buf_1
XFILLER_0_119_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_107_403 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10520_ net748 _03381_ _04708_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10451_ _04705_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_150_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13170_ is_slli_srli_srai decoded_imm_j\[11\] _02065_ VGND VGND VPWR VPWR _06728_
+ sky130_fd_sc_hd__a21o_1
X_10382_ _04668_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12121_ _03123_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12052_ cpuregs\[8\]\[0\] cpuregs\[9\]\[0\] cpuregs\[10\]\[0\] cpuregs\[11\]\[0\]
+ _03107_ _03129_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__mux4_1
Xhold390 cpuregs\[27\]\[28\] VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net1325 _04854_ _05006_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15811_ clknet_leaf_52_clk _01383_ VGND VGND VPWR VPWR cpuregs\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15742_ clknet_leaf_19_clk _01317_ VGND VGND VPWR VPWR cpuregs\[22\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12954_ mem_rdata_q\[9\] net32 _06589_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__mux2_1
X_11905_ _05716_ _01842_ _05717_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__and3b_1
X_15673_ clknet_leaf_145_clk _01248_ VGND VGND VPWR VPWR cpuregs\[29\]\[26\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_230 _03581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12885_ mem_rdata_q\[0\] mem_rdata_q\[1\] VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_241 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ clknet_leaf_147_clk _00282_ VGND VGND VPWR VPWR cpuregs\[21\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ count_cycle\[34\] count_cycle\[35\] net367 VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14555_ clknet_leaf_7_clk _00213_ VGND VGND VPWR VPWR cpuregs\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11767_ count_cycle\[13\] _05620_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13506_ cpuregs\[9\]\[22\] _04865_ _06910_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10718_ _03301_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14486_ clknet_leaf_2_clk _00144_ VGND VGND VPWR VPWR cpuregs\[30\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11698_ _05251_ _05253_ _05494_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13437_ _06876_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer2 _05132_ VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10649_ net724 _03355_ _04804_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13368_ cpuregs\[19\]\[21\] _04863_ _06838_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15107_ clknet_leaf_103_clk _07131_ VGND VGND VPWR VPWR reg_out\[25\] sky130_fd_sc_hd__dfxtp_1
X_12319_ _06067_ _06070_ _06072_ _06076_ _03080_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__a221o_2
XFILLER_0_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13299_ _06803_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15038_ clknet_leaf_122_clk _00696_ VGND VGND VPWR VPWR count_cycle\[21\] sky130_fd_sc_hd__dfxtp_1
X_07860_ _02112_ net248 VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__nand2_1
X_07791_ net181 net213 VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__or2_1
X_09530_ cpuregs\[0\]\[15\] cpuregs\[1\]\[15\] cpuregs\[2\]\[15\] cpuregs\[3\]\[15\]
+ _03439_ _03576_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__mux4_1
X_09461_ _03918_ _03920_ _03923_ _03433_ _03591_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08412_ _02099_ _02965_ _02951_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09392_ _03855_ _03856_ _03446_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_47_846 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08343_ _01880_ _02507_ _02476_ _01913_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08274_ net221 _02867_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_442 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_61_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07225_ mem_do_rinst _01855_ _01858_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07156_ instr_auipc instr_lui VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__or2_2
XFILLER_0_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_483 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07989_ _02590_ _02591_ _02588_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__o21ai_1
X_09728_ _04180_ _04181_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_126_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ decoded_imm\[19\] net181 VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12670_ _03087_ _06412_ _03153_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__a21o_1
X_11621_ _05496_ _05499_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14340_ net896 _03294_ _01789_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11552_ _05434_ _05436_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_42_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10503_ _04733_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14271_ net614 VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__clkbuf_1
X_11483_ _05371_ _05372_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__nor2_1
X_10434_ cpuregs\[21\]\[21\] _03322_ _04695_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__mux2_1
X_13222_ _06525_ decoded_imm_j\[13\] _06738_ mem_rdata_q\[13\] VGND VGND VPWR VPWR
+ _06760_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10365_ net631 _03322_ _04658_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13153_ _01822_ net130 _01818_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_150_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12104_ net250 _05869_ _05863_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__mux2_1
X_13084_ _06683_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__clkbuf_1
X_10296_ _04623_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__clkbuf_1
X_12035_ is_sll_srl_sra _01916_ _01906_ _01908_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13986_ _01611_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__clkbuf_1
X_15725_ clknet_leaf_153_clk _01300_ VGND VGND VPWR VPWR cpuregs\[22\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12937_ _06603_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15656_ clknet_leaf_33_clk _01231_ VGND VGND VPWR VPWR cpuregs\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12868_ is_alu_reg_reg _06528_ _06534_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__and3_1
XFILLER_0_158_678 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_146_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14607_ clknet_leaf_38_clk _00265_ VGND VGND VPWR VPWR cpuregs\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11819_ count_cycle\[28\] _05655_ count_cycle\[29\] VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__a21o_1
X_15587_ clknet_leaf_46_clk _01162_ VGND VGND VPWR VPWR cpuregs\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _01067_ _01068_ _01066_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_99_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14538_ clknet_leaf_48_clk _00196_ VGND VGND VPWR VPWR cpuregs\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14469_ clknet_leaf_137_clk _00127_ VGND VGND VPWR VPWR cpuregs\[12\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_301 VGND VGND VPWR VPWR picorv32_301/HI pcpi_insn[11] sky130_fd_sc_hd__conb_1
XFILLER_0_12_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpicorv32_312 VGND VGND VPWR VPWR picorv32_312/HI pcpi_insn[22] sky130_fd_sc_hd__conb_1
XFILLER_0_51_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_323 VGND VGND VPWR VPWR picorv32_323/HI trace_data[0] sky130_fd_sc_hd__conb_1
Xpicorv32_334 VGND VGND VPWR VPWR picorv32_334/HI trace_data[11] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpicorv32_345 VGND VGND VPWR VPWR picorv32_345/HI trace_data[22] sky130_fd_sc_hd__conb_1
XFILLER_0_12_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpicorv32_356 VGND VGND VPWR VPWR picorv32_356/HI trace_data[33] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_110_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08961_ _03435_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07912_ _02165_ _02466_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_90_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08892_ reg_pc\[29\] _03364_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07843_ net206 VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__clkbuf_4
X_07774_ _02392_ _02393_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_160_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09513_ _03414_ _03973_ _03419_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_157_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_157_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09444_ _03824_ _03906_ _03483_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_818 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_59_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09375_ _02125_ _03479_ _03839_ _03482_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_90_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08326_ _02560_ _02568_ _02445_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08257_ net187 _02852_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07208_ _01866_ _01868_ _01870_ _01872_ _01820_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_178 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08188_ _02237_ net213 _02598_ _02641_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10150_ net1278 _03295_ _04537_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10081_ net918 _03302_ _04498_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13840_ net1002 _06933_ _07100_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_148_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_148_clk sky130_fd_sc_hd__clkbuf_2
X_13771_ _07068_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10983_ _05003_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15510_ clknet_leaf_53_clk _01095_ VGND VGND VPWR VPWR cpuregs\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12722_ _06458_ _06460_ _06461_ _03061_ _03034_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__o221a_1
XFILLER_0_155_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15441_ clknet_leaf_47_clk _01031_ VGND VGND VPWR VPWR cpuregs\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ _05925_ _06395_ _03037_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_26_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11604_ _05461_ _05474_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__and2_1
X_15372_ clknet_leaf_93_clk _00962_ VGND VGND VPWR VPWR latched_rd\[2\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12584_ cpuregs\[0\]\[24\] cpuregs\[1\]\[24\] cpuregs\[2\]\[24\] cpuregs\[3\]\[24\]
+ _06055_ _05829_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_108_553 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14323_ net1355 _03240_ _01778_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11535_ _05419_ _05420_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_156_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14254_ _01752_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__clkbuf_1
X_11466_ _05258_ net651 _05343_ _05357_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13205_ mem_rdata_q\[21\] _06742_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10417_ cpuregs\[21\]\[13\] _03268_ _04684_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__mux2_1
X_14185_ net1098 _06937_ _01710_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11397_ _05276_ _05281_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__nand2_1
X_13136_ _06711_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__clkbuf_1
X_10348_ cpuregs\[28\]\[13\] _03268_ _04647_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__mux2_1
X_10279_ _04614_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__clkbuf_1
X_13067_ net1403 _06513_ _06523_ _06629_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12018_ net53 net84 _05766_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_139_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_139_clk sky130_fd_sc_hd__clkbuf_2
X_13969_ cpuregs\[5\]\[0\] _06923_ _01602_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__mux2_1
X_15708_ clknet_leaf_133_clk _01283_ VGND VGND VPWR VPWR cpuregs\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_07490_ _02018_ _02130_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__or2_2
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15639_ clknet_leaf_128_clk _01214_ VGND VGND VPWR VPWR cpuregs\[23\]\[24\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09160_ cpuregs\[12\]\[4\] cpuregs\[13\]\[4\] cpuregs\[14\]\[4\] cpuregs\[15\]\[4\]
+ _03458_ _03461_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08111_ net175 _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09091_ _03413_ _03563_ _03425_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08042_ _02082_ _02476_ _02598_ _02563_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__a31o_1
XFILLER_0_141_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold901 cpuregs\[14\]\[9\] VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold912 cpuregs\[16\]\[28\] VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 cpuregs\[3\]\[14\] VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold934 cpuregs\[16\]\[30\] VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold945 cpuregs\[5\]\[15\] VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 cpuregs\[18\]\[17\] VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 cpuregs\[30\]\[0\] VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 cpuregs\[16\]\[29\] VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ cpuregs\[16\]\[29\] cpuregs\[17\]\[29\] cpuregs\[18\]\[29\] cpuregs\[19\]\[29\]
+ _03548_ _03549_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__mux4_1
Xhold989 cpuregs\[24\]\[30\] VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08944_ _03418_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_4_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ net705 _03355_ _03315_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__mux2_1
X_07826_ _02444_ _02445_ _02394_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_123_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07757_ _02377_ _02378_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_123_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07688_ _01945_ _02313_ _02314_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__and3_1
X_09427_ _03771_ _03890_ _03670_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09358_ _02082_ _03479_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__nor2_1
X_08309_ net223 _02890_ _02757_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09289_ _03402_ _03756_ _03603_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_138_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11320_ reg_next_pc\[19\] _03304_ _02947_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__mux2_2
XFILLER_0_90_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_498 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_133_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11251_ net466 _05181_ _05036_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_132_375 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_120_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10202_ _04573_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__clkbuf_1
X_11182_ net1008 net405 _05133_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__o21ai_1
X_10133_ net1028 _03241_ _04526_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14941_ clknet_leaf_120_clk _00599_ VGND VGND VPWR VPWR count_instr\[50\] sky130_fd_sc_hd__dfxtp_1
X_10064_ _04486_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__buf_4
X_14872_ clknet_leaf_151_clk _00530_ VGND VGND VPWR VPWR cpuregs\[17\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_13823_ _07095_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13754_ net903 _06983_ _07050_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10966_ _04562_ _04885_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__nor2_4
XFILLER_0_39_930 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_128_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12705_ cpuregs\[20\]\[29\] cpuregs\[21\]\[29\] cpuregs\[22\]\[29\] cpuregs\[23\]\[29\]
+ _03095_ _03144_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13685_ _07022_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__clkbuf_1
X_10897_ _04957_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15424_ clknet_leaf_159_clk _01014_ VGND VGND VPWR VPWR cpuregs\[18\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12636_ cpuregs\[31\]\[26\] _03092_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__or2b_1
XFILLER_0_72_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_884 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15355_ clknet_leaf_68_clk _00945_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dfxtp_1
X_12567_ _06058_ _06313_ _06182_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14306_ _01779_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_318 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11518_ _05031_ reg_next_pc\[13\] VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__or2_1
X_15286_ clknet_leaf_82_clk _00879_ VGND VGND VPWR VPWR decoded_imm\[0\] sky130_fd_sc_hd__dfxtp_2
X_12498_ cpuregs\[12\]\[20\] cpuregs\[13\]\[20\] cpuregs\[14\]\[20\] cpuregs\[15\]\[20\]
+ _03133_ _05994_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__mux4_1
Xhold208 count_cycle\[62\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 count_instr\[30\] VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14237_ net1277 _06989_ _01709_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__mux2_1
X_11449_ _05285_ _05207_ _05341_ _05300_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_896 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14168_ _01707_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__clkbuf_1
X_13119_ _06702_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__clkbuf_1
X_14099_ net726 _06987_ _01637_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__mux2_1
X_08660_ _03168_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__buf_1
X_07611_ reg_pc\[17\] decoded_imm\[17\] VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08591_ _03106_ _03109_ _03035_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07542_ _02178_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_226 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07473_ count_instr\[42\] _01946_ _01947_ count_cycle\[42\] VGND VGND VPWR VPWR _02115_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_516 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09212_ _03448_ _03681_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_456 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_45_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_646 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_115_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09143_ _03609_ _03612_ _03614_ _01870_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_454 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_127_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09074_ _03425_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08025_ _02635_ _02638_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold720 cpuregs\[22\]\[22\] VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 cpuregs\[4\]\[8\] VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 cpuregs\[15\]\[4\] VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold753 cpuregs\[8\]\[22\] VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 cpuregs\[1\]\[28\] VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold775 cpuregs\[5\]\[26\] VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 cpuregs\[23\]\[7\] VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 cpuregs\[6\]\[31\] VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ _03672_ _04422_ _03486_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08927_ _03401_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__buf_8
X_08858_ _03340_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07809_ net188 net220 VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _03277_ _03280_ _03261_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__mux2_4
XFILLER_0_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10820_ net1269 _04875_ _04909_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_209 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10751_ _04878_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_55_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13470_ net1255 _04829_ _06888_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__mux2_1
X_10682_ net1095 _04831_ _04819_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12421_ _06132_ _06165_ _06174_ _06153_ decoded_imm\[16\] VGND VGND VPWR VPWR _06175_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15140_ clknet_leaf_104_clk _00766_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_153_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12352_ cpuregs\[6\]\[14\] cpuregs\[7\]\[14\] _03084_ VGND VGND VPWR VPWR _06108_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11303_ _05194_ net720 _01843_ _05220_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_39_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15071_ clknet_leaf_119_clk _00729_ VGND VGND VPWR VPWR count_cycle\[54\] sky130_fd_sc_hd__dfxtp_1
X_12283_ cpuregs\[20\]\[11\] cpuregs\[21\]\[11\] cpuregs\[22\]\[11\] cpuregs\[23\]\[11\]
+ _05921_ _05922_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__mux4_1
X_14022_ _01630_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__clkbuf_1
X_11234_ net499 net369 _05171_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__a21oi_1
X_11165_ _01884_ _05122_ _05123_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ _04527_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__clkbuf_1
X_11096_ net618 _05073_ _05044_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__o21ai_1
X_14924_ clknet_leaf_116_clk _00582_ VGND VGND VPWR VPWR count_instr\[33\] sky130_fd_sc_hd__dfxtp_1
X_10047_ _04489_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__clkbuf_1
Xhold80 decoded_rd\[3\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 _02444_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
X_14855_ clknet_leaf_130_clk _00513_ VGND VGND VPWR VPWR cpuregs\[20\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_13806_ cpuregs\[3\]\[20\] _06966_ _07086_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14786_ clknet_leaf_125_clk _00444_ VGND VGND VPWR VPWR cpuregs\[16\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11998_ net43 net74 _05785_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13737_ _07027_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_67_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10949_ _04985_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_911 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_45_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13668_ _07013_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15407_ clknet_leaf_92_clk _00997_ VGND VGND VPWR VPWR decoded_imm\[1\] sky130_fd_sc_hd__dfxtp_2
X_12619_ _06357_ _06359_ _06361_ _06363_ _06151_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_14_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_26_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13599_ _03333_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__buf_2
XFILLER_0_42_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_81_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15338_ clknet_leaf_69_clk _00928_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15269_ clknet_leaf_86_clk _00862_ VGND VGND VPWR VPWR decoded_imm_j\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_481 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09830_ _04273_ _04274_ _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09761_ decoded_imm\[22\] net185 VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__or2_1
X_08712_ _03211_ _03212_ _03173_ _03213_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__a2bb2o_2
X_09692_ _04088_ _04116_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer12 _05680_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_1
Xrebuffer23 net381 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_1
X_08643_ mem_rdata_q\[20\] net13 _03018_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__mux2_1
Xrebuffer34 net394 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_1
Xrebuffer45 _05127_ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08574_ cpuregs\[0\]\[3\] cpuregs\[1\]\[3\] cpuregs\[2\]\[3\] cpuregs\[3\]\[3\] _03092_
+ _03087_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07525_ _02162_ _02152_ _02149_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07456_ net202 VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07387_ _01942_ _02030_ _02033_ cpu_state\[6\] VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09126_ _03554_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__buf_8
XFILLER_0_115_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09057_ _03398_ _03529_ _03530_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08008_ net249 _02622_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_131_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold550 cpuregs\[25\]\[6\] VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold561 cpuregs\[10\]\[25\] VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 cpuregs\[4\]\[30\] VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 cpuregs\[6\]\[12\] VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 cpuregs\[13\]\[17\] VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ cpuregs\[0\]\[28\] cpuregs\[1\]\[28\] cpuregs\[2\]\[28\] cpuregs\[3\]\[28\]
+ _03680_ _03443_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__mux4_1
X_12970_ decoded_imm_j\[17\] _01079_ _03021_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__mux2_1
X_11921_ net691 _05726_ _05141_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14640_ clknet_leaf_32_clk _00298_ VGND VGND VPWR VPWR cpuregs\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11852_ net371 _05681_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__nor2_1
X_10803_ net1058 _04858_ _04898_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ clknet_leaf_52_clk _00229_ VGND VGND VPWR VPWR cpuregs\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11783_ count_cycle\[16\] count_cycle\[17\] count_cycle\[18\] _05628_ VGND VGND VPWR
+ VPWR _05634_ sky130_fd_sc_hd__and4_4
Xclkbuf_leaf_52_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_138_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13522_ net1031 _04881_ _06887_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__mux2_1
X_10734_ _03333_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_126_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13453_ _06884_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__clkbuf_1
X_10665_ _04820_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12404_ cpuregs\[0\]\[16\] cpuregs\[1\]\[16\] cpuregs\[2\]\[16\] cpuregs\[3\]\[16\]
+ _06055_ _05909_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__mux4_1
XFILLER_0_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13384_ cpuregs\[19\]\[29\] _04879_ _06838_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_651 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_744 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10596_ _04783_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15123_ clknet_leaf_72_clk _00749_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12335_ _05969_ _06091_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_492 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15054_ clknet_leaf_114_clk _00712_ VGND VGND VPWR VPWR count_cycle\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12266_ _03082_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__buf_4
X_14005_ _01621_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_1
X_11217_ count_instr\[52\] count_instr\[51\] _05156_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__and3_1
Xoutput70 net70 VGND VGND VPWR VPWR mem_la_addr[14] sky130_fd_sc_hd__clkbuf_4
X_12197_ _05871_ _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput81 net81 VGND VGND VPWR VPWR mem_la_addr[25] sky130_fd_sc_hd__buf_2
Xoutput92 net92 VGND VGND VPWR VPWR mem_la_addr[6] sky130_fd_sc_hd__clkbuf_4
X_11148_ net1188 _05109_ _05111_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11079_ count_instr\[10\] _05062_ _05044_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__o21ai_1
X_15956_ clknet_leaf_15_clk _01528_ VGND VGND VPWR VPWR cpuregs\[10\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14907_ clknet_leaf_121_clk _00565_ VGND VGND VPWR VPWR count_instr\[16\] sky130_fd_sc_hd__dfxtp_1
X_15887_ clknet_leaf_14_clk _01459_ VGND VGND VPWR VPWR cpuregs\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14838_ clknet_leaf_0_clk _00496_ VGND VGND VPWR VPWR cpuregs\[20\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_630 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14769_ clknet_leaf_27_clk _00427_ VGND VGND VPWR VPWR cpuregs\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_2
X_07310_ net12 net130 _01960_ _01940_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_551 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_18_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08290_ net222 _02882_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_56 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07241_ _01885_ _01900_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07172_ _01827_ _01828_ _01832_ _01837_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__or4_2
XFILLER_0_152_790 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_111_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09813_ _02306_ _03481_ _04264_ _03483_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__a211o_1
X_09744_ cpuregs\[24\]\[21\] cpuregs\[25\]\[21\] cpuregs\[26\]\[21\] cpuregs\[27\]\[21\]
+ _03808_ _03812_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__mux4_1
X_09675_ cpuregs\[28\]\[19\] cpuregs\[29\]\[19\] cpuregs\[30\]\[19\] cpuregs\[31\]\[19\]
+ _03554_ _03459_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__mux4_1
X_08626_ _03052_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_38_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _03072_ _03076_ _01944_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_2
X_07508_ count_instr\[13\] _02054_ count_cycle\[45\] _02055_ VGND VGND VPWR VPWR _02147_
+ sky130_fd_sc_hd__a22o_1
X_08488_ mem_rdata_q\[15\] net407 _03018_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_702 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_147_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_107_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07439_ latched_is_lh latched_is_lb VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__or2b_2
XFILLER_0_52_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_99_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10450_ net1046 _03374_ _04695_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_278 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09109_ _03413_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__clkbuf_8
X_10381_ net598 _03374_ _04658_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__mux2_1
X_12120_ _05882_ _05883_ _05884_ _05873_ _03083_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12051_ _03061_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__or2_1
Xhold380 cpuregs\[22\]\[20\] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 cpuregs\[10\]\[26\] VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ _05013_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15810_ clknet_leaf_50_clk _01382_ VGND VGND VPWR VPWR cpuregs\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15741_ clknet_leaf_23_clk _01316_ VGND VGND VPWR VPWR cpuregs\[22\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12953_ _06611_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11904_ count_cycle\[55\] _05706_ _05713_ count_cycle\[56\] VGND VGND VPWR VPWR _05717_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15672_ clknet_leaf_131_clk _01247_ VGND VGND VPWR VPWR cpuregs\[29\]\[25\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_220 _06182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12884_ is_alu_reg_imm _06545_ _06566_ _06570_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__a31o_1
*XANTENNA_231 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_242 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14623_ clknet_leaf_122_clk _00281_ VGND VGND VPWR VPWR cpuregs\[21\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11835_ net501 net368 _05669_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_16_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_64_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ clknet_leaf_6_clk _00212_ VGND VGND VPWR VPWR cpuregs\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11766_ _01839_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13505_ _06912_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__clkbuf_1
X_10717_ _04855_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__clkbuf_1
X_14485_ clknet_leaf_1_clk _00143_ VGND VGND VPWR VPWR cpuregs\[30\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11697_ _05253_ _05255_ _05548_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_64_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13436_ net1286 _04863_ _06874_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10648_ _04810_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer3 _05661_ VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13367_ _06839_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__clkbuf_1
X_10579_ net773 _03348_ _04768_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__mux2_1
X_15106_ clknet_leaf_102_clk _07130_ VGND VGND VPWR VPWR reg_out\[24\] sky130_fd_sc_hd__dfxtp_1
X_12318_ _06073_ _06075_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13298_ cpuregs\[18\]\[20\] _04860_ _06802_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__mux2_1
X_15037_ clknet_leaf_122_clk _00695_ VGND VGND VPWR VPWR count_cycle\[20\] sky130_fd_sc_hd__dfxtp_1
X_12249_ _02482_ _06009_ _05863_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07790_ _02237_ net213 VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_79_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15939_ clknet_leaf_51_clk _01511_ VGND VGND VPWR VPWR cpuregs\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_09460_ _03921_ _03922_ _03447_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__mux2_1
X_08411_ reg_next_pc\[9\] reg_out\[9\] _02949_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_35_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09391_ cpuregs\[0\]\[10\] cpuregs\[1\]\[10\] cpuregs\[2\]\[10\] cpuregs\[3\]\[10\]
+ _03456_ _03459_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_16_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08342_ _02251_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_62_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08273_ net220 net246 _02850_ _02757_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__o31a_1
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07224_ _01884_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_115_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07155_ _01822_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__inv_2
XFILLER_0_42_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_495 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07988_ _02603_ _02604_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09727_ _04152_ _04155_ _04153_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ decoded_imm\[19\] net181 VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_143_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _03124_ _03126_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09589_ _04042_ _04044_ _04047_ _03427_ _03490_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_600 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11620_ _05497_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11551_ _05435_ _05424_ _05420_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10502_ net1299 _03322_ _04731_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14270_ _01760_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__clkbuf_1
X_11482_ decoded_imm_j\[11\] _05212_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13221_ decoded_imm\[14\] _06752_ _06735_ _06759_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__o22a_1
X_10433_ _04696_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13152_ _06719_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__clkbuf_1
X_10364_ _04659_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__clkbuf_1
X_12103_ decoded_imm\[4\] _03158_ _01906_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__mux2_1
X_13083_ mem_state\[1\] _06682_ _06680_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__mux2_1
X_10295_ net1197 _03314_ _04622_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12034_ _01923_ _01926_ _05805_ _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__and4b_1
X_13985_ net1239 _06941_ _01602_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15724_ clknet_leaf_154_clk _01299_ VGND VGND VPWR VPWR cpuregs\[22\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12936_ decoded_imm_j\[13\] _01075_ _03169_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15655_ clknet_leaf_55_clk _01230_ VGND VGND VPWR VPWR cpuregs\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12867_ _06544_ _06559_ net242 _06553_ net548 VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11818_ count_cycle\[28\] count_cycle\[29\] _05655_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__and3_1
X_14606_ clknet_leaf_44_clk _00264_ VGND VGND VPWR VPWR cpuregs\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15586_ clknet_leaf_37_clk _01161_ VGND VGND VPWR VPWR cpuregs\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12798_ instr_lui _06513_ _06519_ _06523_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14537_ clknet_leaf_21_clk _00195_ VGND VGND VPWR VPWR cpuregs\[13\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11749_ _05609_ _05610_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_677 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14468_ clknet_leaf_138_clk _00126_ VGND VGND VPWR VPWR cpuregs\[12\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13419_ cpuregs\[24\]\[13\] _04846_ _06863_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__mux2_1
Xpicorv32_302 VGND VGND VPWR VPWR picorv32_302/HI pcpi_insn[12] sky130_fd_sc_hd__conb_1
X_14399_ clknet_leaf_136_clk _00062_ VGND VGND VPWR VPWR cpuregs\[11\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xpicorv32_313 VGND VGND VPWR VPWR picorv32_313/HI pcpi_insn[23] sky130_fd_sc_hd__conb_1
XFILLER_0_24_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_324 VGND VGND VPWR VPWR picorv32_324/HI trace_data[1] sky130_fd_sc_hd__conb_1
Xpicorv32_335 VGND VGND VPWR VPWR picorv32_335/HI trace_data[12] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_346 VGND VGND VPWR VPWR picorv32_346/HI trace_data[23] sky130_fd_sc_hd__conb_1
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpicorv32_357 VGND VGND VPWR VPWR picorv32_357/HI trace_data[34] sky130_fd_sc_hd__conb_1
XFILLER_0_12_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08960_ _00014_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07911_ _02125_ _02475_ _02488_ _02524_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__o221a_1
X_08891_ reg_out\[29\] alu_out_q\[29\] _03176_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07842_ net209 VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__inv_2
X_07773_ net252 net227 VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09512_ cpuregs\[24\]\[14\] cpuregs\[25\]\[14\] cpuregs\[26\]\[14\] cpuregs\[27\]\[14\]
+ _03640_ _03496_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_108_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09443_ _02200_ net243 VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09374_ _02099_ net243 VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_121_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08325_ _02912_ _02913_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_74_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08256_ net246 _02851_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_50_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07207_ _01871_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__buf_4
X_08187_ _02413_ _02781_ _02788_ _02585_ VGND VGND VPWR VPWR alu_out\[18\] sky130_fd_sc_hd__a22o_1
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10080_ _04506_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13770_ net1218 _06931_ _07064_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__mux2_1
X_10982_ cpuregs\[17\]\[7\] _04833_ _04995_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12721_ cpuregs\[0\]\[30\] cpuregs\[1\]\[30\] cpuregs\[2\]\[30\] cpuregs\[3\]\[30\]
+ _05819_ _03086_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_27_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15440_ clknet_leaf_46_clk _01030_ VGND VGND VPWR VPWR cpuregs\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12652_ cpuregs\[6\]\[27\] cpuregs\[7\]\[27\] _03084_ VGND VGND VPWR VPWR _06395_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ decoded_imm_j\[17\] _05228_ _05464_ _05452_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__a31o_1
X_15371_ clknet_leaf_93_clk _00961_ VGND VGND VPWR VPWR latched_rd\[1\] sky130_fd_sc_hd__dfxtp_1
X_12583_ cpuregs\[4\]\[24\] cpuregs\[5\]\[24\] cpuregs\[6\]\[24\] cpuregs\[7\]\[24\]
+ _05908_ _06156_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14322_ _01787_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_340 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_52_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11534_ decoded_imm_j\[15\] _05222_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14253_ net616 VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__clkbuf_1
X_11465_ _05355_ _05356_ _05193_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13204_ decoded_imm\[22\] _06740_ _06737_ _06750_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__o22a_1
XFILLER_0_151_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10416_ _04687_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14184_ _01716_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_36_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11396_ _05276_ _05281_ _05292_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__a21bo_1
X_13135_ net150 net112 _06707_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__mux2_1
X_10347_ _04650_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13066_ is_alu_reg_imm _06513_ _06524_ _06629_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__a22o_1
X_10278_ cpuregs\[2\]\[12\] _03263_ _04611_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12017_ _05795_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13968_ _01601_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__buf_6
XFILLER_0_159_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15707_ clknet_leaf_134_clk _01282_ VGND VGND VPWR VPWR cpuregs\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12919_ _06594_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13899_ _04485_ _01564_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__nor2_4
X_15638_ clknet_leaf_146_clk _01213_ VGND VGND VPWR VPWR cpuregs\[23\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15569_ clknet_leaf_16_clk _01144_ VGND VGND VPWR VPWR cpuregs\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_127_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08110_ _02471_ _02716_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09090_ cpuregs\[16\]\[2\] cpuregs\[17\]\[2\] cpuregs\[18\]\[2\] cpuregs\[19\]\[2\]
+ _03554_ _03459_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__mux4_1
XFILLER_0_141_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08041_ _02585_ _02650_ _02653_ VGND VGND VPWR VPWR alu_out\[7\] sky130_fd_sc_hd__a21o_1
XFILLER_0_153_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold902 cpuregs\[29\]\[3\] VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 cpuregs\[25\]\[3\] VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold924 net159 VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold935 cpuregs\[8\]\[1\] VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 cpuregs\[14\]\[3\] VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 cpuregs\[5\]\[6\] VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 cpuregs\[29\]\[23\] VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _03807_ _04437_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__or2_1
Xhold979 cpuregs\[4\]\[18\] VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_4_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08874_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07825_ net194 net226 VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_511 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07756_ _02365_ _02367_ _02364_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_123_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07687_ _02302_ _02304_ _02312_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__o21ai_1
X_09426_ _02177_ _03770_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09357_ _03475_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_830 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_81_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08308_ _02440_ _02569_ _02898_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ cpuregs\[28\]\[7\] cpuregs\[29\]\[7\] cpuregs\[30\]\[7\] cpuregs\[31\]\[7\]
+ _03640_ _03492_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08239_ _02757_ _02835_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11250_ _05181_ _05182_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_132_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10201_ net1152 _03235_ _04564_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__mux2_1
X_11181_ count_instr\[41\] net1418 VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10132_ _04535_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14940_ clknet_leaf_120_clk _00598_ VGND VGND VPWR VPWR count_instr\[49\] sky130_fd_sc_hd__dfxtp_1
X_10063_ _04497_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14871_ clknet_leaf_151_clk _00529_ VGND VGND VPWR VPWR cpuregs\[17\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_13822_ net670 _06983_ _07086_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_98_875 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13753_ _07058_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__clkbuf_1
X_10965_ _04993_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12704_ _06177_ _06440_ _06442_ _06444_ _06164_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_39_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13684_ cpuregs\[23\]\[27\] _06981_ _07014_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10896_ net671 _04883_ _04922_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__mux2_1
X_12635_ _05969_ _06378_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__or2_1
X_15423_ clknet_leaf_158_clk _01013_ VGND VGND VPWR VPWR cpuregs\[18\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15354_ clknet_leaf_68_clk _00944_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dfxtp_1
X_12566_ cpuregs\[12\]\[23\] cpuregs\[13\]\[23\] cpuregs\[14\]\[23\] cpuregs\[15\]\[23\]
+ _03133_ _03134_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11517_ _05402_ _05403_ _05404_ _05217_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__o2bb2a_1
X_14305_ net841 _03178_ _01778_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15285_ clknet_leaf_92_clk _00878_ VGND VGND VPWR VPWR decoded_imm_j\[3\] sky130_fd_sc_hd__dfxtp_2
X_12497_ _06245_ _06246_ _06014_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold209 cpuregs\[0\]\[10\] VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ _01743_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__clkbuf_1
X_11448_ _05289_ _05336_ _05337_ _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_516 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14167_ net1377 _06987_ _01673_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11379_ decoded_imm_j\[3\] _05195_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__or2_1
X_13118_ net141 net103 _06696_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__mux2_1
X_14098_ _01670_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13049_ _06662_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_53_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07610_ _02198_ _02210_ _02241_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__or3_1
X_08590_ cpuregs\[16\]\[3\] cpuregs\[17\]\[3\] cpuregs\[18\]\[3\] cpuregs\[19\]\[3\]
+ _03107_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_105_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07541_ latched_is_lb latched_is_lh VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_88_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_238 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07472_ _02083_ _02113_ _02085_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09211_ cpuregs\[12\]\[5\] cpuregs\[13\]\[5\] cpuregs\[14\]\[5\] cpuregs\[15\]\[5\]
+ _03680_ _03443_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_102 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_57_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09142_ _03613_ _03611_ _03610_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_658 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09073_ _02044_ _03480_ _03074_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__a21o_1
X_08024_ _02625_ _02637_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold710 count_cycle\[23\] VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_114_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold721 cpuregs\[30\]\[21\] VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold732 cpuregs\[26\]\[29\] VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 cpuregs\[3\]\[6\] VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 count_instr\[14\] VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold765 cpuregs\[31\]\[22\] VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 cpuregs\[15\]\[19\] VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 cpuregs\[1\]\[31\] VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 cpuregs\[9\]\[23\] VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _03474_ _04412_ _04421_ _03528_ reg_pc\[28\] VGND VGND VPWR VPWR _04422_
+ sky130_fd_sc_hd__a32o_1
X_08926_ _03400_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_71_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08857_ _03336_ _03339_ _03293_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07808_ net188 net220 VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _03278_ _03279_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__nor2_1
X_07739_ count_instr\[29\] _01965_ count_cycle\[61\] _02055_ VGND VGND VPWR VPWR _02362_
+ sky130_fd_sc_hd__a22o_1
X_10750_ cpuregs\[26\]\[28\] _04877_ _04861_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09409_ _03437_ _03872_ _03419_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_912 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_80_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10681_ _03220_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12420_ _06167_ _06169_ _06171_ _06173_ _06151_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__a221o_2
X_12351_ _05871_ _06106_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11302_ _01872_ _05219_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_460 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15070_ clknet_leaf_119_clk _00728_ VGND VGND VPWR VPWR count_cycle\[53\] sky130_fd_sc_hd__dfxtp_1
X_12282_ _05879_ _06036_ _06038_ _06040_ _03104_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__a221o_2
XFILLER_0_133_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ cpuregs\[5\]\[25\] _06977_ _01624_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__mux2_1
X_11233_ net499 net369 _05141_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11164_ count_instr\[36\] _05119_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__nand2_1
X_10115_ net1326 _03179_ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__mux2_1
X_11095_ count_instr\[15\] count_instr\[14\] _05072_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__and3_1
X_14923_ clknet_leaf_116_clk _00581_ VGND VGND VPWR VPWR count_instr\[32\] sky130_fd_sc_hd__dfxtp_1
X_10046_ net862 _03189_ _04487_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__mux2_1
Xhold70 instr_add VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 instr_addi VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 count_cycle\[33\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ clknet_leaf_127_clk _00512_ VGND VGND VPWR VPWR cpuregs\[20\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_13805_ _07063_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14785_ clknet_leaf_148_clk _00443_ VGND VGND VPWR VPWR cpuregs\[16\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_11997_ _05766_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_683 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_86_834 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_133_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13736_ _07049_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__clkbuf_1
X_10948_ cpuregs\[20\]\[23\] _04867_ _04981_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_119_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13667_ net737 _06964_ _07003_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_923 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10879_ _04948_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_777 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15406_ clknet_leaf_64_clk _00996_ VGND VGND VPWR VPWR decoded_imm\[2\] sky130_fd_sc_hd__dfxtp_2
X_12618_ _06073_ _06362_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__or2_1
X_13598_ _06972_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15337_ clknet_leaf_69_clk _00927_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dfxtp_1
X_12549_ cpuregs\[31\]\[22\] _03092_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_1 _01566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15268_ clknet_leaf_86_clk _00861_ VGND VGND VPWR VPWR decoded_imm_j\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14219_ net1112 _06971_ _01732_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_128_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15199_ clknet_leaf_70_clk alu_out\[12\] VGND VGND VPWR VPWR alu_out_q\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09760_ decoded_imm\[22\] net185 VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__nand2_1
X_08711_ reg_out\[5\] alu_out_q\[5\] latched_stalu VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__mux2_1
X_09691_ _04079_ _04145_ _03075_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08642_ _01915_ _03122_ _03159_ _01944_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__o22a_1
Xrebuffer13 net396 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_1
Xrebuffer24 _02813_ VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_1
Xrebuffer35 net395 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_1
Xrebuffer46 net1418 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_1
X_08573_ _03091_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_157_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07524_ reg_pc\[13\] decoded_imm\[13\] VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_157_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07455_ _02096_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__xnor2_1
X_07386_ net28 net130 _02032_ _01940_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09125_ _03593_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_118_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_263 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09056_ net182 decoded_imm\[1\] VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__nor2_1
X_08007_ net250 _02609_ _02573_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold540 cpuregs\[2\]\[17\] VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 cpuregs\[31\]\[4\] VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_182 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold562 cpuregs\[4\]\[26\] VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 cpuregs\[23\]\[31\] VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 cpuregs\[29\]\[9\] VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold595 cpuregs\[13\]\[4\] VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__dlygate4sd3_1
X_09958_ cpuregs\[4\]\[28\] cpuregs\[5\]\[28\] cpuregs\[6\]\[28\] cpuregs\[7\]\[28\]
+ _03680_ _03443_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__mux4_1
X_08909_ _03383_ _03384_ _03199_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__mux2_2
X_09889_ _04273_ _04304_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__nand2_1
X_11920_ count_cycle\[60\] count_cycle\[61\] _05724_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11851_ net515 _05678_ _05647_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__o21ai_1
X_10802_ _04907_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__clkbuf_1
X_14570_ clknet_leaf_45_clk _00228_ VGND VGND VPWR VPWR cpuregs\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11782_ _05633_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10733_ _04866_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__clkbuf_1
X_13521_ _06920_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13452_ cpuregs\[24\]\[29\] _04879_ _06874_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__mux2_1
X_10664_ cpuregs\[26\]\[0\] _04817_ _04819_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_904 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12403_ cpuregs\[4\]\[16\] cpuregs\[5\]\[16\] cpuregs\[6\]\[16\] cpuregs\[7\]\[16\]
+ _06011_ _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13383_ _06847_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10595_ net963 _03179_ _04782_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12334_ cpuregs\[24\]\[13\] cpuregs\[25\]\[13\] cpuregs\[26\]\[13\] cpuregs\[27\]\[13\]
+ _05970_ _03108_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_756 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15122_ clknet_leaf_74_clk _00748_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15053_ clknet_leaf_114_clk _00711_ VGND VGND VPWR VPWR count_cycle\[36\] sky130_fd_sc_hd__dfxtp_1
X_12265_ _06023_ _06024_ _05927_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14004_ net801 _06960_ _01613_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__mux2_1
X_11216_ _05158_ _05159_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12196_ cpuregs\[4\]\[8\] cpuregs\[5\]\[8\] _03062_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__mux2_1
Xoutput60 net60 VGND VGND VPWR VPWR mem_addr[5] sky130_fd_sc_hd__clkbuf_4
Xoutput71 net71 VGND VGND VPWR VPWR mem_la_addr[15] sky130_fd_sc_hd__clkbuf_4
Xoutput82 net82 VGND VGND VPWR VPWR mem_la_addr[26] sky130_fd_sc_hd__buf_2
XFILLER_0_128_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xoutput93 net93 VGND VGND VPWR VPWR mem_la_addr[7] sky130_fd_sc_hd__clkbuf_4
X_11147_ count_instr\[31\] net377 _05036_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__a21oi_1
X_11078_ count_instr\[10\] _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__and2_1
X_15955_ clknet_leaf_5_clk _01527_ VGND VGND VPWR VPWR cpuregs\[10\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14906_ clknet_leaf_121_clk _00564_ VGND VGND VPWR VPWR count_instr\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10029_ cpuregs\[4\]\[30\] cpuregs\[5\]\[30\] cpuregs\[6\]\[30\] cpuregs\[7\]\[30\]
+ _03440_ _03451_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__mux4_1
X_15886_ clknet_leaf_15_clk _01458_ VGND VGND VPWR VPWR cpuregs\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_14837_ clknet_leaf_0_clk _00495_ VGND VGND VPWR VPWR cpuregs\[20\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14768_ clknet_leaf_27_clk _00426_ VGND VGND VPWR VPWR cpuregs\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13719_ net840 _06948_ _07039_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_906 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14699_ clknet_leaf_51_clk _00357_ VGND VGND VPWR VPWR cpuregs\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07240_ _00809_ _01899_ _01851_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07171_ _01833_ _01834_ _01835_ _01836_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__or4_1
XFILLER_0_143_246 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_6_669 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_131_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_631 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09812_ _02277_ _03660_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__and2_1
X_09743_ _03446_ _04196_ _03417_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09674_ _03557_ _04129_ _03425_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08625_ _03037_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__buf_6
XFILLER_0_49_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _03075_ _01896_ reg_sh\[2\] VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07507_ count_instr\[45\] _02052_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__and2_1
X_08487_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_714 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07438_ net201 VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_45_572 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_91_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07369_ cpu_state\[3\] cpu_state\[6\] _01953_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__or3_4
XFILLER_0_134_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09108_ _03577_ _03578_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_542 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10380_ _04667_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09039_ cpuregs\[0\]\[1\] cpuregs\[1\]\[1\] cpuregs\[2\]\[1\] cpuregs\[3\]\[1\] _03406_
+ _03410_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__mux4_1
X_12050_ cpuregs\[0\]\[0\] cpuregs\[1\]\[0\] cpuregs\[2\]\[0\] cpuregs\[3\]\[0\] _05819_
+ _03086_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__mux4_1
Xhold370 cpuregs\[21\]\[31\] VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 net146 VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 cpuregs\[30\]\[28\] VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net980 _04852_ _05006_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ clknet_leaf_130_clk _01315_ VGND VGND VPWR VPWR cpuregs\[22\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12952_ net433 _01070_ _06587_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11903_ count_cycle\[55\] count_cycle\[56\] _05714_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__and3_1
X_15671_ clknet_leaf_128_clk _01246_ VGND VGND VPWR VPWR cpuregs\[29\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_210 _03193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12883_ net547 _06541_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__and2_1
*XANTENNA_221 _06182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
*XANTENNA_232 _03581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14622_ clknet_leaf_147_clk _00280_ VGND VGND VPWR VPWR cpuregs\[21\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ net1404 net366 _05622_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_349 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11765_ _05620_ _05621_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__nor2_1
X_14553_ clknet_leaf_9_clk _00211_ VGND VGND VPWR VPWR cpuregs\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_138_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10716_ net1301 _04854_ _04840_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__mux2_1
X_13504_ net1235 _04863_ _06910_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__mux2_1
X_14484_ clknet_leaf_1_clk _00142_ VGND VGND VPWR VPWR cpuregs\[30\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11696_ _05185_ _05567_ _05568_ _05257_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__o211a_1
X_13435_ _06875_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10647_ net1081 _03348_ _04804_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xrebuffer4 _05661_ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13366_ net1202 _04860_ _06838_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10578_ _04773_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_482 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_11_417 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15105_ clknet_leaf_102_clk _07129_ VGND VGND VPWR VPWR reg_out\[23\] sky130_fd_sc_hd__dfxtp_1
X_12317_ cpuregs\[24\]\[12\] cpuregs\[25\]\[12\] cpuregs\[26\]\[12\] cpuregs\[27\]\[12\]
+ _06074_ _05932_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__mux4_1
X_13297_ _06779_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__buf_4
X_15036_ clknet_leaf_122_clk _00694_ VGND VGND VPWR VPWR count_cycle\[19\] sky130_fd_sc_hd__dfxtp_1
X_12248_ _05901_ _05999_ _06008_ _05904_ decoded_imm\[9\] VGND VGND VPWR VPWR _06009_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_139_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12179_ _05912_ _05941_ _03123_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15938_ clknet_leaf_52_clk _01510_ VGND VGND VPWR VPWR cpuregs\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_64_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15869_ clknet_leaf_17_clk _01441_ VGND VGND VPWR VPWR cpuregs\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_817 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08410_ _02964_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_1
X_09390_ cpuregs\[4\]\[10\] cpuregs\[5\]\[10\] cpuregs\[6\]\[10\] cpuregs\[7\]\[10\]
+ _03554_ _03459_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_35_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08341_ _01940_ _02926_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__nand2_2
XFILLER_0_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_100 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_714 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08272_ _02429_ _02861_ _02866_ _02608_ VGND VGND VPWR VPWR alu_out\[25\] sky130_fd_sc_hd__a22o_2
XFILLER_0_144_511 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_509 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07223_ _01839_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07154_ _01820_ _01821_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07987_ net196 _02602_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__or2_1
X_09726_ _04177_ _04179_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ _02222_ _03624_ _04113_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_143_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_940 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_139_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08608_ cpuregs\[4\]\[4\] cpuregs\[5\]\[4\] cpuregs\[6\]\[4\] cpuregs\[7\]\[4\] _03091_
+ _03125_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__mux4_1
X_09588_ _04045_ _04046_ _03647_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08539_ cpuregs\[4\]\[2\] cpuregs\[5\]\[2\] cpuregs\[6\]\[2\] cpuregs\[7\]\[2\] _03051_
+ _03052_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11550_ _05421_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10501_ _04732_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11481_ decoded_imm_j\[11\] _05212_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__nor2_1
X_13220_ _06525_ decoded_imm_j\[14\] _06738_ _06532_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__a22o_1
X_10432_ cpuregs\[21\]\[20\] _03314_ _04695_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_791 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_122_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13151_ net1283 net121 _06684_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__mux2_1
X_10363_ net977 _03314_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__mux2_1
X_12102_ _02502_ _05863_ _05868_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13082_ _01821_ _06675_ _05763_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__a21oi_1
X_10294_ _04599_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12033_ mem_do_prefetch _03389_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13984_ _01610_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__clkbuf_1
X_15723_ clknet_leaf_0_clk _01298_ VGND VGND VPWR VPWR cpuregs\[22\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12935_ _06602_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__clkbuf_1
X_15654_ clknet_leaf_35_clk _01229_ VGND VGND VPWR VPWR cpuregs\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12866_ _06538_ _06559_ net242 _06553_ net602 VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__a32o_1
X_14605_ clknet_leaf_39_clk _00263_ VGND VGND VPWR VPWR cpuregs\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11817_ net509 net384 _05657_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__a21oi_1
X_15585_ clknet_leaf_24_clk _01160_ VGND VGND VPWR VPWR cpuregs\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12797_ _01068_ _01066_ _01067_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ clknet_leaf_59_clk _00194_ VGND VGND VPWR VPWR cpuregs\[13\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_99_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11748_ net779 _05607_ _05169_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14467_ clknet_leaf_98_clk _00125_ VGND VGND VPWR VPWR cpuregs\[12\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11679_ _05246_ _05552_ _05495_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13418_ _06866_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14398_ clknet_leaf_135_clk _00061_ VGND VGND VPWR VPWR cpuregs\[11\]\[24\] sky130_fd_sc_hd__dfxtp_1
Xpicorv32_303 VGND VGND VPWR VPWR picorv32_303/HI pcpi_insn[13] sky130_fd_sc_hd__conb_1
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_314 VGND VGND VPWR VPWR picorv32_314/HI pcpi_insn[24] sky130_fd_sc_hd__conb_1
Xpicorv32_325 VGND VGND VPWR VPWR picorv32_325/HI trace_data[2] sky130_fd_sc_hd__conb_1
XFILLER_0_12_737 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13349_ net1319 _04844_ _06827_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__mux2_1
Xpicorv32_336 VGND VGND VPWR VPWR picorv32_336/HI trace_data[13] sky130_fd_sc_hd__conb_1
XFILLER_0_59_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpicorv32_347 VGND VGND VPWR VPWR picorv32_347/HI trace_data[24] sky130_fd_sc_hd__conb_1
Xpicorv32_358 VGND VGND VPWR VPWR picorv32_358/HI trace_data[35] sky130_fd_sc_hd__conb_1
XFILLER_0_11_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15019_ clknet_leaf_111_clk _00677_ VGND VGND VPWR VPWR count_cycle\[2\] sky130_fd_sc_hd__dfxtp_2
X_07910_ _02486_ _02529_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__nand2_1
X_08890_ _03368_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_90_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07841_ _02425_ _02448_ _02446_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__a2bb2o_1
X_07772_ net252 net227 VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_160_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09511_ _03970_ _03971_ _03579_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09442_ _02154_ _03481_ _03904_ _03616_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09373_ _02044_ _03479_ _03837_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_314 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08324_ _02912_ _02913_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_615 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_7_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08255_ _02757_ _02850_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__and2_1
X_07206_ cpu_state\[1\] VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08186_ _02786_ _02787_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_350 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_772 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09709_ _03593_ _04163_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__or2_1
X_10981_ _05002_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12720_ _05925_ _06459_ _03037_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12651_ _05871_ _06393_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _05463_ _05473_ _05474_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15370_ clknet_leaf_93_clk _00960_ VGND VGND VPWR VPWR latched_rd\[0\] sky130_fd_sc_hd__dfxtp_1
X_12582_ _06328_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14321_ net861 _03234_ _01778_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__mux2_1
X_11533_ decoded_imm_j\[15\] _05222_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11464_ _05273_ _05339_ _05208_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__o21ba_1
X_14252_ _01751_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10415_ cpuregs\[21\]\[12\] _03263_ _04684_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__mux2_1
X_13203_ mem_rdata_q\[22\] _06742_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11395_ _05290_ _05291_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__and2_1
X_14183_ cpuregs\[8\]\[5\] _06935_ _01710_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13134_ _06710_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__clkbuf_1
X_10346_ cpuregs\[28\]\[12\] _03263_ _04647_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__mux2_1
X_13065_ _06670_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__clkbuf_1
X_10277_ _04613_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12016_ net854 net83 _05785_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap2 _02570_ VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__clkbuf_1
X_13967_ _04562_ _01564_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15706_ clknet_leaf_20_clk _01281_ VGND VGND VPWR VPWR cpuregs\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_100_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12918_ mem_rdata_q\[27\] net20 _06589_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_433 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_76_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13898_ latched_rd\[3\] latched_rd\[4\] latched_rd\[2\] VGND VGND VPWR VPWR _01564_
+ sky130_fd_sc_hd__or3b_4
X_15637_ clknet_leaf_146_clk _01212_ VGND VGND VPWR VPWR cpuregs\[23\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12849_ net529 _06554_ _06545_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15568_ clknet_leaf_5_clk _01143_ VGND VGND VPWR VPWR cpuregs\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14519_ clknet_leaf_13_clk _00177_ VGND VGND VPWR VPWR cpuregs\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15499_ clknet_leaf_92_clk _01084_ VGND VGND VPWR VPWR mem_rdata_q\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_119 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08040_ _02066_ _02489_ _02651_ _02652_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold903 cpuregs\[10\]\[14\] VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 cpuregs\[22\]\[10\] VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 cpuregs\[5\]\[18\] VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold936 cpuregs\[18\]\[31\] VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_95 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_141_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold947 cpuregs\[12\]\[12\] VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold958 cpuregs\[1\]\[2\] VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ cpuregs\[20\]\[29\] cpuregs\[21\]\[29\] cpuregs\[22\]\[29\] cpuregs\[23\]\[29\]
+ _03438_ _03812_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__mux4_1
Xhold969 cpuregs\[29\]\[19\] VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__dlygate4sd3_1
X_08942_ _00015_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_4_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08873_ _03261_ _03350_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__o21a_2
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07824_ net194 net226 VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07755_ _02375_ _02376_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_123_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07686_ _02302_ _02304_ _02312_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09425_ _02139_ _03481_ _03888_ _03670_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09356_ _03473_ _03811_ _03821_ _03526_ reg_pc\[9\] VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_23_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_842 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08307_ _02369_ net224 _02618_ _02641_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09287_ _03581_ _03754_ _03426_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08238_ net217 net216 _02813_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_138_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08169_ _02213_ _02770_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__nor2_1
X_10200_ _04572_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11180_ net406 _05134_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10131_ cpuregs\[30\]\[8\] _03235_ _04526_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10062_ net1164 _03241_ _04487_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14870_ clknet_leaf_158_clk _00528_ VGND VGND VPWR VPWR cpuregs\[17\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_13821_ _07094_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13752_ cpuregs\[29\]\[27\] _06981_ _07050_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__mux2_1
X_10964_ net881 _04883_ _04958_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12703_ _05969_ _06443_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13683_ _07021_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__clkbuf_1
X_10895_ _04956_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15422_ clknet_leaf_152_clk _01012_ VGND VGND VPWR VPWR cpuregs\[18\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_12634_ cpuregs\[24\]\[26\] cpuregs\[25\]\[26\] cpuregs\[26\]\[26\] cpuregs\[27\]\[26\]
+ _05970_ _03108_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15353_ clknet_leaf_69_clk _00943_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_648 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12565_ _06310_ _06311_ _06014_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14304_ _01777_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_374 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11516_ _05273_ _05388_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15284_ clknet_leaf_92_clk _00877_ VGND VGND VPWR VPWR decoded_imm_j\[2\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_123_322 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12496_ cpuregs\[0\]\[20\] cpuregs\[1\]\[20\] cpuregs\[2\]\[20\] cpuregs\[3\]\[20\]
+ _06055_ _05829_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14235_ net1132 _06987_ _01709_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11447_ _05206_ _05327_ _05339_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_74_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14166_ _01706_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__clkbuf_1
X_11378_ decoded_imm_j\[3\] _05195_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__nand2_1
X_13117_ _06701_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__clkbuf_1
X_10329_ net1289 _03209_ _04636_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__mux2_1
X_14097_ cpuregs\[6\]\[29\] _06985_ _01660_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__mux2_1
X_13048_ net1005 _04867_ _06658_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14999_ clknet_leaf_87_clk _00657_ VGND VGND VPWR VPWR reg_next_pc\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07540_ net177 VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__buf_4
XFILLER_0_159_753 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07471_ _01846_ _01913_ net19 net2 _01933_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_85_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09210_ _03587_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__buf_8
XFILLER_0_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09141_ decoded_imm\[3\] _01992_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_114 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_133_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09072_ _03482_ _03544_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_115_867 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08023_ _02612_ _02615_ _02624_ _02636_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__a211o_1
Xhold700 cpuregs\[15\]\[28\] VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold711 cpuregs\[27\]\[2\] VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold722 cpuregs\[15\]\[25\] VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 cpuregs\[31\]\[20\] VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 cpuregs\[27\]\[15\] VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 cpuregs\[31\]\[15\] VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 cpuregs\[3\]\[26\] VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 cpuregs\[15\]\[1\] VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 cpuregs\[25\]\[23\] VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 cpuregs\[4\]\[23\] VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _04414_ _04416_ _04418_ _04420_ _03431_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_572 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08925_ _00014_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08856_ _03337_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__nor2_1
X_07807_ net189 net221 VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__nand2_1
X_08787_ reg_pc\[15\] _03272_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ count_instr\[61\] _02052_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07669_ _02262_ _02271_ _02287_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09408_ cpuregs\[8\]\[11\] cpuregs\[9\]\[11\] cpuregs\[10\]\[11\] cpuregs\[11\]\[11\]
+ _03440_ _03451_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__mux4_1
X_10680_ _04830_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09339_ cpuregs\[8\]\[9\] cpuregs\[9\]\[9\] cpuregs\[10\]\[9\] cpuregs\[11\]\[9\]
+ _03586_ _03449_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_90_551 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12350_ cpuregs\[4\]\[14\] cpuregs\[5\]\[14\] _03062_ VGND VGND VPWR VPWR _06106_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11301_ reg_next_pc\[14\] _03270_ _02946_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__mux2_1
X_12281_ _03106_ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11232_ _05168_ _05170_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__nor2_1
X_14020_ _01629_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11163_ count_instr\[36\] _05119_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10114_ _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__clkbuf_8
X_11094_ _05073_ _05074_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__nor2_1
X_14922_ clknet_leaf_117_clk _00580_ VGND VGND VPWR VPWR count_instr\[31\] sky130_fd_sc_hd__dfxtp_1
X_10045_ _04488_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_1
Xhold60 mem_rdata[19] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 net25 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 instr_sra VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ clknet_leaf_144_clk _00511_ VGND VGND VPWR VPWR cpuregs\[20\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold93 reg_next_pc\[24\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ _07085_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__clkbuf_1
X_14784_ clknet_leaf_148_clk _00442_ VGND VGND VPWR VPWR cpuregs\[16\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11996_ _05784_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13735_ net1328 _06964_ _07039_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_846 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_133_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_701 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10947_ _04984_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13666_ _07012_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10878_ net884 _04865_ _04945_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_935 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15405_ clknet_leaf_64_clk _00995_ VGND VGND VPWR VPWR decoded_imm\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_156_789 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12617_ cpuregs\[24\]\[25\] cpuregs\[25\]\[25\] cpuregs\[26\]\[25\] cpuregs\[27\]\[25\]
+ _06074_ _03151_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_306 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13597_ net1124 _06971_ _06967_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_14_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15336_ clknet_leaf_69_clk _00926_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dfxtp_2
X_12548_ _05969_ _06295_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_491 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15267_ clknet_leaf_87_clk _00860_ VGND VGND VPWR VPWR decoded_imm_j\[10\] sky130_fd_sc_hd__dfxtp_1
X_12479_ _06058_ _06229_ _06182_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__o21a_1
*XANTENNA_2 _01638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14218_ _01734_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15198_ clknet_leaf_70_clk alu_out\[11\] VGND VGND VPWR VPWR alu_out_q\[11\] sky130_fd_sc_hd__dfxtp_2
X_14149_ cpuregs\[7\]\[21\] _06969_ _01696_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08710_ reg_pc\[5\] _03206_ _03199_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__o21ai_1
X_09690_ _02237_ _03619_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08641_ _03158_ decoded_imm_j\[4\] is_slli_srli_srai VGND VGND VPWR VPWR _03159_
+ sky130_fd_sc_hd__mux2_1
Xrebuffer14 _05127_ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer25 _05655_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_1
Xrebuffer36 _05667_ VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkbuf_1
Xrebuffer47 _05132_ VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08572_ _03038_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__buf_8
XFILLER_0_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07523_ _02159_ _02160_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_157_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07454_ _02074_ _02079_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07385_ net14 _01937_ _02031_ _01935_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_540 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09124_ cpuregs\[20\]\[3\] cpuregs\[21\]\[3\] cpuregs\[22\]\[3\] cpuregs\[23\]\[3\]
+ _03594_ _03595_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_118_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09055_ _01844_ decoded_imm\[1\] VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08006_ _02613_ _02616_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__nand2_1
Xhold530 cpuregs\[11\]\[28\] VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold541 cpuregs\[31\]\[11\] VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 cpuregs\[6\]\[24\] VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 cpuregs\[12\]\[2\] VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 reg_next_pc\[23\] VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold585 cpuregs\[5\]\[16\] VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 cpuregs\[11\]\[24\] VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ _01977_ _04393_ _04394_ _03397_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_51_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ reg_pc\[31\] _03377_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__xnor2_1
X_09888_ decoded_imm\[26\] net189 VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__xor2_2
X_08839_ reg_out\[22\] alu_out_q\[22\] _03175_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__mux2_1
X_11850_ count_cycle\[37\] count_cycle\[38\] count_cycle\[39\] _05673_ VGND VGND VPWR
+ VPWR _05680_ sky130_fd_sc_hd__and4_1
X_10801_ net775 _04856_ _04898_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__mux2_1
X_11781_ _05631_ _05625_ _05632_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_49_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_712 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13520_ net728 _04879_ _06910_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__mux2_1
X_10732_ net983 _04865_ _04861_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13451_ _06883_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10663_ _04818_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_242 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_24_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12402_ _03047_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_11_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13382_ cpuregs\[19\]\[28\] _04877_ _06838_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10594_ _04781_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__buf_6
XFILLER_0_24_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15121_ clknet_leaf_74_clk _00747_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12333_ _03142_ _06085_ _06089_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15052_ clknet_leaf_115_clk _00710_ VGND VGND VPWR VPWR count_cycle\[35\] sky130_fd_sc_hd__dfxtp_1
X_12264_ cpuregs\[16\]\[10\] cpuregs\[17\]\[10\] cpuregs\[18\]\[10\] cpuregs\[19\]\[10\]
+ _05948_ _05925_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__mux4_1
X_14003_ _01620_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__clkbuf_1
X_11215_ net758 _05156_ _05133_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__o21ai_1
X_12195_ _05957_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__clkbuf_1
Xoutput50 net50 VGND VGND VPWR VPWR mem_addr[25] sky130_fd_sc_hd__buf_2
XFILLER_0_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput61 net61 VGND VGND VPWR VPWR mem_addr[6] sky130_fd_sc_hd__clkbuf_4
Xoutput72 net72 VGND VGND VPWR VPWR mem_la_addr[16] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11146_ _05109_ _05110_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__nor2_1
Xoutput83 net83 VGND VGND VPWR VPWR mem_la_addr[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput94 net94 VGND VGND VPWR VPWR mem_la_addr[8] sky130_fd_sc_hd__clkbuf_4
X_11077_ _05060_ _05058_ _05062_ _05052_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__a211oi_1
X_15954_ clknet_leaf_15_clk _01526_ VGND VGND VPWR VPWR cpuregs\[10\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_14905_ clknet_leaf_121_clk _00563_ VGND VGND VPWR VPWR count_instr\[14\] sky130_fd_sc_hd__dfxtp_1
X_10028_ _03500_ _04472_ _03468_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_69_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ clknet_leaf_8_clk _01457_ VGND VGND VPWR VPWR cpuregs\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14836_ clknet_leaf_2_clk _00494_ VGND VGND VPWR VPWR cpuregs\[20\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_492 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_59_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14767_ clknet_leaf_42_clk _00425_ VGND VGND VPWR VPWR cpuregs\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11979_ net64 net95 _05774_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13718_ _07040_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_315 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14698_ clknet_leaf_54_clk _00356_ VGND VGND VPWR VPWR cpuregs\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13649_ cpuregs\[23\]\[10\] _06945_ _07003_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07170_ instr_sltiu instr_slti instr_bgeu instr_bge VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15319_ clknet_leaf_145_clk _00909_ VGND VGND VPWR VPWR cpuregs\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_120_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_120_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09811_ _03488_ _04262_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__and2_1
X_09742_ cpuregs\[28\]\[21\] cpuregs\[29\]\[21\] cpuregs\[30\]\[21\] cpuregs\[31\]\[21\]
+ _03586_ _03441_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__mux4_1
X_09673_ cpuregs\[16\]\[19\] cpuregs\[17\]\[19\] cpuregs\[18\]\[19\] cpuregs\[19\]\[19\]
+ _03456_ _03441_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08624_ _00011_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_38_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _03074_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__clkbuf_4
X_07506_ _01970_ _02137_ _02138_ _02145_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__a31o_1
XFILLER_0_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08486_ _01857_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__buf_4
X_07437_ _02075_ _02076_ _02080_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07368_ count_instr\[36\] _02013_ count_cycle\[4\] _01951_ _02015_ VGND VGND VPWR
+ VPWR _02016_ sky130_fd_sc_hd__a221o_2
XFILLER_0_45_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09107_ _03552_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_150_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_111_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_111_clk sky130_fd_sc_hd__clkbuf_2
X_07299_ _01950_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_554 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_32_256 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_102_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_180 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09038_ _03493_ _03511_ _03415_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold360 decoded_imm_j\[5\] VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 cpuregs\[25\]\[28\] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 cpuregs\[27\]\[26\] VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _05012_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__clkbuf_1
Xhold393 cpuregs\[12\]\[26\] VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12951_ _06610_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__clkbuf_1
X_11902_ net562 _05714_ _05715_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__a21oi_1
X_15670_ clknet_leaf_145_clk _01245_ VGND VGND VPWR VPWR cpuregs\[29\]\[23\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_200 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12882_ _05041_ _06548_ _06568_ _06529_ net464 VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__a32o_1
*XANTENNA_211 _03193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_222 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14621_ clknet_leaf_155_clk _00279_ VGND VGND VPWR VPWR cpuregs\[21\]\[19\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_233 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11833_ net451 _05664_ _05668_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ clknet_leaf_142_clk _00210_ VGND VGND VPWR VPWR cpuregs\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ net558 _05617_ _05169_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13503_ _06911_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10715_ _03294_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__clkbuf_4
X_14483_ clknet_leaf_32_clk _00141_ VGND VGND VPWR VPWR cpuregs\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11695_ _05031_ net1361 VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13434_ net1350 _04860_ _06874_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10646_ _04809_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer5 _05661_ VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13365_ _06815_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_102_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_102_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10577_ net771 _03341_ _04768_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15104_ clknet_leaf_102_clk _07128_ VGND VGND VPWR VPWR reg_out\[22\] sky130_fd_sc_hd__dfxtp_1
X_12316_ _03046_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_494 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_16084_ net126 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
X_13296_ _06801_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15035_ clknet_leaf_122_clk _00693_ VGND VGND VPWR VPWR count_cycle\[18\] sky130_fd_sc_hd__dfxtp_1
X_12247_ _06001_ _06003_ _06005_ _06007_ _03080_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12178_ cpuregs\[12\]\[7\] cpuregs\[13\]\[7\] cpuregs\[14\]\[7\] cpuregs\[15\]\[7\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__mux4_1
X_11129_ net1412 _05095_ net480 VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15937_ clknet_leaf_20_clk _01509_ VGND VGND VPWR VPWR cpuregs\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15868_ clknet_leaf_142_clk _01440_ VGND VGND VPWR VPWR cpuregs\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_14819_ clknet_leaf_124_clk _00477_ VGND VGND VPWR VPWR cpuregs\[25\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15799_ clknet_leaf_133_clk _01374_ VGND VGND VPWR VPWR cpuregs\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08340_ _01847_ _01913_ _01846_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08271_ _02864_ _02865_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_214 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07222_ _01883_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07153_ mem_do_wdata _01817_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07986_ net196 _02602_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__and2_1
X_09725_ _04178_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__inv_2
X_09656_ _03488_ _04090_ _04094_ _04112_ _03665_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_2_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _03039_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09587_ cpuregs\[0\]\[16\] cpuregs\[1\]\[16\] cpuregs\[2\]\[16\] cpuregs\[3\]\[16\]
+ _03440_ _03451_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_46_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ decoded_imm_j\[3\] decoded_imm_j\[2\] decoded_imm_j\[1\] _03057_ VGND VGND
+ VPWR VPWR _03058_ sky130_fd_sc_hd__or4_4
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_146_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08469_ _02331_ _03005_ _02993_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10500_ net1074 _03314_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11480_ _05263_ net1043 _05358_ _05369_ _05370_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_123_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10431_ _04672_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__buf_4
XFILLER_0_122_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13150_ _06718_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10362_ _04635_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__buf_4
X_12101_ _01906_ _03119_ _05867_ _01841_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__a211o_1
XFILLER_0_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10293_ _04621_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__clkbuf_1
X_13081_ _06681_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__clkbuf_1
X_12032_ _01871_ _01902_ _03389_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__or3_1
Xhold190 count_instr\[52\] VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_155_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13983_ net1169 _06939_ _01602_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__mux2_1
X_15722_ clknet_leaf_0_clk _01297_ VGND VGND VPWR VPWR cpuregs\[22\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12934_ decoded_imm_j\[12\] _01074_ _03169_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15653_ clknet_leaf_33_clk _01228_ VGND VGND VPWR VPWR cpuregs\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12865_ mem_rdata_q\[31\] mem_rdata_q\[30\] mem_rdata_q\[29\] _06563_ VGND VGND VPWR
+ VPWR _06564_ sky130_fd_sc_hd__nor4_1
XFILLER_0_68_440 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_157_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14604_ clknet_leaf_28_clk _00262_ VGND VGND VPWR VPWR cpuregs\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11816_ net1410 net378 _05622_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__o21ai_1
X_15584_ clknet_leaf_45_clk _01159_ VGND VGND VPWR VPWR cpuregs\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12796_ _06522_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_157_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14535_ clknet_leaf_98_clk _00193_ VGND VGND VPWR VPWR cpuregs\[13\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_99_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11747_ count_cycle\[7\] _05607_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14466_ clknet_leaf_136_clk _00124_ VGND VGND VPWR VPWR cpuregs\[12\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11678_ reg_next_pc\[26\] _02999_ _05248_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__a21o_1
X_13417_ cpuregs\[24\]\[12\] _04844_ _06863_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__mux2_1
X_10629_ _04800_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14397_ clknet_leaf_139_clk _00060_ VGND VGND VPWR VPWR cpuregs\[11\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xpicorv32_304 VGND VGND VPWR VPWR picorv32_304/HI pcpi_insn[14] sky130_fd_sc_hd__conb_1
X_13348_ _06829_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__clkbuf_1
Xpicorv32_315 VGND VGND VPWR VPWR picorv32_315/HI pcpi_insn[25] sky130_fd_sc_hd__conb_1
Xpicorv32_326 VGND VGND VPWR VPWR picorv32_326/HI trace_data[3] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpicorv32_337 VGND VGND VPWR VPWR picorv32_337/HI trace_data[14] sky130_fd_sc_hd__conb_1
Xpicorv32_348 VGND VGND VPWR VPWR picorv32_348/HI trace_data[25] sky130_fd_sc_hd__conb_1
Xpicorv32_359 VGND VGND VPWR VPWR picorv32_359/HI trace_valid sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_110_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13279_ cpuregs\[18\]\[11\] _04842_ _06791_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15018_ clknet_leaf_111_clk _00676_ VGND VGND VPWR VPWR count_cycle\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_75_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07840_ _02449_ net224 _02443_ _02457_ _02459_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07771_ _02385_ _02388_ _02391_ _01970_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09510_ cpuregs\[16\]\[14\] cpuregs\[17\]\[14\] cpuregs\[18\]\[14\] cpuregs\[19\]\[14\]
+ _03719_ _03450_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_160_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09441_ _02125_ net243 VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_125_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09372_ _02165_ net243 VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_432 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08323_ _02902_ _02906_ _02904_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_627 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08254_ net218 _02835_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07205_ _01869_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08185_ _02762_ _02766_ _02771_ _02772_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_537 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07969_ net119 _02586_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__xnor2_1
X_09708_ cpuregs\[28\]\[20\] cpuregs\[29\]\[20\] cpuregs\[30\]\[20\] cpuregs\[31\]\[20\]
+ _03463_ _03460_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__mux4_1
X_10980_ cpuregs\[17\]\[6\] _04831_ _04995_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09639_ cpuregs\[16\]\[18\] cpuregs\[17\]\[18\] cpuregs\[18\]\[18\] cpuregs\[19\]\[18\]
+ _03587_ _03442_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__mux4_1
X_12650_ cpuregs\[4\]\[27\] cpuregs\[5\]\[27\] _03051_ VGND VGND VPWR VPWR _06393_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ decoded_imm_j\[20\] _05237_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_26_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12581_ net218 _06327_ _06282_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14320_ _01786_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11532_ _05193_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ net610 VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11463_ _05269_ _05344_ _05354_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13202_ decoded_imm\[23\] _06740_ _06737_ _06749_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__o22a_1
X_10414_ _04686_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14182_ _01715_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__clkbuf_1
X_11394_ decoded_imm_j\[4\] _05197_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_59_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_389 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13133_ net149 net111 _06707_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__mux2_1
X_10345_ _04649_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13064_ net1146 _04883_ _06635_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__mux2_1
X_10276_ net1052 _03255_ _04611_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12015_ _05794_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13966_ _01600_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_401 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15705_ clknet_leaf_17_clk _01280_ VGND VGND VPWR VPWR cpuregs\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_557 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12917_ _06593_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__clkbuf_1
X_13897_ _01563_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_760 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_445 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15636_ clknet_leaf_122_clk _01211_ VGND VGND VPWR VPWR cpuregs\[23\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12848_ net556 _06554_ _06557_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_158_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15567_ clknet_leaf_15_clk _01142_ VGND VGND VPWR VPWR cpuregs\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12779_ _03020_ _01861_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__or2_1
X_14518_ clknet_leaf_13_clk _00176_ VGND VGND VPWR VPWR cpuregs\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_16_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15498_ clknet_leaf_92_clk _01083_ VGND VGND VPWR VPWR mem_rdata_q\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_865 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14449_ clknet_leaf_36_clk _00107_ VGND VGND VPWR VPWR cpuregs\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold904 cpuregs\[2\]\[22\] VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 cpuregs\[7\]\[9\] VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 cpuregs\[18\]\[19\] VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold937 cpuregs\[18\]\[2\] VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold948 cpuregs\[3\]\[18\] VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ _03425_ _04431_ _04433_ _04435_ _00016_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__a221o_1
Xhold959 cpuregs\[20\]\[9\] VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08941_ cpuregs\[8\]\[0\] cpuregs\[9\]\[0\] cpuregs\[10\]\[0\] cpuregs\[11\]\[0\]
+ _03406_ _03410_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__mux4_1
X_08872_ _03351_ _03352_ _03261_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_4_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07823_ _02438_ _02439_ _02442_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07754_ reg_pc\[30\] decoded_imm\[30\] VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_140_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07685_ _02310_ _02311_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_91_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_2
X_09424_ _02112_ _03660_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09355_ _03814_ _03816_ _03818_ _03820_ _03429_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08306_ _02608_ _02894_ _02895_ _02897_ VGND VGND VPWR VPWR alu_out\[28\] sky130_fd_sc_hd__a31o_1
XFILLER_0_118_854 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09286_ cpuregs\[16\]\[7\] cpuregs\[17\]\[7\] cpuregs\[18\]\[7\] cpuregs\[19\]\[7\]
+ _03601_ _03583_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08237_ _02396_ _02826_ _02834_ _02585_ VGND VGND VPWR VPWR alu_out\[22\] sky130_fd_sc_hd__a22o_2
XFILLER_0_90_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08168_ _02213_ _02770_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08099_ _02682_ _02694_ _02695_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10130_ _04534_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ _04496_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13820_ net1204 _06981_ _07086_ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__mux2_1
X_13751_ _07057_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_10963_ _04992_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_82_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12702_ cpuregs\[8\]\[29\] cpuregs\[9\]\[29\] cpuregs\[10\]\[29\] cpuregs\[11\]\[29\]
+ _05970_ _03137_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_905 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13682_ cpuregs\[23\]\[26\] _06979_ _07014_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__mux2_1
X_10894_ net936 _04881_ _04922_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__mux2_1
X_15421_ clknet_leaf_151_clk _01011_ VGND VGND VPWR VPWR cpuregs\[18\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12633_ _03142_ _06372_ _06376_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__or3_1
XFILLER_0_156_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_66_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15352_ clknet_leaf_68_clk _00942_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dfxtp_1
X_12564_ cpuregs\[0\]\[23\] cpuregs\[1\]\[23\] cpuregs\[2\]\[23\] cpuregs\[3\]\[23\]
+ _06055_ _05829_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14303_ _03180_ _04524_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11515_ net361 _05217_ _05387_ _05264_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__a31o_1
X_15283_ clknet_leaf_92_clk _00876_ VGND VGND VPWR VPWR decoded_imm_j\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12495_ cpuregs\[4\]\[20\] cpuregs\[5\]\[20\] cpuregs\[6\]\[20\] cpuregs\[7\]\[20\]
+ _06011_ _06156_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14234_ _01742_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__clkbuf_1
X_11446_ _05288_ _05338_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_879 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14165_ cpuregs\[7\]\[29\] _06985_ _01696_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__mux2_1
X_11377_ _05272_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_150_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13116_ net140 net102 _06696_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__mux2_1
X_10328_ _04640_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__clkbuf_1
X_14096_ _01669_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__clkbuf_1
X_13047_ _06661_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__clkbuf_1
X_10259_ net1275 _03202_ _04600_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_800 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14998_ clknet_leaf_107_clk _00656_ VGND VGND VPWR VPWR reg_next_pc\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13949_ net1158 _06973_ _01588_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_765 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07470_ net172 VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_85_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15619_ clknet_leaf_44_clk _01194_ VGND VGND VPWR VPWR cpuregs\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_09140_ _03610_ _03611_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_733 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09071_ _01844_ _01992_ _03391_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08022_ _02613_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_554 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold701 cpuregs\[5\]\[31\] VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 cpuregs\[11\]\[27\] VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold723 cpuregs\[1\]\[30\] VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold734 cpuregs\[21\]\[10\] VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_877 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold745 cpuregs\[28\]\[27\] VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold756 cpuregs\[8\]\[7\] VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 cpuregs\[29\]\[10\] VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 cpuregs\[15\]\[27\] VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _03500_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__or2_1
Xhold789 cpuregs\[27\]\[10\] VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08924_ _01847_ decoded_imm\[0\] VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__or2_1
X_08855_ reg_pc\[24\] reg_pc\[23\] _03326_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07806_ net189 net221 VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__or2_1
X_08786_ reg_pc\[15\] _03272_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _02018_ _02349_ _02360_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_803 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_67_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_64_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07668_ count_cycle\[24\] _02051_ _02294_ _02295_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09407_ _03869_ _03870_ _03402_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_426 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07599_ reg_pc\[19\] decoded_imm\[19\] VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_48_796 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09338_ _03802_ _03803_ _03552_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_893 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_117_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09269_ _03704_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11300_ _05186_ _05217_ _05218_ _01885_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_153_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12280_ cpuregs\[8\]\[11\] cpuregs\[9\]\[11\] cpuregs\[10\]\[11\] cpuregs\[11\]\[11\]
+ _03150_ _05917_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_120_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11231_ net526 _05165_ _05169_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_56_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_173 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11162_ _05121_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_1
X_10113_ _04522_ _04524_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__nor2_4
X_11093_ net1113 _05072_ _05044_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__o21ai_1
X_15970_ clknet_leaf_75_clk _01542_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_1
X_14921_ clknet_leaf_117_clk _00579_ VGND VGND VPWR VPWR count_instr\[30\] sky130_fd_sc_hd__dfxtp_1
X_10044_ net1287 _03179_ _04487_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__mux2_1
Xhold50 mem_rdata[17] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 net33 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 count_cycle\[0\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkdlybuf4s25_1
X_14852_ clknet_leaf_150_clk _00510_ VGND VGND VPWR VPWR cpuregs\[20\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold83 count_instr\[37\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 instr_andi VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ cpuregs\[3\]\[19\] _06964_ _07075_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__mux2_1
X_14783_ clknet_leaf_124_clk _00441_ VGND VGND VPWR VPWR cpuregs\[16\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11995_ net42 net73 _05774_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_55_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_2
X_13734_ _07048_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__clkbuf_1
X_10946_ net820 _04865_ _04981_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_86_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_156_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13665_ net1391 _06962_ _07003_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__mux2_1
X_10877_ _04947_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_100_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_262 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12616_ _05912_ _06360_ _06193_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__o21a_1
X_15404_ clknet_leaf_91_clk _00994_ VGND VGND VPWR VPWR decoded_imm\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13596_ _03328_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__buf_2
XFILLER_0_26_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_318 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15335_ clknet_leaf_70_clk _00925_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dfxtp_1
X_12547_ cpuregs\[24\]\[22\] cpuregs\[25\]\[22\] cpuregs\[26\]\[22\] cpuregs\[27\]\[22\]
+ _05970_ _03108_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15266_ clknet_leaf_85_clk _00859_ VGND VGND VPWR VPWR decoded_imm_j\[9\] sky130_fd_sc_hd__dfxtp_1
X_12478_ cpuregs\[12\]\[19\] cpuregs\[13\]\[19\] cpuregs\[14\]\[19\] cpuregs\[15\]\[19\]
+ _05913_ _05994_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
*XANTENNA_3 _01674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14217_ net1354 _06969_ _01732_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11429_ _05321_ _05322_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_105_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15197_ clknet_leaf_70_clk alu_out\[10\] VGND VGND VPWR VPWR alu_out_q\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_10_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14148_ _01697_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14079_ net1032 _06966_ _01660_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08640_ _03080_ _03141_ _03157_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_87_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer15 _05127_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_1
Xrebuffer26 _05168_ VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_1
Xrebuffer37 net397 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_1
X_08571_ _03061_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_46_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07522_ reg_pc\[14\] decoded_imm\[14\] VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_157_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07453_ _02094_ _02095_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07384_ net5 net22 _01844_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09123_ _03459_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_287 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09054_ _03527_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_641 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08005_ _02608_ _02616_ _02617_ _02620_ _02498_ VGND VGND VPWR VPWR alu_out\[4\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold520 cpuregs\[28\]\[5\] VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 cpuregs\[16\]\[31\] VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 cpuregs\[1\]\[10\] VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold553 cpuregs\[10\]\[12\] VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_860 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold564 cpuregs\[8\]\[0\] VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 cpuregs\[21\]\[24\] VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 cpuregs\[29\]\[0\] VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 instr_lw VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__dlygate4sd3_1
X_09956_ _04399_ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_51_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ reg_out\[31\] alu_out_q\[31\] _03176_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__mux2_1
X_09887_ _04266_ _04335_ _03075_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__o21ai_1
X_08838_ _03323_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08769_ net1215 _03263_ _03249_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_2
X_10800_ _04906_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__clkbuf_1
X_11780_ count_cycle\[16\] _05628_ count_cycle\[17\] VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10731_ _03328_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13450_ net846 _04877_ _06874_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_82_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10662_ _04524_ _04744_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__nor2_4
XFILLER_0_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12401_ _06155_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__clkbuf_1
X_13381_ _06846_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10593_ _03183_ _04481_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__nor2_2
XFILLER_0_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15120_ clknet_leaf_74_clk _00746_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_1
X_12332_ _05845_ _06086_ _06088_ _03139_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15051_ clknet_leaf_115_clk _00709_ VGND VGND VPWR VPWR count_cycle\[34\] sky130_fd_sc_hd__dfxtp_1
X_12263_ _03061_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14002_ net944 _06958_ _01613_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__mux2_1
X_11214_ count_instr\[51\] _05156_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__and2_1
X_12194_ _02489_ _05956_ _05863_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__mux2_1
Xoutput40 net40 VGND VGND VPWR VPWR mem_addr[15] sky130_fd_sc_hd__clkbuf_4
Xoutput51 net51 VGND VGND VPWR VPWR mem_addr[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput62 net62 VGND VGND VPWR VPWR mem_addr[7] sky130_fd_sc_hd__clkbuf_4
Xoutput73 net73 VGND VGND VPWR VPWR mem_la_addr[17] sky130_fd_sc_hd__clkbuf_4
X_11145_ net578 _05107_ _05090_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__o21ai_1
Xoutput84 net84 VGND VGND VPWR VPWR mem_la_addr[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput95 net95 VGND VGND VPWR VPWR mem_la_addr[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11076_ count_instr\[7\] count_instr\[6\] _05051_ _05061_ VGND VGND VPWR VPWR _05062_
+ sky130_fd_sc_hd__and4_1
X_15953_ clknet_leaf_12_clk _01525_ VGND VGND VPWR VPWR cpuregs\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_14904_ clknet_leaf_102_clk net468 VGND VGND VPWR VPWR count_instr\[13\] sky130_fd_sc_hd__dfxtp_1
X_10027_ cpuregs\[8\]\[30\] cpuregs\[9\]\[30\] cpuregs\[10\]\[30\] cpuregs\[11\]\[30\]
+ _03680_ _03443_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_69_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ clknet_leaf_11_clk _01456_ VGND VGND VPWR VPWR cpuregs\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ clknet_leaf_29_clk _00493_ VGND VGND VPWR VPWR cpuregs\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_814 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_28_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_19_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14766_ clknet_leaf_42_clk _00424_ VGND VGND VPWR VPWR cpuregs\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11978_ _05775_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_82_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13717_ net1126 _06945_ _07039_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__mux2_1
X_10929_ cpuregs\[20\]\[14\] _04848_ _04970_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14697_ clknet_leaf_18_clk _00355_ VGND VGND VPWR VPWR cpuregs\[27\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_711 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_73_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13648_ _06991_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__buf_4
XFILLER_0_27_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_755 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13579_ _06959_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_30_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15318_ clknet_leaf_141_clk _00908_ VGND VGND VPWR VPWR cpuregs\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15249_ clknet_leaf_76_clk _00842_ VGND VGND VPWR VPWR instr_sltu sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09810_ _03574_ _04252_ _04261_ _03527_ reg_pc\[23\] VGND VGND VPWR VPWR _04262_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09741_ _03435_ _04194_ _03425_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09672_ _03446_ _04127_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__or2_1
X_08623_ _03123_ _03127_ _03131_ _03136_ _03140_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_19_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08554_ _03073_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_38_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07505_ _01977_ _02139_ _02141_ _01928_ _02144_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__a221o_1
X_08485_ _03016_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_1
XFILLER_0_147_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07436_ _01893_ _02079_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07367_ count_instr\[4\] _01965_ count_cycle\[36\] _02014_ VGND VGND VPWR VPWR _02015_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09106_ cpuregs\[0\]\[3\] cpuregs\[1\]\[3\] cpuregs\[2\]\[3\] cpuregs\[3\]\[3\] _03439_
+ _03576_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_150_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07298_ instr_rdinstrh instr_rdcycleh instr_rdinstr VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__nor3_2
XFILLER_0_21_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_566 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09037_ cpuregs\[6\]\[1\] cpuregs\[7\]\[1\] _03406_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_68_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold350 reg_pc\[22\] VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 reg_pc\[14\] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold372 cpuregs\[11\]\[7\] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 cpuregs\[23\]\[23\] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold394 cpuregs\[22\]\[24\] VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__dlygate4sd3_1
X_09939_ _04384_ _04385_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_148_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_12950_ mem_rdata_q\[8\] net31 _06589_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__mux2_1
Xhold1050 _01915_ VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ count_cycle\[55\] _05714_ _01905_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12881_ _05041_ _06547_ _06568_ _06529_ net481 VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__a32o_1
*XANTENNA_201 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_212 _03401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
*XANTENNA_223 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11832_ _05036_ net365 VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__nor2_1
X_14620_ clknet_leaf_155_clk _00278_ VGND VGND VPWR VPWR cpuregs\[21\]\[18\] sky130_fd_sc_hd__dfxtp_1
*XANTENNA_234 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ clknet_leaf_14_clk _00209_ VGND VGND VPWR VPWR cpuregs\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11763_ net531 count_cycle\[11\] count_cycle\[12\] _05613_ VGND VGND VPWR VPWR _05620_
+ sky130_fd_sc_hd__and4_4
XTAP_TAPCELL_ROW_64_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10714_ _04853_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__clkbuf_1
X_13502_ net1009 _04860_ _06910_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14482_ clknet_leaf_55_clk _00140_ VGND VGND VPWR VPWR cpuregs\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11694_ _05253_ _05566_ _05032_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13433_ _06851_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__buf_4
X_10645_ net927 _03341_ _04804_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_91_680 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13364_ _06837_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer6 _05667_ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
X_10576_ _04772_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12315_ _03045_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__clkbuf_4
X_15103_ clknet_leaf_102_clk _07127_ VGND VGND VPWR VPWR reg_out\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16083_ net125 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_2
X_13295_ net1285 _04858_ _06791_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15034_ clknet_leaf_122_clk _00692_ VGND VGND VPWR VPWR count_cycle\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_791 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12246_ _03149_ _06006_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12177_ _05938_ _05939_ _03124_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__mux2_1
X_11128_ count_instr\[25\] count_instr\[24\] VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11059_ net462 VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__inv_2
X_15936_ clknet_leaf_58_clk _01508_ VGND VGND VPWR VPWR cpuregs\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15867_ clknet_leaf_132_clk _01439_ VGND VGND VPWR VPWR cpuregs\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_14818_ clknet_leaf_127_clk _00476_ VGND VGND VPWR VPWR cpuregs\[25\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15798_ clknet_leaf_140_clk _01373_ VGND VGND VPWR VPWR cpuregs\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14749_ clknet_leaf_156_clk _00407_ VGND VGND VPWR VPWR cpuregs\[26\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_08270_ _02849_ _02855_ _02853_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07221_ instr_sltu instr_sltiu net455 VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_226 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_719 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07152_ net414 VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_112_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07985_ net251 _02601_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__xnor2_1
X_09724_ decoded_imm\[21\] net184 VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__nor2_1
X_09655_ reg_pc\[18\] _03528_ _04111_ _03626_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_143_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08606_ _03037_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_2_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09586_ cpuregs\[4\]\[16\] cpuregs\[5\]\[16\] cpuregs\[6\]\[16\] cpuregs\[7\]\[16\]
+ _03440_ _03451_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__mux4_1
X_08537_ decoded_imm_j\[11\] decoded_imm_j\[4\] VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_46_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_38_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08468_ reg_next_pc\[26\] reg_out\[26\] _02991_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_362 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_80_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07419_ _02061_ _02063_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08399_ reg_next_pc\[5\] reg_out\[5\] _02949_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10430_ _04694_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_900 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_116_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10361_ _04657_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12100_ decoded_imm\[3\] _01906_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13080_ mem_state\[0\] _06676_ _06680_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__mux2_1
X_10292_ cpuregs\[2\]\[19\] _03307_ _04611_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_103_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12031_ _05803_ _05036_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__nor2_2
Xhold180 reg_next_pc\[30\] VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 count_cycle\[19\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13982_ _01609_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__clkbuf_1
X_15721_ clknet_leaf_0_clk _01296_ VGND VGND VPWR VPWR cpuregs\[22\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_12933_ _06601_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15652_ clknet_leaf_43_clk _01227_ VGND VGND VPWR VPWR cpuregs\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12864_ mem_rdata_q\[28\] mem_rdata_q\[27\] mem_rdata_q\[26\] mem_rdata_q\[25\] VGND
+ VGND VPWR VPWR _06563_ sky130_fd_sc_hd__or4_2
XFILLER_0_96_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14603_ clknet_leaf_53_clk _00261_ VGND VGND VPWR VPWR cpuregs\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11815_ _05655_ _05656_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12795_ mem_rdata_q\[5\] net28 _01857_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15583_ clknet_leaf_45_clk _01158_ VGND VGND VPWR VPWR cpuregs\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11746_ _05607_ _05608_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__nor2_1
X_14534_ clknet_leaf_97_clk _00192_ VGND VGND VPWR VPWR cpuregs\[13\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_800 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14465_ clknet_leaf_136_clk _00123_ VGND VGND VPWR VPWR cpuregs\[12\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_11677_ _05549_ _05550_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_546 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13416_ _06865_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__clkbuf_1
X_10628_ cpuregs\[15\]\[16\] _03287_ _04793_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14396_ clknet_leaf_141_clk _00059_ VGND VGND VPWR VPWR cpuregs\[11\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13347_ cpuregs\[19\]\[11\] _04842_ _06827_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__mux2_1
Xpicorv32_305 VGND VGND VPWR VPWR picorv32_305/HI pcpi_insn[15] sky130_fd_sc_hd__conb_1
XFILLER_0_3_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xpicorv32_316 VGND VGND VPWR VPWR picorv32_316/HI pcpi_insn[26] sky130_fd_sc_hd__conb_1
X_10559_ _04763_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__clkbuf_1
Xpicorv32_327 VGND VGND VPWR VPWR picorv32_327/HI trace_data[4] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_338 VGND VGND VPWR VPWR picorv32_338/HI trace_data[15] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_94_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_349 VGND VGND VPWR VPWR picorv32_349/HI trace_data[26] sky130_fd_sc_hd__conb_1
X_13278_ _06792_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15017_ clknet_leaf_111_clk _00675_ VGND VGND VPWR VPWR count_cycle\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_110_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12229_ _05990_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_783 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_75_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07770_ _02389_ _02390_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_160_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15919_ clknet_leaf_18_clk _01491_ VGND VGND VPWR VPWR cpuregs\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_160_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09440_ _03651_ _03901_ _03902_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_125_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09371_ _03767_ _03830_ _03834_ _03795_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_91_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08322_ _02910_ _02911_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_682 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_129_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08253_ _02756_ net237 net236 _02848_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_145_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07204_ cpu_state\[6\] cpu_state\[5\] VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_41_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_61_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08184_ _02784_ _02785_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_549 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_160_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_15_577 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_113_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput230 net230 VGND VGND VPWR VPWR pcpi_rs2[5] sky130_fd_sc_hd__buf_2
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07968_ net97 net108 instr_sub VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__o21ba_1
X_09707_ _03746_ _04161_ _03419_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__o21a_1
X_07899_ _02496_ _02497_ net250 VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__a21bo_1
X_09638_ cpuregs\[20\]\[18\] cpuregs\[21\]\[18\] cpuregs\[22\]\[18\] cpuregs\[23\]\[18\]
+ _03594_ _03442_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_569 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09569_ _02177_ net243 VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11600_ _05185_ _05479_ _05480_ _05257_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _06132_ _06317_ _06326_ _06153_ decoded_imm\[23\] VGND VGND VPWR VPWR _06327_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_108_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11531_ _05186_ _05416_ _05417_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14250_ _01750_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__clkbuf_1
X_11462_ _05352_ _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_156_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13201_ net484 _06742_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__and2_1
X_10413_ net1015 _03255_ _04684_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__mux2_1
X_14181_ cpuregs\[8\]\[4\] _06933_ _01710_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11393_ decoded_imm_j\[4\] _05197_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_763 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13132_ _06709_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__clkbuf_1
X_10344_ net1341 _03255_ _04647_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13063_ _06669_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__clkbuf_1
X_10275_ _04612_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__clkbuf_1
X_12014_ net51 net82 _05785_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13965_ net1247 _06989_ _01565_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__mux2_1
X_15704_ clknet_leaf_130_clk _01279_ VGND VGND VPWR VPWR cpuregs\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12916_ decoded_imm_j\[6\] _01088_ _03169_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13896_ net676 _06989_ _07099_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15635_ clknet_leaf_147_clk _01210_ VGND VGND VPWR VPWR cpuregs\[23\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12847_ is_lb_lh_lw_lbu_lhu _06531_ _06543_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__and3_1
XFILLER_0_158_457 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_29_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15566_ clknet_leaf_11_clk _01141_ VGND VGND VPWR VPWR cpuregs\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12778_ latched_is_lb _06509_ _06511_ _05257_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_120_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14517_ clknet_leaf_31_clk _00175_ VGND VGND VPWR VPWR cpuregs\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11729_ net431 net435 _05141_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_71_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15497_ clknet_leaf_93_clk _01082_ VGND VGND VPWR VPWR mem_rdata_q\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14448_ clknet_leaf_33_clk _00106_ VGND VGND VPWR VPWR cpuregs\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_825 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_4_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_25_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_769 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold905 cpuregs\[23\]\[0\] VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ clknet_leaf_38_clk _00042_ VGND VGND VPWR VPWR cpuregs\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold916 cpuregs\[2\]\[3\] VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 cpuregs\[24\]\[21\] VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold938 cpuregs\[16\]\[6\] VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold949 cpuregs\[9\]\[18\] VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_23_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08940_ _03414_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_788 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08871_ reg_pc\[26\] reg_pc\[25\] _03338_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_127_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07822_ _02440_ _02441_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07753_ reg_pc\[30\] decoded_imm\[30\] VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_140_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07684_ reg_pc\[25\] decoded_imm\[25\] VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_140_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09423_ _03488_ _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09354_ _03435_ _03819_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08305_ _02595_ _02896_ _02438_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__o21ba_1
X_09285_ _03454_ _03752_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_797 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_118_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08236_ _02831_ _02833_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_814 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08167_ net211 _02769_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08098_ _02704_ _02705_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10060_ net818 _03235_ _04487_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13750_ cpuregs\[29\]\[26\] _06979_ _07050_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__mux2_1
X_10962_ cpuregs\[20\]\[30\] _04881_ _04958_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__mux2_1
X_12701_ _03143_ _06441_ _06182_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__o21a_1
X_13681_ _07020_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__clkbuf_1
X_10893_ _04955_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15420_ clknet_leaf_158_clk _01010_ VGND VGND VPWR VPWR cpuregs\[18\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12632_ _05845_ _06373_ _06375_ _03139_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15351_ clknet_leaf_68_clk _00941_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12563_ cpuregs\[4\]\[23\] cpuregs\[5\]\[23\] cpuregs\[6\]\[23\] cpuregs\[7\]\[23\]
+ _06011_ _06156_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14302_ _01776_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__clkbuf_1
X_11514_ _05289_ _05400_ _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__nand3_1
XFILLER_0_25_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_600 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_53_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15282_ clknet_leaf_93_clk _00875_ VGND VGND VPWR VPWR decoded_imm_j\[11\] sky130_fd_sc_hd__dfxtp_2
X_12494_ _06244_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14233_ net804 _06985_ _01732_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__mux2_1
X_11445_ _05204_ _05206_ _05312_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_151_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14164_ _01705_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_74_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_165 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11376_ _05263_ net1329 _05268_ _05274_ _05257_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__o221a_1
X_13115_ _06700_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10327_ net1280 _03202_ _04636_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__mux2_1
X_14095_ net870 _06983_ _01660_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__mux2_1
X_13046_ net885 _04865_ _06658_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__mux2_1
X_10258_ _04603_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__clkbuf_1
X_10189_ net1064 _03194_ _04564_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_812 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14997_ clknet_leaf_86_clk _00655_ VGND VGND VPWR VPWR reg_next_pc\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13948_ _01591_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13879_ _01554_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_265 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15618_ clknet_leaf_39_clk _01193_ VGND VGND VPWR VPWR cpuregs\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15549_ clknet_leaf_81_clk _00022_ VGND VGND VPWR VPWR cpu_state\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09070_ _03540_ _03541_ _03539_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_184 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08021_ _02633_ _02634_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_566 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold702 cpuregs\[30\]\[29\] VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 cpuregs\[1\]\[16\] VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_688 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold724 cpuregs\[20\]\[2\] VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 cpuregs\[22\]\[27\] VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 cpuregs\[17\]\[14\] VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold757 cpuregs\[7\]\[17\] VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 cpuregs\[23\]\[9\] VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ cpuregs\[24\]\[28\] cpuregs\[25\]\[28\] cpuregs\[26\]\[28\] cpuregs\[27\]\[28\]
+ _03636_ _03637_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold779 reg_next_pc\[3\] VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08923_ net171 decoded_imm\[0\] VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08854_ reg_pc\[23\] _03326_ reg_pc\[24\] VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__a21oi_1
X_07805_ _02395_ _02404_ _02408_ _02423_ _02424_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__o221a_1
X_08785_ reg_out\[15\] alu_out_q\[15\] _03175_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ _02058_ _02357_ _02359_ _01968_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07667_ count_instr\[56\] _02052_ _02055_ count_cycle\[56\] VGND VGND VPWR VPWR _02295_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09406_ cpuregs\[0\]\[11\] cpuregs\[1\]\[11\] cpuregs\[2\]\[11\] cpuregs\[3\]\[11\]
+ _03405_ _03496_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_137_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07598_ count_cycle\[19\] _02051_ _02229_ _02230_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_63_712 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09337_ cpuregs\[0\]\[9\] cpuregs\[1\]\[9\] cpuregs\[2\]\[9\] cpuregs\[3\]\[9\] _03800_
+ _03407_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_909 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_118_652 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09268_ _03734_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__or2b_1
XFILLER_0_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_406 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08219_ _02816_ _02817_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_153_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09199_ _02008_ _03660_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__and2_1
X_11230_ _05040_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_56_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_176 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11161_ _05119_ _05113_ _05120_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__and3b_1
XFILLER_0_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10112_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__clkbuf_8
X_11092_ count_instr\[14\] _05072_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__and2_1
X_14920_ clknet_leaf_117_clk _00578_ VGND VGND VPWR VPWR count_instr\[29\] sky130_fd_sc_hd__dfxtp_1
X_10043_ _04486_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__clkbuf_8
Xhold51 mem_rdata[20] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 mem_rdata[16] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ clknet_leaf_122_clk _00509_ VGND VGND VPWR VPWR cpuregs\[20\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold73 mem_wordsize\[0\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold84 mem_rdata_q\[27\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 count_cycle\[54\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _07084_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14782_ clknet_leaf_148_clk _00440_ VGND VGND VPWR VPWR cpuregs\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11994_ _05783_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__clkbuf_1
X_13733_ cpuregs\[29\]\[18\] _06962_ _07039_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__mux2_1
X_10945_ _04983_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_917 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13664_ _07011_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__clkbuf_1
X_10876_ net958 _04863_ _04945_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15403_ clknet_leaf_82_clk _00993_ VGND VGND VPWR VPWR decoded_imm\[5\] sky130_fd_sc_hd__dfxtp_2
X_12615_ cpuregs\[28\]\[25\] cpuregs\[29\]\[25\] cpuregs\[30\]\[25\] cpuregs\[31\]\[25\]
+ _06191_ _05914_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13595_ _06970_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15334_ clknet_leaf_70_clk _00924_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dfxtp_2
X_12546_ _03142_ _06289_ _06293_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_266 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_81_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15265_ clknet_leaf_90_clk _00858_ VGND VGND VPWR VPWR decoded_imm_j\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12477_ _06226_ _06227_ _06014_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
*XANTENNA_4 _01823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14216_ _01733_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__clkbuf_1
X_11428_ decoded_imm_j\[7\] _05204_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15196_ clknet_leaf_70_clk alu_out\[9\] VGND VGND VPWR VPWR alu_out_q\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_837 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_14147_ net1000 _06966_ _01696_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__mux2_1
X_11359_ _05258_ reg_pc\[30\] _05239_ _05260_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__o211a_1
X_14078_ _01637_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__buf_4
X_13029_ net1006 _04848_ _06647_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__mux2_1
Xrebuffer16 _05116_ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_1
Xrebuffer27 _05116_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_1
X_08570_ _03083_ _03088_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__nor2_1
Xrebuffer38 net398 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07521_ reg_pc\[14\] decoded_imm\[14\] VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_157_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07452_ reg_pc\[9\] decoded_imm\[9\] VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_937 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_07383_ net198 VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09122_ _03456_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__buf_8
XFILLER_0_161_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_33_918 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_09053_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_135_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_430 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_143_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_352 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_603 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_08004_ _02595_ _02619_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_142_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold510 cpuregs\[25\]\[5\] VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold521 cpuregs\[11\]\[8\] VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 cpuregs\[20\]\[1\] VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap240 _02570_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__buf_1
Xhold543 cpuregs\[7\]\[11\] VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 cpuregs\[26\]\[26\] VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
Xhold565 cpuregs\[10\]\[16\] VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 cpuregs\[8\]\[9\] VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold587 cpuregs\[24\]\[5\] VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 cpuregs\[5\]\[23\] VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09955_ _04400_ _04401_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_51_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08906_ _03382_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__clkbuf_1
X_09886_ _02316_ _03617_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__nor2_1
X_08837_ net1352 _03322_ _03315_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__mux2_1
X_08768_ _03262_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__clkbuf_4
X_07719_ count_instr\[27\] _01949_ count_cycle\[59\] _01947_ VGND VGND VPWR VPWR _02344_
+ sky130_fd_sc_hd__a22o_1
X_08699_ net1183 _03202_ _03185_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10730_ _04864_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10661_ _03178_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_706 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_12400_ net209 _06154_ _06052_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__mux2_1
X_13380_ net877 _04875_ _06838_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10592_ _04780_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12331_ _03042_ _06087_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_132 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_35_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15050_ clknet_leaf_115_clk _00708_ VGND VGND VPWR VPWR count_cycle\[33\] sky130_fd_sc_hd__dfxtp_1
X_12262_ _03143_ _06021_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__or2_1
X_11213_ _05156_ _05157_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__nor2_1
X_14001_ _01619_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12193_ _05901_ _05945_ _05955_ _05904_ decoded_imm\[7\] VGND VGND VPWR VPWR _05956_
+ sky130_fd_sc_hd__a32o_1
Xoutput41 net41 VGND VGND VPWR VPWR mem_addr[16] sky130_fd_sc_hd__clkbuf_4
Xoutput52 net52 VGND VGND VPWR VPWR mem_addr[27] sky130_fd_sc_hd__clkbuf_4
X_11144_ count_instr\[30\] count_instr\[29\] count_instr\[28\] _05103_ VGND VGND VPWR
+ VPWR _05109_ sky130_fd_sc_hd__and4_1
Xoutput63 net63 VGND VGND VPWR VPWR mem_addr[8] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 VGND VGND VPWR VPWR mem_la_addr[18] sky130_fd_sc_hd__buf_2
Xoutput85 net85 VGND VGND VPWR VPWR mem_la_addr[29] sky130_fd_sc_hd__buf_2
Xoutput96 net96 VGND VGND VPWR VPWR mem_la_read sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_11075_ count_instr\[9\] count_instr\[8\] VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__and2_1
X_15952_ clknet_leaf_16_clk _01524_ VGND VGND VPWR VPWR cpuregs\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_14903_ clknet_leaf_102_clk _00561_ VGND VGND VPWR VPWR count_instr\[12\] sky130_fd_sc_hd__dfxtp_1
X_10026_ _03448_ _04470_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__or2_1
X_15883_ clknet_leaf_30_clk _01455_ VGND VGND VPWR VPWR cpuregs\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ clknet_leaf_58_clk _00492_ VGND VGND VPWR VPWR cpuregs\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14765_ clknet_leaf_26_clk _00423_ VGND VGND VPWR VPWR cpuregs\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11977_ net63 net94 _05774_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13716_ _07027_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_82_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10928_ _04974_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14696_ clknet_leaf_24_clk _00354_ VGND VGND VPWR VPWR cpuregs\[27\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13647_ _07002_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__clkbuf_1
X_10859_ cpuregs\[25\]\[13\] _04846_ _04934_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_767 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_13578_ net798 _06958_ _06946_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15317_ clknet_leaf_133_clk _00907_ VGND VGND VPWR VPWR cpuregs\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12529_ cpuregs\[24\]\[21\] cpuregs\[25\]\[21\] cpuregs\[26\]\[21\] cpuregs\[27\]\[21\]
+ _06074_ _03151_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_597 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_15248_ clknet_leaf_76_clk _00841_ VGND VGND VPWR VPWR instr_slt sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15179_ clknet_leaf_61_clk _00804_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_130_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09740_ cpuregs\[16\]\[21\] cpuregs\[17\]\[21\] cpuregs\[18\]\[21\] cpuregs\[19\]\[21\]
+ _03548_ _03549_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__mux4_1
.ends picorv32_m

