* Spice description of nts_x1
* Spice driver version 1586745115
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:16

* INTERF cmd i nq vdd vss 


.subckt nts_x1 5 6 4 1 8 
* NET 1 = vdd
* NET 4 = nq
* NET 5 = cmd
* NET 6 = i
* NET 8 = vss
Mtr_00006 4 3 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 1 5 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00004 2 6 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00003 4 5 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 8 5 3 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 7 6 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C8 1 8 2.22211e-15
C6 3 8 1.32368e-15
C5 4 8 2.15173e-15
C4 5 8 2.68055e-15
C3 6 8 2.34207e-15
C1 8 8 1.86659e-15
.ends nts_x1

