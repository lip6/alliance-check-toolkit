* MacroLib

* NPN_05v5_W1u00L1u00
.subckt NPN_05v5_W1u00L1u00 collector base emitter
Xnpn collector base emitter sky130_fd_pr__npn_05v5_W1p00L1p00
.ends NPN_05v5_W1u00L1u00

* NPN_05v5_W1u00L2u00
.subckt NPN_05v5_W1u00L2u00 collector base emitter
Xnpn collector base emitter sky130_fd_pr__npn_05v5_W1p00L2p00
.ends NPN_05v5_W1u00L2u00

* PNP_05v5_W0u68L0u68
.subckt PNP_05v5_W0u68L0u68 collector base emitter
Xpnp collector base emitter sky130_fd_pr__pnp_05v5_W0p68L0p68
.ends PNP_05v5_W0u68L0u68

* PNP_05v5_W3u40L3u40
.subckt PNP_05v5_W3u40L3u40 collector base emitter
Xpnp collector base emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
.ends PNP_05v5_W3u40L3u40
