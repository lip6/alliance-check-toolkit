* Spice description of mx2_x4
* Spice driver version -990253285
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:45

* INTERF cmd i0 i1 q vdd vss 


.subckt mx2_x4 10 5 6 4 3 11 
* NET 3 = vdd
* NET 4 = q
* NET 5 = i0
* NET 6 = i1
* NET 10 = cmd
* NET 11 = vss
Mtr_00014 4 9 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 3 6 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00012 2 5 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00011 3 10 12 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00010 1 12 9 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00009 9 10 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00008 3 9 4 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 4 9 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00006 11 6 8 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00005 9 12 7 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00004 7 5 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00003 11 10 12 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00002 11 9 4 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 8 10 9 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
C10 3 11 4.11856e-15
C9 4 11 2.15173e-15
C8 5 11 1.77589e-15
C7 6 11 2.47522e-15
C4 9 11 2.17098e-15
C3 10 11 2.98806e-15
C2 11 11 3.15255e-15
C1 12 11 2.72381e-15
.ends mx2_x4

