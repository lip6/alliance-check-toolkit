* Spice description of a3_x4
* Spice driver version 533778203
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:30

* INTERF i0 i1 i2 q vdd vss 


.subckt a3_x4 6 7 2 4 1 5 
* NET 1 = vdd
* NET 2 = i2
* NET 4 = q
* NET 5 = vss
* NET 6 = i0
* NET 7 = i1
Mtr_00010 1 9 4 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 4 9 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 1 2 9 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 9 7 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 1 6 9 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00005 5 9 4 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 4 9 5 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 5 2 3 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 3 7 8 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 8 6 9 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C9 1 5 2.94067e-15
C8 2 5 1.49465e-15
C6 4 5 2.15173e-15
C5 5 5 2.35713e-15
C4 6 5 1.45814e-15
C3 7 5 1.45814e-15
C1 9 5 2.88673e-15
.ends a3_x4

