-- no model for and2_x1
