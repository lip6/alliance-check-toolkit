* npn_s
.param
+ dkisnpn1x1=5.9826e-01 dkbfnpn1x1=4.7271e-01
+ dkisnpn1x2=6.2301e-01 dkbfnpn1x2=4.6386e-01
+ dkisnpnpolyhv=0.591 dkbfnpnpolyhv=0.479
