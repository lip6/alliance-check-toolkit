* Coriolis Structural SPICE Driver
* Generated on Sep 25, 2024, 13:06
* Cell/Subckt "arlet6502_cts_r".
* 
* INTERF vss
* INTERF vdd
* INTERF reset
* INTERF clk
* INTERF WE
* INTERF RDY
* INTERF NMI
* INTERF IRQ
* INTERF DO[7]
* INTERF DO[6]
* INTERF DO[5]
* INTERF DO[4]
* INTERF DO[3]
* INTERF DO[2]
* INTERF DO[1]
* INTERF DO[0]
* INTERF DI[7]
* INTERF DI[6]
* INTERF DI[5]
* INTERF DI[4]
* INTERF DI[3]
* INTERF DI[2]
* INTERF DI[1]
* INTERF DI[0]
* INTERF A[9]
* INTERF A[8]
* INTERF A[7]
* INTERF A[6]
* INTERF A[5]
* INTERF A[4]
* INTERF A[3]
* INTERF A[2]
* INTERF A[15]
* INTERF A[14]
* INTERF A[13]
* INTERF A[12]
* INTERF A[11]
* INTERF A[10]
* INTERF A[1]
* INTERF A[0]

* Terminal models (aka standard cells) used througout all the hierarchy.
.include decap_w0.spi
.include tie.spi
.include nand2_x0.spi
.include mux2_x1.spi
.include and2_x1.spi
.include buf_x4.spi
.include and4_x1.spi
.include and21nor_x0.spi
.include or2_x1.spi
.include or21nand_x0.spi
.include nand3_x0.spi
.include nand4_x0.spi
.include and3_x1.spi
.include dff_x1.spi
.include nor4_x0.spi
.include inv_x0.spi
.include nor2_x0.spi
.include nexor2_x0.spi
.include or3_x1.spi
.include xor2_x0.spi
.include nor3_x0.spi
.include or4_x1.spi
.include diode_w1.spi

* Non-terminal models (part of the user's design hierarchy).

.subckt arlet6502_cts_r 0 1 23 83 1914 1918 1919 2074 2075 2076 2077 2078 2079 2080 2081 2082 2083 2084 2085 2086 2087 2088 2089 2090 2091 2092 2093 2094 2095 2096 2097 2098 2099 2100 2101 2102 2103 2104 2105 2106
* NET     0 = vss
* NET     1 = vdd
* NET     2 = reset_root_tr_tr_0
* NET     3 = reset_root_tr_tl_0
* NET     4 = reset_root_tr_br_0
* NET     5 = reset_root_tr_bl_0
* NET     6 = reset_root_tr_0
* NET     7 = reset_root_tl_tr_0
* NET     8 = reset_root_tl_tl_0
* NET     9 = reset_root_tl_br_0
* NET    10 = reset_root_tl_bl_0
* NET    11 = reset_root_tl_0
* NET    12 = reset_root_br_tr_0
* NET    13 = reset_root_br_tl_0
* NET    14 = reset_root_br_br_0
* NET    15 = reset_root_br_bl_0
* NET    16 = reset_root_br_0
* NET    17 = reset_root_bl_tr_0
* NET    18 = reset_root_bl_tl_0
* NET    19 = reset_root_bl_br_0
* NET    20 = reset_root_bl_bl_0
* NET    21 = reset_root_bl_0
* NET    22 = reset_root_0
* NET    23 = reset
* NET    24 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[5]
* NET    25 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[4]
* NET    26 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[3]
* NET    27 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[2]
* NET    28 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[1]
* NET    29 = flatten_MOS6502_auto_fsm_map_cc_288_map_fsm_1405_Y[0]
* NET    30 = clk_root_tr_tr_2
* NET    31 = clk_root_tr_tr_1
* NET    32 = clk_root_tr_tr_0
* NET    33 = clk_root_tr_tl_2
* NET    34 = clk_root_tr_tl_1
* NET    35 = clk_root_tr_tl_0
* NET    36 = clk_root_tr_br_2
* NET    37 = clk_root_tr_br_1
* NET    38 = clk_root_tr_br_0
* NET    39 = clk_root_tr_bl_2
* NET    40 = clk_root_tr_bl_1
* NET    41 = clk_root_tr_bl_0
* NET    42 = clk_root_tr_0
* NET    43 = clk_root_tl_tr_2
* NET    44 = clk_root_tl_tr_1
* NET    45 = clk_root_tl_tr_0
* NET    46 = clk_root_tl_tl_2
* NET    47 = clk_root_tl_tl_1
* NET    48 = clk_root_tl_tl_0
* NET    49 = clk_root_tl_br_2
* NET    50 = clk_root_tl_br_1
* NET    51 = clk_root_tl_br_0
* NET    52 = clk_root_tl_bl_2
* NET    53 = clk_root_tl_bl_1
* NET    54 = clk_root_tl_bl_0
* NET    55 = clk_root_tl_0
* NET    56 = clk_root_br_tr_2
* NET    57 = clk_root_br_tr_1
* NET    58 = clk_root_br_tr_0
* NET    59 = clk_root_br_tl_2
* NET    60 = clk_root_br_tl_1
* NET    61 = clk_root_br_tl_0
* NET    62 = clk_root_br_br_2
* NET    63 = clk_root_br_br_1
* NET    64 = clk_root_br_br_0
* NET    65 = clk_root_br_bl_2
* NET    66 = clk_root_br_bl_1
* NET    67 = clk_root_br_bl_0
* NET    68 = clk_root_br_0
* NET    69 = clk_root_bl_tr_2
* NET    70 = clk_root_bl_tr_1
* NET    71 = clk_root_bl_tr_0
* NET    72 = clk_root_bl_tl_2
* NET    73 = clk_root_bl_tl_1
* NET    74 = clk_root_bl_tl_0
* NET    75 = clk_root_bl_br_2
* NET    76 = clk_root_bl_br_1
* NET    77 = clk_root_bl_br_0
* NET    78 = clk_root_bl_bl_2
* NET    79 = clk_root_bl_bl_1
* NET    80 = clk_root_bl_bl_0
* NET    81 = clk_root_bl_0
* NET    82 = clk_root_0
* NET    83 = clk
* NET    84 = blockagenet
* NET    85 = abc_11867_new_n999
* NET    86 = abc_11867_new_n998
* NET    87 = abc_11867_new_n997
* NET    88 = abc_11867_new_n996
* NET    89 = abc_11867_new_n995
* NET    90 = abc_11867_new_n994
* NET    91 = abc_11867_new_n993
* NET    92 = abc_11867_new_n992
* NET    93 = abc_11867_new_n991
* NET    94 = abc_11867_new_n990
* NET    95 = abc_11867_new_n988
* NET    96 = abc_11867_new_n987
* NET    97 = abc_11867_new_n986
* NET    98 = abc_11867_new_n985
* NET    99 = abc_11867_new_n984
* NET   100 = abc_11867_new_n983
* NET   101 = abc_11867_new_n982
* NET   102 = abc_11867_new_n981
* NET   103 = abc_11867_new_n980
* NET   104 = abc_11867_new_n979
* NET   105 = abc_11867_new_n977
* NET   106 = abc_11867_new_n976
* NET   107 = abc_11867_new_n975
* NET   108 = abc_11867_new_n974
* NET   109 = abc_11867_new_n973
* NET   110 = abc_11867_new_n972
* NET   111 = abc_11867_new_n971
* NET   112 = abc_11867_new_n970
* NET   113 = abc_11867_new_n969
* NET   114 = abc_11867_new_n968
* NET   115 = abc_11867_new_n967
* NET   116 = abc_11867_new_n966
* NET   117 = abc_11867_new_n965
* NET   118 = abc_11867_new_n964
* NET   119 = abc_11867_new_n963
* NET   120 = abc_11867_new_n962
* NET   121 = abc_11867_new_n961
* NET   122 = abc_11867_new_n959
* NET   123 = abc_11867_new_n958
* NET   124 = abc_11867_new_n957
* NET   125 = abc_11867_new_n956
* NET   126 = abc_11867_new_n955
* NET   127 = abc_11867_new_n954
* NET   128 = abc_11867_new_n953
* NET   129 = abc_11867_new_n952
* NET   130 = abc_11867_new_n951
* NET   131 = abc_11867_new_n950
* NET   132 = abc_11867_new_n949
* NET   133 = abc_11867_new_n948
* NET   134 = abc_11867_new_n946
* NET   135 = abc_11867_new_n945
* NET   136 = abc_11867_new_n944
* NET   137 = abc_11867_new_n943
* NET   138 = abc_11867_new_n942
* NET   139 = abc_11867_new_n941
* NET   140 = abc_11867_new_n940
* NET   141 = abc_11867_new_n939
* NET   142 = abc_11867_new_n938
* NET   143 = abc_11867_new_n937
* NET   144 = abc_11867_new_n936
* NET   145 = abc_11867_new_n935
* NET   146 = abc_11867_new_n933
* NET   147 = abc_11867_new_n932
* NET   148 = abc_11867_new_n931
* NET   149 = abc_11867_new_n930
* NET   150 = abc_11867_new_n929
* NET   151 = abc_11867_new_n928
* NET   152 = abc_11867_new_n927
* NET   153 = abc_11867_new_n926
* NET   154 = abc_11867_new_n925
* NET   155 = abc_11867_new_n924
* NET   156 = abc_11867_new_n923
* NET   157 = abc_11867_new_n922
* NET   158 = abc_11867_new_n920
* NET   159 = abc_11867_new_n919
* NET   160 = abc_11867_new_n918
* NET   161 = abc_11867_new_n917
* NET   162 = abc_11867_new_n916
* NET   163 = abc_11867_new_n915
* NET   164 = abc_11867_new_n914
* NET   165 = abc_11867_new_n913
* NET   166 = abc_11867_new_n912
* NET   167 = abc_11867_new_n911
* NET   168 = abc_11867_new_n910
* NET   169 = abc_11867_new_n909
* NET   170 = abc_11867_new_n908
* NET   171 = abc_11867_new_n907
* NET   172 = abc_11867_new_n906
* NET   173 = abc_11867_new_n905
* NET   174 = abc_11867_new_n904
* NET   175 = abc_11867_new_n903
* NET   176 = abc_11867_new_n902
* NET   177 = abc_11867_new_n901
* NET   178 = abc_11867_new_n900
* NET   179 = abc_11867_new_n899
* NET   180 = abc_11867_new_n898
* NET   181 = abc_11867_new_n897
* NET   182 = abc_11867_new_n896
* NET   183 = abc_11867_new_n895
* NET   184 = abc_11867_new_n894
* NET   185 = abc_11867_new_n893
* NET   186 = abc_11867_new_n892
* NET   187 = abc_11867_new_n891
* NET   188 = abc_11867_new_n890
* NET   189 = abc_11867_new_n889
* NET   190 = abc_11867_new_n888
* NET   191 = abc_11867_new_n887
* NET   192 = abc_11867_new_n886
* NET   193 = abc_11867_new_n885
* NET   194 = abc_11867_new_n884
* NET   195 = abc_11867_new_n883
* NET   196 = abc_11867_new_n882
* NET   197 = abc_11867_new_n881
* NET   198 = abc_11867_new_n880
* NET   199 = abc_11867_new_n879
* NET   200 = abc_11867_new_n878
* NET   201 = abc_11867_new_n876
* NET   202 = abc_11867_new_n875
* NET   203 = abc_11867_new_n874
* NET   204 = abc_11867_new_n873
* NET   205 = abc_11867_new_n872
* NET   206 = abc_11867_new_n871
* NET   207 = abc_11867_new_n870
* NET   208 = abc_11867_new_n869
* NET   209 = abc_11867_new_n868
* NET   210 = abc_11867_new_n867
* NET   211 = abc_11867_new_n866
* NET   212 = abc_11867_new_n865
* NET   213 = abc_11867_new_n863
* NET   214 = abc_11867_new_n862
* NET   215 = abc_11867_new_n861
* NET   216 = abc_11867_new_n860
* NET   217 = abc_11867_new_n859
* NET   218 = abc_11867_new_n858
* NET   219 = abc_11867_new_n857
* NET   220 = abc_11867_new_n856
* NET   221 = abc_11867_new_n855
* NET   222 = abc_11867_new_n854
* NET   223 = abc_11867_new_n853
* NET   224 = abc_11867_new_n851
* NET   225 = abc_11867_new_n850
* NET   226 = abc_11867_new_n849
* NET   227 = abc_11867_new_n848
* NET   228 = abc_11867_new_n847
* NET   229 = abc_11867_new_n846
* NET   230 = abc_11867_new_n845
* NET   231 = abc_11867_new_n844
* NET   232 = abc_11867_new_n843
* NET   233 = abc_11867_new_n841
* NET   234 = abc_11867_new_n840
* NET   235 = abc_11867_new_n839
* NET   236 = abc_11867_new_n838
* NET   237 = abc_11867_new_n837
* NET   238 = abc_11867_new_n836
* NET   239 = abc_11867_new_n835
* NET   240 = abc_11867_new_n834
* NET   241 = abc_11867_new_n833
* NET   242 = abc_11867_new_n832
* NET   243 = abc_11867_new_n831
* NET   244 = abc_11867_new_n830
* NET   245 = abc_11867_new_n829
* NET   246 = abc_11867_new_n828
* NET   247 = abc_11867_new_n827
* NET   248 = abc_11867_new_n826
* NET   249 = abc_11867_new_n825
* NET   250 = abc_11867_new_n824
* NET   251 = abc_11867_new_n823
* NET   252 = abc_11867_new_n822
* NET   253 = abc_11867_new_n821
* NET   254 = abc_11867_new_n820
* NET   255 = abc_11867_new_n819
* NET   256 = abc_11867_new_n818
* NET   257 = abc_11867_new_n817
* NET   258 = abc_11867_new_n816
* NET   259 = abc_11867_new_n815
* NET   260 = abc_11867_new_n814
* NET   261 = abc_11867_new_n813
* NET   262 = abc_11867_new_n811
* NET   263 = abc_11867_new_n810
* NET   264 = abc_11867_new_n809
* NET   265 = abc_11867_new_n808
* NET   266 = abc_11867_new_n807
* NET   267 = abc_11867_new_n806
* NET   268 = abc_11867_new_n805
* NET   269 = abc_11867_new_n804
* NET   270 = abc_11867_new_n803
* NET   271 = abc_11867_new_n802
* NET   272 = abc_11867_new_n801
* NET   273 = abc_11867_new_n800
* NET   274 = abc_11867_new_n799
* NET   275 = abc_11867_new_n798
* NET   276 = abc_11867_new_n797
* NET   277 = abc_11867_new_n796
* NET   278 = abc_11867_new_n795
* NET   279 = abc_11867_new_n794
* NET   280 = abc_11867_new_n793
* NET   281 = abc_11867_new_n792
* NET   282 = abc_11867_new_n791
* NET   283 = abc_11867_new_n790
* NET   284 = abc_11867_new_n789
* NET   285 = abc_11867_new_n788
* NET   286 = abc_11867_new_n787
* NET   287 = abc_11867_new_n786
* NET   288 = abc_11867_new_n785
* NET   289 = abc_11867_new_n784
* NET   290 = abc_11867_new_n783
* NET   291 = abc_11867_new_n782
* NET   292 = abc_11867_new_n781
* NET   293 = abc_11867_new_n780
* NET   294 = abc_11867_new_n779
* NET   295 = abc_11867_new_n778
* NET   296 = abc_11867_new_n777
* NET   297 = abc_11867_new_n776
* NET   298 = abc_11867_new_n775
* NET   299 = abc_11867_new_n774
* NET   300 = abc_11867_new_n773
* NET   301 = abc_11867_new_n772
* NET   302 = abc_11867_new_n771
* NET   303 = abc_11867_new_n770
* NET   304 = abc_11867_new_n769
* NET   305 = abc_11867_new_n768
* NET   306 = abc_11867_new_n767
* NET   307 = abc_11867_new_n766
* NET   308 = abc_11867_new_n765
* NET   309 = abc_11867_new_n764
* NET   310 = abc_11867_new_n763
* NET   311 = abc_11867_new_n762
* NET   312 = abc_11867_new_n761
* NET   313 = abc_11867_new_n760
* NET   314 = abc_11867_new_n759
* NET   315 = abc_11867_new_n758
* NET   316 = abc_11867_new_n757
* NET   317 = abc_11867_new_n756
* NET   318 = abc_11867_new_n754
* NET   319 = abc_11867_new_n753
* NET   320 = abc_11867_new_n752
* NET   321 = abc_11867_new_n751
* NET   322 = abc_11867_new_n750
* NET   323 = abc_11867_new_n749
* NET   324 = abc_11867_new_n748
* NET   325 = abc_11867_new_n747
* NET   326 = abc_11867_new_n746
* NET   327 = abc_11867_new_n745
* NET   328 = abc_11867_new_n744
* NET   329 = abc_11867_new_n743
* NET   330 = abc_11867_new_n742
* NET   331 = abc_11867_new_n741
* NET   332 = abc_11867_new_n740
* NET   333 = abc_11867_new_n739
* NET   334 = abc_11867_new_n738
* NET   335 = abc_11867_new_n737
* NET   336 = abc_11867_new_n736
* NET   337 = abc_11867_new_n735
* NET   338 = abc_11867_new_n734
* NET   339 = abc_11867_new_n733
* NET   340 = abc_11867_new_n732
* NET   341 = abc_11867_new_n731
* NET   342 = abc_11867_new_n730
* NET   343 = abc_11867_new_n729
* NET   344 = abc_11867_new_n728
* NET   345 = abc_11867_new_n727
* NET   346 = abc_11867_new_n726
* NET   347 = abc_11867_new_n725
* NET   348 = abc_11867_new_n724
* NET   349 = abc_11867_new_n723
* NET   350 = abc_11867_new_n722
* NET   351 = abc_11867_new_n721
* NET   352 = abc_11867_new_n720
* NET   353 = abc_11867_new_n719
* NET   354 = abc_11867_new_n718
* NET   355 = abc_11867_new_n717
* NET   356 = abc_11867_new_n716
* NET   357 = abc_11867_new_n715
* NET   358 = abc_11867_new_n714
* NET   359 = abc_11867_new_n713
* NET   360 = abc_11867_new_n712
* NET   361 = abc_11867_new_n711
* NET   362 = abc_11867_new_n710
* NET   363 = abc_11867_new_n709
* NET   364 = abc_11867_new_n708
* NET   365 = abc_11867_new_n707
* NET   366 = abc_11867_new_n706
* NET   367 = abc_11867_new_n705
* NET   368 = abc_11867_new_n704
* NET   369 = abc_11867_new_n703
* NET   370 = abc_11867_new_n702
* NET   371 = abc_11867_new_n701
* NET   372 = abc_11867_new_n700
* NET   373 = abc_11867_new_n699
* NET   374 = abc_11867_new_n698
* NET   375 = abc_11867_new_n697
* NET   376 = abc_11867_new_n696
* NET   377 = abc_11867_new_n695
* NET   378 = abc_11867_new_n694
* NET   379 = abc_11867_new_n693
* NET   380 = abc_11867_new_n692
* NET   381 = abc_11867_new_n691
* NET   382 = abc_11867_new_n690
* NET   383 = abc_11867_new_n689
* NET   384 = abc_11867_new_n688
* NET   385 = abc_11867_new_n687
* NET   386 = abc_11867_new_n686
* NET   387 = abc_11867_new_n685
* NET   388 = abc_11867_new_n683
* NET   389 = abc_11867_new_n682
* NET   390 = abc_11867_new_n681
* NET   391 = abc_11867_new_n680
* NET   392 = abc_11867_new_n679
* NET   393 = abc_11867_new_n678
* NET   394 = abc_11867_new_n677
* NET   395 = abc_11867_new_n676
* NET   396 = abc_11867_new_n675
* NET   397 = abc_11867_new_n674
* NET   398 = abc_11867_new_n673
* NET   399 = abc_11867_new_n672
* NET   400 = abc_11867_new_n671
* NET   401 = abc_11867_new_n670
* NET   402 = abc_11867_new_n669
* NET   403 = abc_11867_new_n668
* NET   404 = abc_11867_new_n667
* NET   405 = abc_11867_new_n666
* NET   406 = abc_11867_new_n665
* NET   407 = abc_11867_new_n664
* NET   408 = abc_11867_new_n663
* NET   409 = abc_11867_new_n662
* NET   410 = abc_11867_new_n661
* NET   411 = abc_11867_new_n660
* NET   412 = abc_11867_new_n659
* NET   413 = abc_11867_new_n658
* NET   414 = abc_11867_new_n657
* NET   415 = abc_11867_new_n656
* NET   416 = abc_11867_new_n655
* NET   417 = abc_11867_new_n654
* NET   418 = abc_11867_new_n653
* NET   419 = abc_11867_new_n652
* NET   420 = abc_11867_new_n651
* NET   421 = abc_11867_new_n650
* NET   422 = abc_11867_new_n649
* NET   423 = abc_11867_new_n648
* NET   424 = abc_11867_new_n647
* NET   425 = abc_11867_new_n646
* NET   426 = abc_11867_new_n645
* NET   427 = abc_11867_new_n644
* NET   428 = abc_11867_new_n643
* NET   429 = abc_11867_new_n642
* NET   430 = abc_11867_new_n641
* NET   431 = abc_11867_new_n640
* NET   432 = abc_11867_new_n639
* NET   433 = abc_11867_new_n638
* NET   434 = abc_11867_new_n637
* NET   435 = abc_11867_new_n636
* NET   436 = abc_11867_new_n635
* NET   437 = abc_11867_new_n634
* NET   438 = abc_11867_new_n633
* NET   439 = abc_11867_new_n632
* NET   440 = abc_11867_new_n631
* NET   441 = abc_11867_new_n630
* NET   442 = abc_11867_new_n629
* NET   443 = abc_11867_new_n628
* NET   444 = abc_11867_new_n627
* NET   445 = abc_11867_new_n626
* NET   446 = abc_11867_new_n625
* NET   447 = abc_11867_new_n624
* NET   448 = abc_11867_new_n623
* NET   449 = abc_11867_new_n622
* NET   450 = abc_11867_new_n621
* NET   451 = abc_11867_new_n620
* NET   452 = abc_11867_new_n619
* NET   453 = abc_11867_new_n618
* NET   454 = abc_11867_new_n617
* NET   455 = abc_11867_new_n616
* NET   456 = abc_11867_new_n615
* NET   457 = abc_11867_new_n614
* NET   458 = abc_11867_new_n613
* NET   459 = abc_11867_new_n612
* NET   460 = abc_11867_new_n611
* NET   461 = abc_11867_new_n610
* NET   462 = abc_11867_new_n609
* NET   463 = abc_11867_new_n608
* NET   464 = abc_11867_new_n607
* NET   465 = abc_11867_new_n606
* NET   466 = abc_11867_new_n605
* NET   467 = abc_11867_new_n604
* NET   468 = abc_11867_new_n603
* NET   469 = abc_11867_new_n602
* NET   470 = abc_11867_new_n601
* NET   471 = abc_11867_new_n600
* NET   472 = abc_11867_new_n599
* NET   473 = abc_11867_new_n598
* NET   474 = abc_11867_new_n597
* NET   475 = abc_11867_new_n596
* NET   476 = abc_11867_new_n595
* NET   477 = abc_11867_new_n594
* NET   478 = abc_11867_new_n593
* NET   479 = abc_11867_new_n592
* NET   480 = abc_11867_new_n591
* NET   481 = abc_11867_new_n590
* NET   482 = abc_11867_new_n589
* NET   483 = abc_11867_new_n588
* NET   484 = abc_11867_new_n587
* NET   485 = abc_11867_new_n586
* NET   486 = abc_11867_new_n585
* NET   487 = abc_11867_new_n584
* NET   488 = abc_11867_new_n583_hfns_2
* NET   489 = abc_11867_new_n583_hfns_1
* NET   490 = abc_11867_new_n583_hfns_0
* NET   491 = abc_11867_new_n583
* NET   492 = abc_11867_new_n582
* NET   493 = abc_11867_new_n581
* NET   494 = abc_11867_new_n580
* NET   495 = abc_11867_new_n579
* NET   496 = abc_11867_new_n578
* NET   497 = abc_11867_new_n577
* NET   498 = abc_11867_new_n576
* NET   499 = abc_11867_new_n575
* NET   500 = abc_11867_new_n574
* NET   501 = abc_11867_new_n573
* NET   502 = abc_11867_new_n572
* NET   503 = abc_11867_new_n571
* NET   504 = abc_11867_new_n570
* NET   505 = abc_11867_new_n569
* NET   506 = abc_11867_new_n568
* NET   507 = abc_11867_new_n567
* NET   508 = abc_11867_new_n566
* NET   509 = abc_11867_new_n565
* NET   510 = abc_11867_new_n564
* NET   511 = abc_11867_new_n563
* NET   512 = abc_11867_new_n562
* NET   513 = abc_11867_new_n561
* NET   514 = abc_11867_new_n560
* NET   515 = abc_11867_new_n559
* NET   516 = abc_11867_new_n558
* NET   517 = abc_11867_new_n557
* NET   518 = abc_11867_new_n556
* NET   519 = abc_11867_new_n555
* NET   520 = abc_11867_new_n554
* NET   521 = abc_11867_new_n553
* NET   522 = abc_11867_new_n552
* NET   523 = abc_11867_new_n551
* NET   524 = abc_11867_new_n550
* NET   525 = abc_11867_new_n549
* NET   526 = abc_11867_new_n548
* NET   527 = abc_11867_new_n547
* NET   528 = abc_11867_new_n546
* NET   529 = abc_11867_new_n545
* NET   530 = abc_11867_new_n544
* NET   531 = abc_11867_new_n543_hfns_2
* NET   532 = abc_11867_new_n543_hfns_1
* NET   533 = abc_11867_new_n543_hfns_0
* NET   534 = abc_11867_new_n543
* NET   535 = abc_11867_new_n542
* NET   536 = abc_11867_new_n541
* NET   537 = abc_11867_new_n540
* NET   538 = abc_11867_new_n539
* NET   539 = abc_11867_new_n538
* NET   540 = abc_11867_new_n537
* NET   541 = abc_11867_new_n536
* NET   542 = abc_11867_new_n535
* NET   543 = abc_11867_new_n534
* NET   544 = abc_11867_new_n533
* NET   545 = abc_11867_new_n532
* NET   546 = abc_11867_new_n531
* NET   547 = abc_11867_new_n530
* NET   548 = abc_11867_new_n529
* NET   549 = abc_11867_new_n528
* NET   550 = abc_11867_new_n527
* NET   551 = abc_11867_new_n526
* NET   552 = abc_11867_new_n525
* NET   553 = abc_11867_new_n524
* NET   554 = abc_11867_new_n523
* NET   555 = abc_11867_new_n522_hfns_3
* NET   556 = abc_11867_new_n522_hfns_2
* NET   557 = abc_11867_new_n522_hfns_1
* NET   558 = abc_11867_new_n522_hfns_0
* NET   559 = abc_11867_new_n522
* NET   560 = abc_11867_new_n521
* NET   561 = abc_11867_new_n520
* NET   562 = abc_11867_new_n519
* NET   563 = abc_11867_new_n518
* NET   564 = abc_11867_new_n517
* NET   565 = abc_11867_new_n516
* NET   566 = abc_11867_new_n515
* NET   567 = abc_11867_new_n514
* NET   568 = abc_11867_new_n513
* NET   569 = abc_11867_new_n512
* NET   570 = abc_11867_new_n511
* NET   571 = abc_11867_new_n510
* NET   572 = abc_11867_new_n509
* NET   573 = abc_11867_new_n508
* NET   574 = abc_11867_new_n507
* NET   575 = abc_11867_new_n506
* NET   576 = abc_11867_new_n505
* NET   577 = abc_11867_new_n504
* NET   578 = abc_11867_new_n503
* NET   579 = abc_11867_new_n502
* NET   580 = abc_11867_new_n501
* NET   581 = abc_11867_new_n500
* NET   582 = abc_11867_new_n499
* NET   583 = abc_11867_new_n498
* NET   584 = abc_11867_new_n497
* NET   585 = abc_11867_new_n496
* NET   586 = abc_11867_new_n495
* NET   587 = abc_11867_new_n494
* NET   588 = abc_11867_new_n493
* NET   589 = abc_11867_new_n492
* NET   590 = abc_11867_new_n491
* NET   591 = abc_11867_new_n490
* NET   592 = abc_11867_new_n489
* NET   593 = abc_11867_new_n488_hfns_2
* NET   594 = abc_11867_new_n488_hfns_1
* NET   595 = abc_11867_new_n488_hfns_0
* NET   596 = abc_11867_new_n488
* NET   597 = abc_11867_new_n487
* NET   598 = abc_11867_new_n486
* NET   599 = abc_11867_new_n485
* NET   600 = abc_11867_new_n484
* NET   601 = abc_11867_new_n483
* NET   602 = abc_11867_new_n482
* NET   603 = abc_11867_new_n481
* NET   604 = abc_11867_new_n480
* NET   605 = abc_11867_new_n479
* NET   606 = abc_11867_new_n478
* NET   607 = abc_11867_new_n477_hfns_3
* NET   608 = abc_11867_new_n477_hfns_2
* NET   609 = abc_11867_new_n477_hfns_1
* NET   610 = abc_11867_new_n477_hfns_0
* NET   611 = abc_11867_new_n477
* NET   612 = abc_11867_new_n476
* NET   613 = abc_11867_new_n475
* NET   614 = abc_11867_new_n474
* NET   615 = abc_11867_new_n473_hfns_2
* NET   616 = abc_11867_new_n473_hfns_1
* NET   617 = abc_11867_new_n473_hfns_0
* NET   618 = abc_11867_new_n473
* NET   619 = abc_11867_new_n472
* NET   620 = abc_11867_new_n471
* NET   621 = abc_11867_new_n470
* NET   622 = abc_11867_new_n469
* NET   623 = abc_11867_new_n468
* NET   624 = abc_11867_new_n467
* NET   625 = abc_11867_new_n466
* NET   626 = abc_11867_new_n465
* NET   627 = abc_11867_new_n464
* NET   628 = abc_11867_new_n463
* NET   629 = abc_11867_new_n462
* NET   630 = abc_11867_new_n461
* NET   631 = abc_11867_new_n460
* NET   632 = abc_11867_new_n459
* NET   633 = abc_11867_new_n458
* NET   634 = abc_11867_new_n457
* NET   635 = abc_11867_new_n456
* NET   636 = abc_11867_new_n455
* NET   637 = abc_11867_new_n454
* NET   638 = abc_11867_new_n453
* NET   639 = abc_11867_new_n452
* NET   640 = abc_11867_new_n451
* NET   641 = abc_11867_new_n450
* NET   642 = abc_11867_new_n449
* NET   643 = abc_11867_new_n448
* NET   644 = abc_11867_new_n447
* NET   645 = abc_11867_new_n446
* NET   646 = abc_11867_new_n445
* NET   647 = abc_11867_new_n444
* NET   648 = abc_11867_new_n443
* NET   649 = abc_11867_new_n442
* NET   650 = abc_11867_new_n441
* NET   651 = abc_11867_new_n440
* NET   652 = abc_11867_new_n439
* NET   653 = abc_11867_new_n438
* NET   654 = abc_11867_new_n437
* NET   655 = abc_11867_new_n436
* NET   656 = abc_11867_new_n435
* NET   657 = abc_11867_new_n434
* NET   658 = abc_11867_new_n433_hfns_3
* NET   659 = abc_11867_new_n433_hfns_2
* NET   660 = abc_11867_new_n433_hfns_1
* NET   661 = abc_11867_new_n433_hfns_0
* NET   662 = abc_11867_new_n433
* NET   663 = abc_11867_new_n432
* NET   664 = abc_11867_new_n431_hfns_2
* NET   665 = abc_11867_new_n431_hfns_1
* NET   666 = abc_11867_new_n431_hfns_0
* NET   667 = abc_11867_new_n431
* NET   668 = abc_11867_new_n430_hfns_2
* NET   669 = abc_11867_new_n430_hfns_1
* NET   670 = abc_11867_new_n430_hfns_0
* NET   671 = abc_11867_new_n430
* NET   672 = abc_11867_new_n429_hfns_2
* NET   673 = abc_11867_new_n429_hfns_1
* NET   674 = abc_11867_new_n429_hfns_0
* NET   675 = abc_11867_new_n429
* NET   676 = abc_11867_new_n428
* NET   677 = abc_11867_new_n427_hfns_5
* NET   678 = abc_11867_new_n427_hfns_4
* NET   679 = abc_11867_new_n427_hfns_3
* NET   680 = abc_11867_new_n427_hfns_2
* NET   681 = abc_11867_new_n427_hfns_1
* NET   682 = abc_11867_new_n427_hfns_0
* NET   683 = abc_11867_new_n427
* NET   684 = abc_11867_new_n426
* NET   685 = abc_11867_new_n425_hfns_2
* NET   686 = abc_11867_new_n425_hfns_1
* NET   687 = abc_11867_new_n425_hfns_0
* NET   688 = abc_11867_new_n425
* NET   689 = abc_11867_new_n423
* NET   690 = abc_11867_new_n421
* NET   691 = abc_11867_new_n419
* NET   692 = abc_11867_new_n417
* NET   693 = abc_11867_new_n415
* NET   694 = abc_11867_new_n413
* NET   695 = abc_11867_new_n411
* NET   696 = abc_11867_new_n409
* NET   697 = abc_11867_new_n408
* NET   698 = abc_11867_new_n407
* NET   699 = abc_11867_new_n406
* NET   700 = abc_11867_new_n405
* NET   701 = abc_11867_new_n404
* NET   702 = abc_11867_new_n403
* NET   703 = abc_11867_new_n402
* NET   704 = abc_11867_new_n401
* NET   705 = abc_11867_new_n400
* NET   706 = abc_11867_new_n399
* NET   707 = abc_11867_new_n398
* NET   708 = abc_11867_new_n397
* NET   709 = abc_11867_new_n396
* NET   710 = abc_11867_new_n395
* NET   711 = abc_11867_new_n394
* NET   712 = abc_11867_new_n393
* NET   713 = abc_11867_new_n392
* NET   714 = abc_11867_new_n391
* NET   715 = abc_11867_new_n390
* NET   716 = abc_11867_new_n389
* NET   717 = abc_11867_new_n388
* NET   718 = abc_11867_new_n387
* NET   719 = abc_11867_new_n386
* NET   720 = abc_11867_new_n385
* NET   721 = abc_11867_new_n384
* NET   722 = abc_11867_new_n383
* NET   723 = abc_11867_new_n382
* NET   724 = abc_11867_new_n381
* NET   725 = abc_11867_new_n380
* NET   726 = abc_11867_new_n379
* NET   727 = abc_11867_new_n378
* NET   728 = abc_11867_new_n377
* NET   729 = abc_11867_new_n376
* NET   730 = abc_11867_new_n375
* NET   731 = abc_11867_new_n374
* NET   732 = abc_11867_new_n373
* NET   733 = abc_11867_new_n372
* NET   734 = abc_11867_new_n371
* NET   735 = abc_11867_new_n370
* NET   736 = abc_11867_new_n369
* NET   737 = abc_11867_new_n368
* NET   738 = abc_11867_new_n367
* NET   739 = abc_11867_new_n366
* NET   740 = abc_11867_new_n365
* NET   741 = abc_11867_new_n364
* NET   742 = abc_11867_new_n363
* NET   743 = abc_11867_new_n362
* NET   744 = abc_11867_new_n361
* NET   745 = abc_11867_new_n360
* NET   746 = abc_11867_new_n359
* NET   747 = abc_11867_new_n358
* NET   748 = abc_11867_new_n357
* NET   749 = abc_11867_new_n356
* NET   750 = abc_11867_new_n355
* NET   751 = abc_11867_new_n354
* NET   752 = abc_11867_new_n353
* NET   753 = abc_11867_new_n352
* NET   754 = abc_11867_new_n351
* NET   755 = abc_11867_new_n350
* NET   756 = abc_11867_new_n349
* NET   757 = abc_11867_new_n348
* NET   758 = abc_11867_new_n347
* NET   759 = abc_11867_new_n346
* NET   760 = abc_11867_new_n345
* NET   761 = abc_11867_new_n344
* NET   762 = abc_11867_new_n343
* NET   763 = abc_11867_new_n342
* NET   764 = abc_11867_new_n341
* NET   765 = abc_11867_new_n340
* NET   766 = abc_11867_new_n339
* NET   767 = abc_11867_new_n338
* NET   768 = abc_11867_new_n337
* NET   769 = abc_11867_new_n336
* NET   770 = abc_11867_new_n335
* NET   771 = abc_11867_new_n334
* NET   772 = abc_11867_new_n333_hfns_3
* NET   773 = abc_11867_new_n333_hfns_2
* NET   774 = abc_11867_new_n333_hfns_1
* NET   775 = abc_11867_new_n333_hfns_0
* NET   776 = abc_11867_new_n333
* NET   777 = abc_11867_new_n332
* NET   778 = abc_11867_new_n331
* NET   779 = abc_11867_new_n330
* NET   780 = abc_11867_new_n329
* NET   781 = abc_11867_new_n328
* NET   782 = abc_11867_new_n327
* NET   783 = abc_11867_new_n326
* NET   784 = abc_11867_new_n325
* NET   785 = abc_11867_new_n324
* NET   786 = abc_11867_new_n323
* NET   787 = abc_11867_new_n2135
* NET   788 = abc_11867_new_n2134
* NET   789 = abc_11867_new_n2133
* NET   790 = abc_11867_new_n2128
* NET   791 = abc_11867_new_n2127
* NET   792 = abc_11867_new_n2126
* NET   793 = abc_11867_new_n2124
* NET   794 = abc_11867_new_n2123
* NET   795 = abc_11867_new_n2122
* NET   796 = abc_11867_new_n2121
* NET   797 = abc_11867_new_n2120
* NET   798 = abc_11867_new_n2119
* NET   799 = abc_11867_new_n2118
* NET   800 = abc_11867_new_n2117
* NET   801 = abc_11867_new_n2116
* NET   802 = abc_11867_new_n2115
* NET   803 = abc_11867_new_n2114
* NET   804 = abc_11867_new_n2113
* NET   805 = abc_11867_new_n2112
* NET   806 = abc_11867_new_n2111
* NET   807 = abc_11867_new_n2110
* NET   808 = abc_11867_new_n2109
* NET   809 = abc_11867_new_n2108
* NET   810 = abc_11867_new_n2107
* NET   811 = abc_11867_new_n2106
* NET   812 = abc_11867_new_n2105
* NET   813 = abc_11867_new_n2104
* NET   814 = abc_11867_new_n2103
* NET   815 = abc_11867_new_n2102
* NET   816 = abc_11867_new_n2101
* NET   817 = abc_11867_new_n2100
* NET   818 = abc_11867_new_n2099
* NET   819 = abc_11867_new_n2098
* NET   820 = abc_11867_new_n2097
* NET   821 = abc_11867_new_n2096
* NET   822 = abc_11867_new_n2095
* NET   823 = abc_11867_new_n2094
* NET   824 = abc_11867_new_n2093
* NET   825 = abc_11867_new_n2092
* NET   826 = abc_11867_new_n2091
* NET   827 = abc_11867_new_n2090
* NET   828 = abc_11867_new_n2089
* NET   829 = abc_11867_new_n2088
* NET   830 = abc_11867_new_n2087
* NET   831 = abc_11867_new_n2086
* NET   832 = abc_11867_new_n2085
* NET   833 = abc_11867_new_n2084
* NET   834 = abc_11867_new_n2083
* NET   835 = abc_11867_new_n2082
* NET   836 = abc_11867_new_n2081
* NET   837 = abc_11867_new_n2080
* NET   838 = abc_11867_new_n2079
* NET   839 = abc_11867_new_n2078
* NET   840 = abc_11867_new_n2077
* NET   841 = abc_11867_new_n2076
* NET   842 = abc_11867_new_n2075
* NET   843 = abc_11867_new_n2074
* NET   844 = abc_11867_new_n2073
* NET   845 = abc_11867_new_n2072
* NET   846 = abc_11867_new_n2071
* NET   847 = abc_11867_new_n2070
* NET   848 = abc_11867_new_n2069
* NET   849 = abc_11867_new_n2068
* NET   850 = abc_11867_new_n2067
* NET   851 = abc_11867_new_n2066
* NET   852 = abc_11867_new_n2065
* NET   853 = abc_11867_new_n2064
* NET   854 = abc_11867_new_n2063
* NET   855 = abc_11867_new_n2062
* NET   856 = abc_11867_new_n2061
* NET   857 = abc_11867_new_n2060
* NET   858 = abc_11867_new_n2059
* NET   859 = abc_11867_new_n2058
* NET   860 = abc_11867_new_n2057
* NET   861 = abc_11867_new_n2056
* NET   862 = abc_11867_new_n2055
* NET   863 = abc_11867_new_n2054
* NET   864 = abc_11867_new_n2053
* NET   865 = abc_11867_new_n2052
* NET   866 = abc_11867_new_n2051
* NET   867 = abc_11867_new_n2050
* NET   868 = abc_11867_new_n2049
* NET   869 = abc_11867_new_n2048
* NET   870 = abc_11867_new_n2047
* NET   871 = abc_11867_new_n2046
* NET   872 = abc_11867_new_n2045
* NET   873 = abc_11867_new_n2044
* NET   874 = abc_11867_new_n2043
* NET   875 = abc_11867_new_n2042
* NET   876 = abc_11867_new_n2041
* NET   877 = abc_11867_new_n2040
* NET   878 = abc_11867_new_n2039
* NET   879 = abc_11867_new_n2038
* NET   880 = abc_11867_new_n2037
* NET   881 = abc_11867_new_n2036
* NET   882 = abc_11867_new_n2035
* NET   883 = abc_11867_new_n2034
* NET   884 = abc_11867_new_n2033
* NET   885 = abc_11867_new_n2032
* NET   886 = abc_11867_new_n2031
* NET   887 = abc_11867_new_n2030
* NET   888 = abc_11867_new_n2029
* NET   889 = abc_11867_new_n2028
* NET   890 = abc_11867_new_n2027
* NET   891 = abc_11867_new_n2026
* NET   892 = abc_11867_new_n2025
* NET   893 = abc_11867_new_n2024
* NET   894 = abc_11867_new_n2023
* NET   895 = abc_11867_new_n2022
* NET   896 = abc_11867_new_n2021
* NET   897 = abc_11867_new_n2020
* NET   898 = abc_11867_new_n2019
* NET   899 = abc_11867_new_n2018
* NET   900 = abc_11867_new_n2017
* NET   901 = abc_11867_new_n2016
* NET   902 = abc_11867_new_n2015
* NET   903 = abc_11867_new_n2014
* NET   904 = abc_11867_new_n2013
* NET   905 = abc_11867_new_n2012
* NET   906 = abc_11867_new_n2011
* NET   907 = abc_11867_new_n2010
* NET   908 = abc_11867_new_n2009
* NET   909 = abc_11867_new_n2008
* NET   910 = abc_11867_new_n2007
* NET   911 = abc_11867_new_n2006
* NET   912 = abc_11867_new_n2005
* NET   913 = abc_11867_new_n2004
* NET   914 = abc_11867_new_n2003
* NET   915 = abc_11867_new_n2002
* NET   916 = abc_11867_new_n2001
* NET   917 = abc_11867_new_n2000
* NET   918 = abc_11867_new_n1999
* NET   919 = abc_11867_new_n1998
* NET   920 = abc_11867_new_n1997
* NET   921 = abc_11867_new_n1996
* NET   922 = abc_11867_new_n1995
* NET   923 = abc_11867_new_n1994
* NET   924 = abc_11867_new_n1993
* NET   925 = abc_11867_new_n1992
* NET   926 = abc_11867_new_n1991
* NET   927 = abc_11867_new_n1990
* NET   928 = abc_11867_new_n1989
* NET   929 = abc_11867_new_n1988
* NET   930 = abc_11867_new_n1987
* NET   931 = abc_11867_new_n1986
* NET   932 = abc_11867_new_n1985
* NET   933 = abc_11867_new_n1984
* NET   934 = abc_11867_new_n1983
* NET   935 = abc_11867_new_n1982
* NET   936 = abc_11867_new_n1981
* NET   937 = abc_11867_new_n1980
* NET   938 = abc_11867_new_n1979
* NET   939 = abc_11867_new_n1978
* NET   940 = abc_11867_new_n1977
* NET   941 = abc_11867_new_n1976
* NET   942 = abc_11867_new_n1975
* NET   943 = abc_11867_new_n1974
* NET   944 = abc_11867_new_n1973
* NET   945 = abc_11867_new_n1972
* NET   946 = abc_11867_new_n1971
* NET   947 = abc_11867_new_n1970
* NET   948 = abc_11867_new_n1969
* NET   949 = abc_11867_new_n1968
* NET   950 = abc_11867_new_n1967
* NET   951 = abc_11867_new_n1966
* NET   952 = abc_11867_new_n1965
* NET   953 = abc_11867_new_n1964
* NET   954 = abc_11867_new_n1963
* NET   955 = abc_11867_new_n1962
* NET   956 = abc_11867_new_n1961
* NET   957 = abc_11867_new_n1960
* NET   958 = abc_11867_new_n1959
* NET   959 = abc_11867_new_n1958
* NET   960 = abc_11867_new_n1957
* NET   961 = abc_11867_new_n1956
* NET   962 = abc_11867_new_n1955
* NET   963 = abc_11867_new_n1954
* NET   964 = abc_11867_new_n1953
* NET   965 = abc_11867_new_n1952
* NET   966 = abc_11867_new_n1951
* NET   967 = abc_11867_new_n1950
* NET   968 = abc_11867_new_n1949
* NET   969 = abc_11867_new_n1948
* NET   970 = abc_11867_new_n1947
* NET   971 = abc_11867_new_n1946
* NET   972 = abc_11867_new_n1945
* NET   973 = abc_11867_new_n1944
* NET   974 = abc_11867_new_n1943
* NET   975 = abc_11867_new_n1942
* NET   976 = abc_11867_new_n1941
* NET   977 = abc_11867_new_n1940
* NET   978 = abc_11867_new_n1939
* NET   979 = abc_11867_new_n1938
* NET   980 = abc_11867_new_n1937
* NET   981 = abc_11867_new_n1936
* NET   982 = abc_11867_new_n1935
* NET   983 = abc_11867_new_n1934
* NET   984 = abc_11867_new_n1933
* NET   985 = abc_11867_new_n1932
* NET   986 = abc_11867_new_n1931
* NET   987 = abc_11867_new_n1930
* NET   988 = abc_11867_new_n1929
* NET   989 = abc_11867_new_n1928
* NET   990 = abc_11867_new_n1927
* NET   991 = abc_11867_new_n1926
* NET   992 = abc_11867_new_n1925
* NET   993 = abc_11867_new_n1924
* NET   994 = abc_11867_new_n1923
* NET   995 = abc_11867_new_n1922
* NET   996 = abc_11867_new_n1921
* NET   997 = abc_11867_new_n1920
* NET   998 = abc_11867_new_n1919
* NET   999 = abc_11867_new_n1918
* NET  1000 = abc_11867_new_n1917
* NET  1001 = abc_11867_new_n1916
* NET  1002 = abc_11867_new_n1915
* NET  1003 = abc_11867_new_n1914
* NET  1004 = abc_11867_new_n1913
* NET  1005 = abc_11867_new_n1912
* NET  1006 = abc_11867_new_n1911
* NET  1007 = abc_11867_new_n1910
* NET  1008 = abc_11867_new_n1909
* NET  1009 = abc_11867_new_n1908
* NET  1010 = abc_11867_new_n1907
* NET  1011 = abc_11867_new_n1906
* NET  1012 = abc_11867_new_n1905
* NET  1013 = abc_11867_new_n1904
* NET  1014 = abc_11867_new_n1903
* NET  1015 = abc_11867_new_n1902
* NET  1016 = abc_11867_new_n1901
* NET  1017 = abc_11867_new_n1900
* NET  1018 = abc_11867_new_n1899
* NET  1019 = abc_11867_new_n1898
* NET  1020 = abc_11867_new_n1897
* NET  1021 = abc_11867_new_n1896
* NET  1022 = abc_11867_new_n1895
* NET  1023 = abc_11867_new_n1894
* NET  1024 = abc_11867_new_n1893
* NET  1025 = abc_11867_new_n1892
* NET  1026 = abc_11867_new_n1891
* NET  1027 = abc_11867_new_n1890
* NET  1028 = abc_11867_new_n1889
* NET  1029 = abc_11867_new_n1888
* NET  1030 = abc_11867_new_n1887
* NET  1031 = abc_11867_new_n1886
* NET  1032 = abc_11867_new_n1885
* NET  1033 = abc_11867_new_n1884
* NET  1034 = abc_11867_new_n1883
* NET  1035 = abc_11867_new_n1882
* NET  1036 = abc_11867_new_n1881
* NET  1037 = abc_11867_new_n1880
* NET  1038 = abc_11867_new_n1879
* NET  1039 = abc_11867_new_n1878
* NET  1040 = abc_11867_new_n1877
* NET  1041 = abc_11867_new_n1876
* NET  1042 = abc_11867_new_n1875
* NET  1043 = abc_11867_new_n1874
* NET  1044 = abc_11867_new_n1873
* NET  1045 = abc_11867_new_n1872
* NET  1046 = abc_11867_new_n1871
* NET  1047 = abc_11867_new_n1870
* NET  1048 = abc_11867_new_n1869
* NET  1049 = abc_11867_new_n1868
* NET  1050 = abc_11867_new_n1867
* NET  1051 = abc_11867_new_n1866
* NET  1052 = abc_11867_new_n1865
* NET  1053 = abc_11867_new_n1864
* NET  1054 = abc_11867_new_n1863
* NET  1055 = abc_11867_new_n1862
* NET  1056 = abc_11867_new_n1861
* NET  1057 = abc_11867_new_n1860
* NET  1058 = abc_11867_new_n1859
* NET  1059 = abc_11867_new_n1858
* NET  1060 = abc_11867_new_n1857
* NET  1061 = abc_11867_new_n1856
* NET  1062 = abc_11867_new_n1854
* NET  1063 = abc_11867_new_n1853
* NET  1064 = abc_11867_new_n1852
* NET  1065 = abc_11867_new_n1851
* NET  1066 = abc_11867_new_n1850
* NET  1067 = abc_11867_new_n1849
* NET  1068 = abc_11867_new_n1848_hfns_2
* NET  1069 = abc_11867_new_n1848_hfns_1
* NET  1070 = abc_11867_new_n1848_hfns_0
* NET  1071 = abc_11867_new_n1848
* NET  1072 = abc_11867_new_n1847
* NET  1073 = abc_11867_new_n1846
* NET  1074 = abc_11867_new_n1845
* NET  1075 = abc_11867_new_n1844
* NET  1076 = abc_11867_new_n1843
* NET  1077 = abc_11867_new_n1842
* NET  1078 = abc_11867_new_n1841
* NET  1079 = abc_11867_new_n1840
* NET  1080 = abc_11867_new_n1839
* NET  1081 = abc_11867_new_n1838
* NET  1082 = abc_11867_new_n1837
* NET  1083 = abc_11867_new_n1836
* NET  1084 = abc_11867_new_n1835
* NET  1085 = abc_11867_new_n1834
* NET  1086 = abc_11867_new_n1833
* NET  1087 = abc_11867_new_n1832
* NET  1088 = abc_11867_new_n1831
* NET  1089 = abc_11867_new_n1830
* NET  1090 = abc_11867_new_n1829
* NET  1091 = abc_11867_new_n1828
* NET  1092 = abc_11867_new_n1827
* NET  1093 = abc_11867_new_n1826
* NET  1094 = abc_11867_new_n1825
* NET  1095 = abc_11867_new_n1824
* NET  1096 = abc_11867_new_n1823
* NET  1097 = abc_11867_new_n1822
* NET  1098 = abc_11867_new_n1821
* NET  1099 = abc_11867_new_n1820
* NET  1100 = abc_11867_new_n1819
* NET  1101 = abc_11867_new_n1818
* NET  1102 = abc_11867_new_n1817
* NET  1103 = abc_11867_new_n1816
* NET  1104 = abc_11867_new_n1815
* NET  1105 = abc_11867_new_n1814
* NET  1106 = abc_11867_new_n1813
* NET  1107 = abc_11867_new_n1812
* NET  1108 = abc_11867_new_n1811
* NET  1109 = abc_11867_new_n1810
* NET  1110 = abc_11867_new_n1809
* NET  1111 = abc_11867_new_n1808
* NET  1112 = abc_11867_new_n1807
* NET  1113 = abc_11867_new_n1806
* NET  1114 = abc_11867_new_n1805
* NET  1115 = abc_11867_new_n1804
* NET  1116 = abc_11867_new_n1803
* NET  1117 = abc_11867_new_n1802
* NET  1118 = abc_11867_new_n1801
* NET  1119 = abc_11867_new_n1800
* NET  1120 = abc_11867_new_n1799
* NET  1121 = abc_11867_new_n1798
* NET  1122 = abc_11867_new_n1797
* NET  1123 = abc_11867_new_n1796
* NET  1124 = abc_11867_new_n1795
* NET  1125 = abc_11867_new_n1794
* NET  1126 = abc_11867_new_n1793
* NET  1127 = abc_11867_new_n1792
* NET  1128 = abc_11867_new_n1791
* NET  1129 = abc_11867_new_n1790
* NET  1130 = abc_11867_new_n1789
* NET  1131 = abc_11867_new_n1788
* NET  1132 = abc_11867_new_n1787
* NET  1133 = abc_11867_new_n1786
* NET  1134 = abc_11867_new_n1785
* NET  1135 = abc_11867_new_n1784
* NET  1136 = abc_11867_new_n1783
* NET  1137 = abc_11867_new_n1782
* NET  1138 = abc_11867_new_n1781
* NET  1139 = abc_11867_new_n1780
* NET  1140 = abc_11867_new_n1779
* NET  1141 = abc_11867_new_n1778
* NET  1142 = abc_11867_new_n1777
* NET  1143 = abc_11867_new_n1776
* NET  1144 = abc_11867_new_n1775
* NET  1145 = abc_11867_new_n1773
* NET  1146 = abc_11867_new_n1772
* NET  1147 = abc_11867_new_n1771
* NET  1148 = abc_11867_new_n1770
* NET  1149 = abc_11867_new_n1769
* NET  1150 = abc_11867_new_n1768
* NET  1151 = abc_11867_new_n1767
* NET  1152 = abc_11867_new_n1766
* NET  1153 = abc_11867_new_n1765
* NET  1154 = abc_11867_new_n1764
* NET  1155 = abc_11867_new_n1763
* NET  1156 = abc_11867_new_n1761
* NET  1157 = abc_11867_new_n1760
* NET  1158 = abc_11867_new_n1759
* NET  1159 = abc_11867_new_n1758
* NET  1160 = abc_11867_new_n1757
* NET  1161 = abc_11867_new_n1756
* NET  1162 = abc_11867_new_n1755
* NET  1163 = abc_11867_new_n1754
* NET  1164 = abc_11867_new_n1753
* NET  1165 = abc_11867_new_n1752
* NET  1166 = abc_11867_new_n1751
* NET  1167 = abc_11867_new_n1749
* NET  1168 = abc_11867_new_n1748
* NET  1169 = abc_11867_new_n1747
* NET  1170 = abc_11867_new_n1746
* NET  1171 = abc_11867_new_n1745
* NET  1172 = abc_11867_new_n1744
* NET  1173 = abc_11867_new_n1743
* NET  1174 = abc_11867_new_n1742
* NET  1175 = abc_11867_new_n1741
* NET  1176 = abc_11867_new_n1740
* NET  1177 = abc_11867_new_n1739
* NET  1178 = abc_11867_new_n1738
* NET  1179 = abc_11867_new_n1737
* NET  1180 = abc_11867_new_n1735
* NET  1181 = abc_11867_new_n1734
* NET  1182 = abc_11867_new_n1733
* NET  1183 = abc_11867_new_n1732
* NET  1184 = abc_11867_new_n1731
* NET  1185 = abc_11867_new_n1730
* NET  1186 = abc_11867_new_n1729
* NET  1187 = abc_11867_new_n1728
* NET  1188 = abc_11867_new_n1727
* NET  1189 = abc_11867_new_n1726
* NET  1190 = abc_11867_new_n1725
* NET  1191 = abc_11867_new_n1724
* NET  1192 = abc_11867_new_n1723
* NET  1193 = abc_11867_new_n1721
* NET  1194 = abc_11867_new_n1720
* NET  1195 = abc_11867_new_n1719
* NET  1196 = abc_11867_new_n1718
* NET  1197 = abc_11867_new_n1717
* NET  1198 = abc_11867_new_n1716
* NET  1199 = abc_11867_new_n1715
* NET  1200 = abc_11867_new_n1714
* NET  1201 = abc_11867_new_n1713
* NET  1202 = abc_11867_new_n1712
* NET  1203 = abc_11867_new_n1711
* NET  1204 = abc_11867_new_n1710
* NET  1205 = abc_11867_new_n1708
* NET  1206 = abc_11867_new_n1707
* NET  1207 = abc_11867_new_n1706
* NET  1208 = abc_11867_new_n1705
* NET  1209 = abc_11867_new_n1704
* NET  1210 = abc_11867_new_n1703
* NET  1211 = abc_11867_new_n1702
* NET  1212 = abc_11867_new_n1701
* NET  1213 = abc_11867_new_n1700
* NET  1214 = abc_11867_new_n1699
* NET  1215 = abc_11867_new_n1698
* NET  1216 = abc_11867_new_n1697
* NET  1217 = abc_11867_new_n1696
* NET  1218 = abc_11867_new_n1694
* NET  1219 = abc_11867_new_n1693
* NET  1220 = abc_11867_new_n1692
* NET  1221 = abc_11867_new_n1691
* NET  1222 = abc_11867_new_n1690
* NET  1223 = abc_11867_new_n1689
* NET  1224 = abc_11867_new_n1688
* NET  1225 = abc_11867_new_n1687
* NET  1226 = abc_11867_new_n1686
* NET  1227 = abc_11867_new_n1685
* NET  1228 = abc_11867_new_n1684
* NET  1229 = abc_11867_new_n1683
* NET  1230 = abc_11867_new_n1682
* NET  1231 = abc_11867_new_n1680
* NET  1232 = abc_11867_new_n1679
* NET  1233 = abc_11867_new_n1678
* NET  1234 = abc_11867_new_n1677
* NET  1235 = abc_11867_new_n1676
* NET  1236 = abc_11867_new_n1675
* NET  1237 = abc_11867_new_n1674
* NET  1238 = abc_11867_new_n1673
* NET  1239 = abc_11867_new_n1672
* NET  1240 = abc_11867_new_n1671
* NET  1241 = abc_11867_new_n1670
* NET  1242 = abc_11867_new_n1669
* NET  1243 = abc_11867_new_n1667
* NET  1244 = abc_11867_new_n1666
* NET  1245 = abc_11867_new_n1665
* NET  1246 = abc_11867_new_n1664
* NET  1247 = abc_11867_new_n1663
* NET  1248 = abc_11867_new_n1662
* NET  1249 = abc_11867_new_n1661
* NET  1250 = abc_11867_new_n1660
* NET  1251 = abc_11867_new_n1659
* NET  1252 = abc_11867_new_n1658
* NET  1253 = abc_11867_new_n1657
* NET  1254 = abc_11867_new_n1655
* NET  1255 = abc_11867_new_n1654
* NET  1256 = abc_11867_new_n1653
* NET  1257 = abc_11867_new_n1652
* NET  1258 = abc_11867_new_n1651
* NET  1259 = abc_11867_new_n1650
* NET  1260 = abc_11867_new_n1649
* NET  1261 = abc_11867_new_n1648
* NET  1262 = abc_11867_new_n1647
* NET  1263 = abc_11867_new_n1645
* NET  1264 = abc_11867_new_n1644
* NET  1265 = abc_11867_new_n1643
* NET  1266 = abc_11867_new_n1642
* NET  1267 = abc_11867_new_n1641
* NET  1268 = abc_11867_new_n1640
* NET  1269 = abc_11867_new_n1639
* NET  1270 = abc_11867_new_n1638
* NET  1271 = abc_11867_new_n1637
* NET  1272 = abc_11867_new_n1635
* NET  1273 = abc_11867_new_n1634
* NET  1274 = abc_11867_new_n1633
* NET  1275 = abc_11867_new_n1632
* NET  1276 = abc_11867_new_n1631
* NET  1277 = abc_11867_new_n1630
* NET  1278 = abc_11867_new_n1629
* NET  1279 = abc_11867_new_n1628
* NET  1280 = abc_11867_new_n1627
* NET  1281 = abc_11867_new_n1626
* NET  1282 = abc_11867_new_n1624
* NET  1283 = abc_11867_new_n1623
* NET  1284 = abc_11867_new_n1622
* NET  1285 = abc_11867_new_n1621
* NET  1286 = abc_11867_new_n1620
* NET  1287 = abc_11867_new_n1619
* NET  1288 = abc_11867_new_n1618
* NET  1289 = abc_11867_new_n1617
* NET  1290 = abc_11867_new_n1616
* NET  1291 = abc_11867_new_n1614
* NET  1292 = abc_11867_new_n1613
* NET  1293 = abc_11867_new_n1612
* NET  1294 = abc_11867_new_n1611
* NET  1295 = abc_11867_new_n1610
* NET  1296 = abc_11867_new_n1609
* NET  1297 = abc_11867_new_n1608
* NET  1298 = abc_11867_new_n1607
* NET  1299 = abc_11867_new_n1606
* NET  1300 = abc_11867_new_n1605
* NET  1301 = abc_11867_new_n1603
* NET  1302 = abc_11867_new_n1602
* NET  1303 = abc_11867_new_n1601
* NET  1304 = abc_11867_new_n1600
* NET  1305 = abc_11867_new_n1599
* NET  1306 = abc_11867_new_n1598
* NET  1307 = abc_11867_new_n1597
* NET  1308 = abc_11867_new_n1596
* NET  1309 = abc_11867_new_n1595
* NET  1310 = abc_11867_new_n1593
* NET  1311 = abc_11867_new_n1592
* NET  1312 = abc_11867_new_n1591
* NET  1313 = abc_11867_new_n1590
* NET  1314 = abc_11867_new_n1589
* NET  1315 = abc_11867_new_n1588
* NET  1316 = abc_11867_new_n1587
* NET  1317 = abc_11867_new_n1586
* NET  1318 = abc_11867_new_n1585
* NET  1319 = abc_11867_new_n1584
* NET  1320 = abc_11867_new_n1583
* NET  1321 = abc_11867_new_n1582
* NET  1322 = abc_11867_new_n1581
* NET  1323 = abc_11867_new_n1580
* NET  1324 = abc_11867_new_n1579
* NET  1325 = abc_11867_new_n1578
* NET  1326 = abc_11867_new_n1577
* NET  1327 = abc_11867_new_n1576
* NET  1328 = abc_11867_new_n1575
* NET  1329 = abc_11867_new_n1574
* NET  1330 = abc_11867_new_n1573
* NET  1331 = abc_11867_new_n1572
* NET  1332 = abc_11867_new_n1571
* NET  1333 = abc_11867_new_n1570
* NET  1334 = abc_11867_new_n1553
* NET  1335 = abc_11867_new_n1552
* NET  1336 = abc_11867_new_n1551
* NET  1337 = abc_11867_new_n1550
* NET  1338 = abc_11867_new_n1549
* NET  1339 = abc_11867_new_n1548
* NET  1340 = abc_11867_new_n1547
* NET  1341 = abc_11867_new_n1546
* NET  1342 = abc_11867_new_n1545
* NET  1343 = abc_11867_new_n1544
* NET  1344 = abc_11867_new_n1543
* NET  1345 = abc_11867_new_n1542
* NET  1346 = abc_11867_new_n1541
* NET  1347 = abc_11867_new_n1540
* NET  1348 = abc_11867_new_n1539
* NET  1349 = abc_11867_new_n1538
* NET  1350 = abc_11867_new_n1537
* NET  1351 = abc_11867_new_n1536
* NET  1352 = abc_11867_new_n1535
* NET  1353 = abc_11867_new_n1534
* NET  1354 = abc_11867_new_n1533
* NET  1355 = abc_11867_new_n1532
* NET  1356 = abc_11867_new_n1531
* NET  1357 = abc_11867_new_n1530
* NET  1358 = abc_11867_new_n1529
* NET  1359 = abc_11867_new_n1528
* NET  1360 = abc_11867_new_n1527
* NET  1361 = abc_11867_new_n1526
* NET  1362 = abc_11867_new_n1525
* NET  1363 = abc_11867_new_n1524
* NET  1364 = abc_11867_new_n1523
* NET  1365 = abc_11867_new_n1522
* NET  1366 = abc_11867_new_n1521
* NET  1367 = abc_11867_new_n1520
* NET  1368 = abc_11867_new_n1519
* NET  1369 = abc_11867_new_n1518
* NET  1370 = abc_11867_new_n1517
* NET  1371 = abc_11867_new_n1516
* NET  1372 = abc_11867_new_n1515
* NET  1373 = abc_11867_new_n1514
* NET  1374 = abc_11867_new_n1513
* NET  1375 = abc_11867_new_n1512
* NET  1376 = abc_11867_new_n1511
* NET  1377 = abc_11867_new_n1510
* NET  1378 = abc_11867_new_n1509
* NET  1379 = abc_11867_new_n1508
* NET  1380 = abc_11867_new_n1507
* NET  1381 = abc_11867_new_n1504
* NET  1382 = abc_11867_new_n1503
* NET  1383 = abc_11867_new_n1502
* NET  1384 = abc_11867_new_n1501
* NET  1385 = abc_11867_new_n1500
* NET  1386 = abc_11867_new_n1499
* NET  1387 = abc_11867_new_n1498
* NET  1388 = abc_11867_new_n1497
* NET  1389 = abc_11867_new_n1496
* NET  1390 = abc_11867_new_n1495
* NET  1391 = abc_11867_new_n1494
* NET  1392 = abc_11867_new_n1493
* NET  1393 = abc_11867_new_n1492
* NET  1394 = abc_11867_new_n1491
* NET  1395 = abc_11867_new_n1489
* NET  1396 = abc_11867_new_n1488
* NET  1397 = abc_11867_new_n1487
* NET  1398 = abc_11867_new_n1486
* NET  1399 = abc_11867_new_n1485
* NET  1400 = abc_11867_new_n1484
* NET  1401 = abc_11867_new_n1483
* NET  1402 = abc_11867_new_n1482
* NET  1403 = abc_11867_new_n1481
* NET  1404 = abc_11867_new_n1479
* NET  1405 = abc_11867_new_n1478
* NET  1406 = abc_11867_new_n1477
* NET  1407 = abc_11867_new_n1476
* NET  1408 = abc_11867_new_n1475
* NET  1409 = abc_11867_new_n1474
* NET  1410 = abc_11867_new_n1473
* NET  1411 = abc_11867_new_n1471
* NET  1412 = abc_11867_new_n1470
* NET  1413 = abc_11867_new_n1469
* NET  1414 = abc_11867_new_n1468
* NET  1415 = abc_11867_new_n1467
* NET  1416 = abc_11867_new_n1465
* NET  1417 = abc_11867_new_n1464
* NET  1418 = abc_11867_new_n1463
* NET  1419 = abc_11867_new_n1462
* NET  1420 = abc_11867_new_n1461
* NET  1421 = abc_11867_new_n1460
* NET  1422 = abc_11867_new_n1459
* NET  1423 = abc_11867_new_n1458
* NET  1424 = abc_11867_new_n1457
* NET  1425 = abc_11867_new_n1455
* NET  1426 = abc_11867_new_n1454
* NET  1427 = abc_11867_new_n1453
* NET  1428 = abc_11867_new_n1452
* NET  1429 = abc_11867_new_n1451
* NET  1430 = abc_11867_new_n1450
* NET  1431 = abc_11867_new_n1449
* NET  1432 = abc_11867_new_n1448
* NET  1433 = abc_11867_new_n1447
* NET  1434 = abc_11867_new_n1446
* NET  1435 = abc_11867_new_n1445
* NET  1436 = abc_11867_new_n1444
* NET  1437 = abc_11867_new_n1443
* NET  1438 = abc_11867_new_n1434
* NET  1439 = abc_11867_new_n1432
* NET  1440 = abc_11867_new_n1431
* NET  1441 = abc_11867_new_n1430
* NET  1442 = abc_11867_new_n1429
* NET  1443 = abc_11867_new_n1428
* NET  1444 = abc_11867_new_n1426
* NET  1445 = abc_11867_new_n1425
* NET  1446 = abc_11867_new_n1424
* NET  1447 = abc_11867_new_n1423
* NET  1448 = abc_11867_new_n1422
* NET  1449 = abc_11867_new_n1421
* NET  1450 = abc_11867_new_n1420
* NET  1451 = abc_11867_new_n1419
* NET  1452 = abc_11867_new_n1418
* NET  1453 = abc_11867_new_n1417
* NET  1454 = abc_11867_new_n1416
* NET  1455 = abc_11867_new_n1415
* NET  1456 = abc_11867_new_n1414
* NET  1457 = abc_11867_new_n1413
* NET  1458 = abc_11867_new_n1410
* NET  1459 = abc_11867_new_n1409
* NET  1460 = abc_11867_new_n1408
* NET  1461 = abc_11867_new_n1407
* NET  1462 = abc_11867_new_n1406
* NET  1463 = abc_11867_new_n1404
* NET  1464 = abc_11867_new_n1403
* NET  1465 = abc_11867_new_n1402
* NET  1466 = abc_11867_new_n1401
* NET  1467 = abc_11867_new_n1400
* NET  1468 = abc_11867_new_n1399
* NET  1469 = abc_11867_new_n1397
* NET  1470 = abc_11867_new_n1396
* NET  1471 = abc_11867_new_n1395
* NET  1472 = abc_11867_new_n1394
* NET  1473 = abc_11867_new_n1393
* NET  1474 = abc_11867_new_n1392
* NET  1475 = abc_11867_new_n1391
* NET  1476 = abc_11867_new_n1390
* NET  1477 = abc_11867_new_n1389
* NET  1478 = abc_11867_new_n1387
* NET  1479 = abc_11867_new_n1386
* NET  1480 = abc_11867_new_n1385
* NET  1481 = abc_11867_new_n1384
* NET  1482 = abc_11867_new_n1383
* NET  1483 = abc_11867_new_n1382
* NET  1484 = abc_11867_new_n1381
* NET  1485 = abc_11867_new_n1380
* NET  1486 = abc_11867_new_n1378
* NET  1487 = abc_11867_new_n1377
* NET  1488 = abc_11867_new_n1376
* NET  1489 = abc_11867_new_n1374
* NET  1490 = abc_11867_new_n1373
* NET  1491 = abc_11867_new_n1372
* NET  1492 = abc_11867_new_n1371
* NET  1493 = abc_11867_new_n1369
* NET  1494 = abc_11867_new_n1368
* NET  1495 = abc_11867_new_n1366
* NET  1496 = abc_11867_new_n1365
* NET  1497 = abc_11867_new_n1363
* NET  1498 = abc_11867_new_n1362
* NET  1499 = abc_11867_new_n1361
* NET  1500 = abc_11867_new_n1358
* NET  1501 = abc_11867_new_n1357
* NET  1502 = abc_11867_new_n1356
* NET  1503 = abc_11867_new_n1355
* NET  1504 = abc_11867_new_n1353
* NET  1505 = abc_11867_new_n1352
* NET  1506 = abc_11867_new_n1351
* NET  1507 = abc_11867_new_n1350
* NET  1508 = abc_11867_new_n1349
* NET  1509 = abc_11867_new_n1348
* NET  1510 = abc_11867_new_n1347
* NET  1511 = abc_11867_new_n1345
* NET  1512 = abc_11867_new_n1344
* NET  1513 = abc_11867_new_n1341
* NET  1514 = abc_11867_new_n1340
* NET  1515 = abc_11867_new_n1339
* NET  1516 = abc_11867_new_n1338
* NET  1517 = abc_11867_new_n1337
* NET  1518 = abc_11867_new_n1334
* NET  1519 = abc_11867_new_n1333
* NET  1520 = abc_11867_new_n1332
* NET  1521 = abc_11867_new_n1331
* NET  1522 = abc_11867_new_n1330
* NET  1523 = abc_11867_new_n1329
* NET  1524 = abc_11867_new_n1328
* NET  1525 = abc_11867_new_n1327
* NET  1526 = abc_11867_new_n1326
* NET  1527 = abc_11867_new_n1325
* NET  1528 = abc_11867_new_n1324
* NET  1529 = abc_11867_new_n1323
* NET  1530 = abc_11867_new_n1322
* NET  1531 = abc_11867_new_n1321
* NET  1532 = abc_11867_new_n1320
* NET  1533 = abc_11867_new_n1319
* NET  1534 = abc_11867_new_n1317
* NET  1535 = abc_11867_new_n1316
* NET  1536 = abc_11867_new_n1315
* NET  1537 = abc_11867_new_n1314
* NET  1538 = abc_11867_new_n1313
* NET  1539 = abc_11867_new_n1311
* NET  1540 = abc_11867_new_n1310
* NET  1541 = abc_11867_new_n1309
* NET  1542 = abc_11867_new_n1308
* NET  1543 = abc_11867_new_n1307
* NET  1544 = abc_11867_new_n1306
* NET  1545 = abc_11867_new_n1305
* NET  1546 = abc_11867_new_n1304
* NET  1547 = abc_11867_new_n1303
* NET  1548 = abc_11867_new_n1302
* NET  1549 = abc_11867_new_n1301
* NET  1550 = abc_11867_new_n1299
* NET  1551 = abc_11867_new_n1298
* NET  1552 = abc_11867_new_n1297
* NET  1553 = abc_11867_new_n1295
* NET  1554 = abc_11867_new_n1294
* NET  1555 = abc_11867_new_n1293
* NET  1556 = abc_11867_new_n1292
* NET  1557 = abc_11867_new_n1290
* NET  1558 = abc_11867_new_n1289
* NET  1559 = abc_11867_new_n1287
* NET  1560 = abc_11867_new_n1286
* NET  1561 = abc_11867_new_n1284
* NET  1562 = abc_11867_new_n1282
* NET  1563 = abc_11867_new_n1281
* NET  1564 = abc_11867_new_n1280
* NET  1565 = abc_11867_new_n1278
* NET  1566 = abc_11867_new_n1277
* NET  1567 = abc_11867_new_n1276
* NET  1568 = abc_11867_new_n1275
* NET  1569 = abc_11867_new_n1273
* NET  1570 = abc_11867_new_n1272
* NET  1571 = abc_11867_new_n1271
* NET  1572 = abc_11867_new_n1269
* NET  1573 = abc_11867_new_n1267
* NET  1574 = abc_11867_new_n1266
* NET  1575 = abc_11867_new_n1265
* NET  1576 = abc_11867_new_n1264
* NET  1577 = abc_11867_new_n1259
* NET  1578 = abc_11867_new_n1250
* NET  1579 = abc_11867_new_n1241
* NET  1580 = abc_11867_new_n1232
* NET  1581 = abc_11867_new_n1230
* NET  1582 = abc_11867_new_n1229
* NET  1583 = abc_11867_new_n1228
* NET  1584 = abc_11867_new_n1227
* NET  1585 = abc_11867_new_n1226
* NET  1586 = abc_11867_new_n1224
* NET  1587 = abc_11867_new_n1223
* NET  1588 = abc_11867_new_n1222
* NET  1589 = abc_11867_new_n1221
* NET  1590 = abc_11867_new_n1220
* NET  1591 = abc_11867_new_n1219
* NET  1592 = abc_11867_new_n1218
* NET  1593 = abc_11867_new_n1216
* NET  1594 = abc_11867_new_n1215
* NET  1595 = abc_11867_new_n1214
* NET  1596 = abc_11867_new_n1213
* NET  1597 = abc_11867_new_n1212
* NET  1598 = abc_11867_new_n1211
* NET  1599 = abc_11867_new_n1209
* NET  1600 = abc_11867_new_n1207
* NET  1601 = abc_11867_new_n1206
* NET  1602 = abc_11867_new_n1205
* NET  1603 = abc_11867_new_n1204
* NET  1604 = abc_11867_new_n1203
* NET  1605 = abc_11867_new_n1201
* NET  1606 = abc_11867_new_n1200
* NET  1607 = abc_11867_new_n1199
* NET  1608 = abc_11867_new_n1198
* NET  1609 = abc_11867_new_n1197
* NET  1610 = abc_11867_new_n1196
* NET  1611 = abc_11867_new_n1195
* NET  1612 = abc_11867_new_n1193
* NET  1613 = abc_11867_new_n1192
* NET  1614 = abc_11867_new_n1191
* NET  1615 = abc_11867_new_n1190
* NET  1616 = abc_11867_new_n1189
* NET  1617 = abc_11867_new_n1188
* NET  1618 = abc_11867_new_n1186
* NET  1619 = abc_11867_new_n1185
* NET  1620 = abc_11867_new_n1184
* NET  1621 = abc_11867_new_n1183
* NET  1622 = abc_11867_new_n1182
* NET  1623 = abc_11867_new_n1181
* NET  1624 = abc_11867_new_n1180
* NET  1625 = abc_11867_new_n1179
* NET  1626 = abc_11867_new_n1176
* NET  1627 = abc_11867_new_n1175
* NET  1628 = abc_11867_new_n1174
* NET  1629 = abc_11867_new_n1173
* NET  1630 = abc_11867_new_n1172
* NET  1631 = abc_11867_new_n1171
* NET  1632 = abc_11867_new_n1170
* NET  1633 = abc_11867_new_n1168
* NET  1634 = abc_11867_new_n1167
* NET  1635 = abc_11867_new_n1166
* NET  1636 = abc_11867_new_n1165
* NET  1637 = abc_11867_new_n1164
* NET  1638 = abc_11867_new_n1163
* NET  1639 = abc_11867_new_n1162
* NET  1640 = abc_11867_new_n1160
* NET  1641 = abc_11867_new_n1159
* NET  1642 = abc_11867_new_n1158
* NET  1643 = abc_11867_new_n1157
* NET  1644 = abc_11867_new_n1156
* NET  1645 = abc_11867_new_n1155
* NET  1646 = abc_11867_new_n1154
* NET  1647 = abc_11867_new_n1152
* NET  1648 = abc_11867_new_n1151
* NET  1649 = abc_11867_new_n1150
* NET  1650 = abc_11867_new_n1149
* NET  1651 = abc_11867_new_n1148
* NET  1652 = abc_11867_new_n1147
* NET  1653 = abc_11867_new_n1146
* NET  1654 = abc_11867_new_n1144
* NET  1655 = abc_11867_new_n1143
* NET  1656 = abc_11867_new_n1142
* NET  1657 = abc_11867_new_n1141
* NET  1658 = abc_11867_new_n1140
* NET  1659 = abc_11867_new_n1139
* NET  1660 = abc_11867_new_n1138
* NET  1661 = abc_11867_new_n1136
* NET  1662 = abc_11867_new_n1135
* NET  1663 = abc_11867_new_n1134
* NET  1664 = abc_11867_new_n1133
* NET  1665 = abc_11867_new_n1132
* NET  1666 = abc_11867_new_n1131
* NET  1667 = abc_11867_new_n1130
* NET  1668 = abc_11867_new_n1128
* NET  1669 = abc_11867_new_n1127
* NET  1670 = abc_11867_new_n1126
* NET  1671 = abc_11867_new_n1125
* NET  1672 = abc_11867_new_n1124
* NET  1673 = abc_11867_new_n1123
* NET  1674 = abc_11867_new_n1122
* NET  1675 = abc_11867_new_n1120
* NET  1676 = abc_11867_new_n1119
* NET  1677 = abc_11867_new_n1118
* NET  1678 = abc_11867_new_n1117
* NET  1679 = abc_11867_new_n1116
* NET  1680 = abc_11867_new_n1115
* NET  1681 = abc_11867_new_n1114
* NET  1682 = abc_11867_new_n1113
* NET  1683 = abc_11867_new_n1112
* NET  1684 = abc_11867_new_n1110
* NET  1685 = abc_11867_new_n1109
* NET  1686 = abc_11867_new_n1108
* NET  1687 = abc_11867_new_n1107
* NET  1688 = abc_11867_new_n1106
* NET  1689 = abc_11867_new_n1105
* NET  1690 = abc_11867_new_n1104
* NET  1691 = abc_11867_new_n1102
* NET  1692 = abc_11867_new_n1101
* NET  1693 = abc_11867_new_n1100
* NET  1694 = abc_11867_new_n1099
* NET  1695 = abc_11867_new_n1098
* NET  1696 = abc_11867_new_n1097
* NET  1697 = abc_11867_new_n1096
* NET  1698 = abc_11867_new_n1094
* NET  1699 = abc_11867_new_n1093
* NET  1700 = abc_11867_new_n1092
* NET  1701 = abc_11867_new_n1091
* NET  1702 = abc_11867_new_n1090
* NET  1703 = abc_11867_new_n1089
* NET  1704 = abc_11867_new_n1088
* NET  1705 = abc_11867_new_n1086
* NET  1706 = abc_11867_new_n1085
* NET  1707 = abc_11867_new_n1084
* NET  1708 = abc_11867_new_n1083
* NET  1709 = abc_11867_new_n1082
* NET  1710 = abc_11867_new_n1081
* NET  1711 = abc_11867_new_n1080
* NET  1712 = abc_11867_new_n1078
* NET  1713 = abc_11867_new_n1077
* NET  1714 = abc_11867_new_n1076
* NET  1715 = abc_11867_new_n1075
* NET  1716 = abc_11867_new_n1074
* NET  1717 = abc_11867_new_n1073
* NET  1718 = abc_11867_new_n1072
* NET  1719 = abc_11867_new_n1070
* NET  1720 = abc_11867_new_n1069
* NET  1721 = abc_11867_new_n1068
* NET  1722 = abc_11867_new_n1067
* NET  1723 = abc_11867_new_n1066
* NET  1724 = abc_11867_new_n1065
* NET  1725 = abc_11867_new_n1064
* NET  1726 = abc_11867_new_n1062
* NET  1727 = abc_11867_new_n1061
* NET  1728 = abc_11867_new_n1060
* NET  1729 = abc_11867_new_n1059
* NET  1730 = abc_11867_new_n1058
* NET  1731 = abc_11867_new_n1057
* NET  1732 = abc_11867_new_n1056
* NET  1733 = abc_11867_new_n1054
* NET  1734 = abc_11867_new_n1053
* NET  1735 = abc_11867_new_n1052
* NET  1736 = abc_11867_new_n1051
* NET  1737 = abc_11867_new_n1050
* NET  1738 = abc_11867_new_n1049
* NET  1739 = abc_11867_new_n1048
* NET  1740 = abc_11867_new_n1047
* NET  1741 = abc_11867_new_n1046
* NET  1742 = abc_11867_new_n1045
* NET  1743 = abc_11867_new_n1044
* NET  1744 = abc_11867_new_n1043
* NET  1745 = abc_11867_new_n1042
* NET  1746 = abc_11867_new_n1041
* NET  1747 = abc_11867_new_n1040
* NET  1748 = abc_11867_new_n1039
* NET  1749 = abc_11867_new_n1038
* NET  1750 = abc_11867_new_n1037
* NET  1751 = abc_11867_new_n1036
* NET  1752 = abc_11867_new_n1035
* NET  1753 = abc_11867_new_n1034
* NET  1754 = abc_11867_new_n1033
* NET  1755 = abc_11867_new_n1032
* NET  1756 = abc_11867_new_n1031
* NET  1757 = abc_11867_new_n1030
* NET  1758 = abc_11867_new_n1029
* NET  1759 = abc_11867_new_n1028
* NET  1760 = abc_11867_new_n1027
* NET  1761 = abc_11867_new_n1026
* NET  1762 = abc_11867_new_n1025
* NET  1763 = abc_11867_new_n1024
* NET  1764 = abc_11867_new_n1023
* NET  1765 = abc_11867_new_n1022
* NET  1766 = abc_11867_new_n1021
* NET  1767 = abc_11867_new_n1020
* NET  1768 = abc_11867_new_n1019
* NET  1769 = abc_11867_new_n1018
* NET  1770 = abc_11867_new_n1016
* NET  1771 = abc_11867_new_n1015
* NET  1772 = abc_11867_new_n1014
* NET  1773 = abc_11867_new_n1013
* NET  1774 = abc_11867_new_n1012
* NET  1775 = abc_11867_new_n1011
* NET  1776 = abc_11867_new_n1010
* NET  1777 = abc_11867_new_n1009
* NET  1778 = abc_11867_new_n1008
* NET  1779 = abc_11867_new_n1007
* NET  1780 = abc_11867_new_n1006
* NET  1781 = abc_11867_new_n1005
* NET  1782 = abc_11867_new_n1004
* NET  1783 = abc_11867_new_n1003
* NET  1784 = abc_11867_new_n1002
* NET  1785 = abc_11867_new_n1000
* NET  1786 = abc_11867_flatten_MOS6502_0_adj_bcd_0_0
* NET  1787 = abc_11867_auto_rtlil_cc_2608_MuxGate_11866
* NET  1788 = abc_11867_auto_rtlil_cc_2608_MuxGate_11864
* NET  1789 = abc_11867_auto_rtlil_cc_2608_MuxGate_11862
* NET  1790 = abc_11867_auto_rtlil_cc_2608_MuxGate_11860
* NET  1791 = abc_11867_auto_rtlil_cc_2608_MuxGate_11858
* NET  1792 = abc_11867_auto_rtlil_cc_2608_MuxGate_11856
* NET  1793 = abc_11867_auto_rtlil_cc_2608_MuxGate_11854
* NET  1794 = abc_11867_auto_rtlil_cc_2608_MuxGate_11852
* NET  1795 = abc_11867_auto_rtlil_cc_2608_MuxGate_11850
* NET  1796 = abc_11867_auto_rtlil_cc_2608_MuxGate_11848
* NET  1797 = abc_11867_auto_rtlil_cc_2608_MuxGate_11846
* NET  1798 = abc_11867_auto_rtlil_cc_2608_MuxGate_11844
* NET  1799 = abc_11867_auto_rtlil_cc_2608_MuxGate_11842
* NET  1800 = abc_11867_auto_rtlil_cc_2608_MuxGate_11840
* NET  1801 = abc_11867_auto_rtlil_cc_2608_MuxGate_11838
* NET  1802 = abc_11867_auto_rtlil_cc_2608_MuxGate_11836
* NET  1803 = abc_11867_auto_rtlil_cc_2608_MuxGate_11834
* NET  1804 = abc_11867_auto_rtlil_cc_2608_MuxGate_11832
* NET  1805 = abc_11867_auto_rtlil_cc_2608_MuxGate_11830
* NET  1806 = abc_11867_auto_rtlil_cc_2608_MuxGate_11828
* NET  1807 = abc_11867_auto_rtlil_cc_2608_MuxGate_11826
* NET  1808 = abc_11867_auto_rtlil_cc_2608_MuxGate_11824
* NET  1809 = abc_11867_auto_rtlil_cc_2608_MuxGate_11822
* NET  1810 = abc_11867_auto_rtlil_cc_2608_MuxGate_11820
* NET  1811 = abc_11867_auto_rtlil_cc_2608_MuxGate_11818
* NET  1812 = abc_11867_auto_rtlil_cc_2608_MuxGate_11816
* NET  1813 = abc_11867_auto_rtlil_cc_2608_MuxGate_11814
* NET  1814 = abc_11867_auto_rtlil_cc_2608_MuxGate_11812
* NET  1815 = abc_11867_auto_rtlil_cc_2608_MuxGate_11810
* NET  1816 = abc_11867_auto_rtlil_cc_2608_MuxGate_11808
* NET  1817 = abc_11867_auto_rtlil_cc_2608_MuxGate_11806
* NET  1818 = abc_11867_auto_rtlil_cc_2608_MuxGate_11804
* NET  1819 = abc_11867_auto_rtlil_cc_2608_MuxGate_11802
* NET  1820 = abc_11867_auto_rtlil_cc_2608_MuxGate_11800
* NET  1821 = abc_11867_auto_rtlil_cc_2608_MuxGate_11798
* NET  1822 = abc_11867_auto_rtlil_cc_2608_MuxGate_11796
* NET  1823 = abc_11867_auto_rtlil_cc_2608_MuxGate_11794
* NET  1824 = abc_11867_auto_rtlil_cc_2608_MuxGate_11792
* NET  1825 = abc_11867_auto_rtlil_cc_2608_MuxGate_11790
* NET  1826 = abc_11867_auto_rtlil_cc_2608_MuxGate_11788
* NET  1827 = abc_11867_auto_rtlil_cc_2608_MuxGate_11786
* NET  1828 = abc_11867_auto_rtlil_cc_2608_MuxGate_11784
* NET  1829 = abc_11867_auto_rtlil_cc_2608_MuxGate_11782
* NET  1830 = abc_11867_auto_rtlil_cc_2608_MuxGate_11780
* NET  1831 = abc_11867_auto_rtlil_cc_2608_MuxGate_11778
* NET  1832 = abc_11867_auto_rtlil_cc_2608_MuxGate_11776
* NET  1833 = abc_11867_auto_rtlil_cc_2608_MuxGate_11774
* NET  1834 = abc_11867_auto_rtlil_cc_2608_MuxGate_11772
* NET  1835 = abc_11867_auto_rtlil_cc_2608_MuxGate_11770
* NET  1836 = abc_11867_auto_rtlil_cc_2608_MuxGate_11768
* NET  1837 = abc_11867_auto_rtlil_cc_2608_MuxGate_11764
* NET  1838 = abc_11867_auto_rtlil_cc_2608_MuxGate_11762
* NET  1839 = abc_11867_auto_rtlil_cc_2608_MuxGate_11760
* NET  1840 = abc_11867_auto_rtlil_cc_2608_MuxGate_11758
* NET  1841 = abc_11867_auto_rtlil_cc_2608_MuxGate_11756
* NET  1842 = abc_11867_auto_rtlil_cc_2608_MuxGate_11754
* NET  1843 = abc_11867_auto_rtlil_cc_2608_MuxGate_11752
* NET  1844 = abc_11867_auto_rtlil_cc_2608_MuxGate_11750
* NET  1845 = abc_11867_auto_rtlil_cc_2608_MuxGate_11748
* NET  1846 = abc_11867_auto_rtlil_cc_2608_MuxGate_11746
* NET  1847 = abc_11867_auto_rtlil_cc_2608_MuxGate_11742
* NET  1848 = abc_11867_auto_rtlil_cc_2608_MuxGate_11740
* NET  1849 = abc_11867_auto_rtlil_cc_2608_MuxGate_11736
* NET  1850 = abc_11867_auto_rtlil_cc_2608_MuxGate_11734
* NET  1851 = abc_11867_auto_rtlil_cc_2608_MuxGate_11732
* NET  1852 = abc_11867_auto_rtlil_cc_2608_MuxGate_11730
* NET  1853 = abc_11867_auto_rtlil_cc_2608_MuxGate_11728
* NET  1854 = abc_11867_auto_rtlil_cc_2608_MuxGate_11726
* NET  1855 = abc_11867_auto_rtlil_cc_2608_MuxGate_11724
* NET  1856 = abc_11867_auto_rtlil_cc_2608_MuxGate_11722
* NET  1857 = abc_11867_auto_rtlil_cc_2608_MuxGate_11720
* NET  1858 = abc_11867_auto_rtlil_cc_2608_MuxGate_11718
* NET  1859 = abc_11867_auto_rtlil_cc_2608_MuxGate_11716
* NET  1860 = abc_11867_auto_rtlil_cc_2608_MuxGate_11714
* NET  1861 = abc_11867_auto_rtlil_cc_2608_MuxGate_11710
* NET  1862 = abc_11867_auto_rtlil_cc_2608_MuxGate_11708
* NET  1863 = abc_11867_auto_rtlil_cc_2608_MuxGate_11706
* NET  1864 = abc_11867_auto_rtlil_cc_2608_MuxGate_11704
* NET  1865 = abc_11867_auto_rtlil_cc_2608_MuxGate_11702
* NET  1866 = abc_11867_auto_rtlil_cc_2608_MuxGate_11700
* NET  1867 = abc_11867_auto_rtlil_cc_2608_MuxGate_11698
* NET  1868 = abc_11867_auto_rtlil_cc_2608_MuxGate_11696
* NET  1869 = abc_11867_auto_rtlil_cc_2608_MuxGate_11694
* NET  1870 = abc_11867_auto_rtlil_cc_2608_MuxGate_11692
* NET  1871 = abc_11867_auto_rtlil_cc_2608_MuxGate_11690
* NET  1872 = abc_11867_auto_rtlil_cc_2608_MuxGate_11688
* NET  1873 = abc_11867_auto_rtlil_cc_2608_MuxGate_11686
* NET  1874 = abc_11867_auto_rtlil_cc_2608_MuxGate_11684
* NET  1875 = abc_11867_auto_rtlil_cc_2608_MuxGate_11682
* NET  1876 = abc_11867_auto_rtlil_cc_2608_MuxGate_11680
* NET  1877 = abc_11867_auto_rtlil_cc_2608_MuxGate_11678
* NET  1878 = abc_11867_auto_rtlil_cc_2608_MuxGate_11676
* NET  1879 = abc_11867_auto_rtlil_cc_2608_MuxGate_11674
* NET  1880 = abc_11867_auto_rtlil_cc_2608_MuxGate_11672
* NET  1881 = abc_11867_auto_rtlil_cc_2608_MuxGate_11670
* NET  1882 = abc_11867_auto_rtlil_cc_2608_MuxGate_11666
* NET  1883 = abc_11867_auto_rtlil_cc_2608_MuxGate_11664
* NET  1884 = abc_11867_auto_rtlil_cc_2608_MuxGate_11662
* NET  1885 = abc_11867_auto_rtlil_cc_2608_MuxGate_11660
* NET  1886 = abc_11867_auto_rtlil_cc_2608_MuxGate_11658
* NET  1887 = abc_11867_auto_rtlil_cc_2608_MuxGate_11656
* NET  1888 = abc_11867_auto_rtlil_cc_2608_MuxGate_11654
* NET  1889 = abc_11867_auto_rtlil_cc_2608_MuxGate_11652
* NET  1890 = abc_11867_auto_rtlil_cc_2608_MuxGate_11650
* NET  1891 = abc_11867_auto_rtlil_cc_2608_MuxGate_11648
* NET  1892 = abc_11867_auto_rtlil_cc_2608_MuxGate_11646
* NET  1893 = abc_11867_auto_rtlil_cc_2608_MuxGate_11644
* NET  1894 = abc_11867_auto_rtlil_cc_2608_MuxGate_11642
* NET  1895 = abc_11867_auto_rtlil_cc_2608_MuxGate_11640
* NET  1896 = abc_11867_auto_rtlil_cc_2608_MuxGate_11638
* NET  1897 = abc_11867_auto_rtlil_cc_2608_MuxGate_11636
* NET  1898 = abc_11867_auto_rtlil_cc_2608_MuxGate_11634
* NET  1899 = abc_11867_auto_rtlil_cc_2608_MuxGate_11632
* NET  1900 = abc_11867_auto_rtlil_cc_2608_MuxGate_11630
* NET  1901 = abc_11867_auto_rtlil_cc_2608_MuxGate_11628
* NET  1902 = abc_11867_auto_rtlil_cc_2608_MuxGate_11626
* NET  1903 = abc_11867_auto_rtlil_cc_2608_MuxGate_11624
* NET  1904 = abc_11867_auto_rtlil_cc_2608_MuxGate_11622
* NET  1905 = abc_11867_auto_rtlil_cc_2608_MuxGate_11620
* NET  1906 = abc_11867_auto_rtlil_cc_2608_MuxGate_11618
* NET  1907 = abc_11867_auto_rtlil_cc_2608_MuxGate_11616
* NET  1908 = abc_11867_auto_rtlil_cc_2608_MuxGate_11614
* NET  1909 = abc_11867_auto_rtlil_cc_2608_MuxGate_11612
* NET  1910 = abc_11867_auto_rtlil_cc_2608_MuxGate_11610
* NET  1911 = abc_11867_auto_rtlil_cc_2608_MuxGate_11608
* NET  1912 = abc_11867_auto_rtlil_cc_2608_MuxGate_11606
* NET  1913 = abc_11867_auto_rtlil_cc_2608_MuxGate_11604
* NET  1914 = WE
* NET  1915 = RDY_hfns_2
* NET  1916 = RDY_hfns_1
* NET  1917 = RDY_hfns_0
* NET  1918 = RDY
* NET  1919 = NMI
* NET  1920 = MOS6502_write_back
* NET  1921 = MOS6502_store
* NET  1922 = MOS6502_state_bit0_hfns_2
* NET  1923 = MOS6502_state_bit0_hfns_1
* NET  1924 = MOS6502_state_bit0_hfns_0
* NET  1925 = MOS6502_state[5]
* NET  1926 = MOS6502_state[4]
* NET  1927 = MOS6502_state[3]
* NET  1928 = MOS6502_state[2]
* NET  1929 = MOS6502_state[1]
* NET  1930 = MOS6502_state[0]
* NET  1931 = MOS6502_src_reg[1]
* NET  1932 = MOS6502_src_reg[0]
* NET  1933 = MOS6502_shift_right
* NET  1934 = MOS6502_shift
* NET  1935 = MOS6502_sei
* NET  1936 = MOS6502_sed
* NET  1937 = MOS6502_sec
* NET  1938 = MOS6502_rotate
* NET  1939 = MOS6502_res
* NET  1940 = MOS6502_plp
* NET  1941 = MOS6502_php
* NET  1942 = MOS6502_op[3]
* NET  1943 = MOS6502_op[2]
* NET  1944 = MOS6502_op[1]
* NET  1945 = MOS6502_op[0]
* NET  1946 = MOS6502_load_reg
* NET  1947 = MOS6502_load_only
* NET  1948 = MOS6502_index_y
* NET  1949 = MOS6502_inc
* NET  1950 = MOS6502_dst_reg[1]
* NET  1951 = MOS6502_dst_reg[0]
* NET  1952 = MOS6502_cond_code[2]
* NET  1953 = MOS6502_cond_code[1]
* NET  1954 = MOS6502_cond_code[0]
* NET  1955 = MOS6502_compare
* NET  1956 = MOS6502_clv
* NET  1957 = MOS6502_cli
* NET  1958 = MOS6502_cld
* NET  1959 = MOS6502_clc
* NET  1960 = MOS6502_bit_ins
* NET  1961 = MOS6502_backwards
* NET  1962 = MOS6502_adj_bcd
* NET  1963 = MOS6502_adc_sbc
* NET  1964 = MOS6502_adc_bcd
* NET  1965 = MOS6502_Z
* NET  1966 = MOS6502_V
* NET  1967 = MOS6502_PC[9]
* NET  1968 = MOS6502_PC[8]
* NET  1969 = MOS6502_PC[7]
* NET  1970 = MOS6502_PC[6]
* NET  1971 = MOS6502_PC[5]
* NET  1972 = MOS6502_PC[4]
* NET  1973 = MOS6502_PC[3]
* NET  1974 = MOS6502_PC[2]
* NET  1975 = MOS6502_PC[15]
* NET  1976 = MOS6502_PC[14]
* NET  1977 = MOS6502_PC[13]
* NET  1978 = MOS6502_PC[12]
* NET  1979 = MOS6502_PC[11]
* NET  1980 = MOS6502_PC[10]
* NET  1981 = MOS6502_PC[1]
* NET  1982 = MOS6502_PC[0]
* NET  1983 = MOS6502_NMI_edge
* NET  1984 = MOS6502_NMI_1
* NET  1985 = MOS6502_N
* NET  1986 = MOS6502_IRHOLD_valid
* NET  1987 = MOS6502_IRHOLD[7]
* NET  1988 = MOS6502_IRHOLD[6]
* NET  1989 = MOS6502_IRHOLD[5]
* NET  1990 = MOS6502_IRHOLD[4]
* NET  1991 = MOS6502_IRHOLD[3]
* NET  1992 = MOS6502_IRHOLD[2]
* NET  1993 = MOS6502_IRHOLD[1]
* NET  1994 = MOS6502_IRHOLD[0]
* NET  1995 = MOS6502_I
* NET  1996 = MOS6502_DIMUX[7]
* NET  1997 = MOS6502_DIMUX[6]
* NET  1998 = MOS6502_DIMUX[5]
* NET  1999 = MOS6502_DIMUX[4]
* NET  2000 = MOS6502_DIMUX[3]
* NET  2001 = MOS6502_DIMUX[2]
* NET  2002 = MOS6502_DIMUX[1]
* NET  2003 = MOS6502_DIMUX[0]
* NET  2004 = MOS6502_DIHOLD[7]
* NET  2005 = MOS6502_DIHOLD[6]
* NET  2006 = MOS6502_DIHOLD[5]
* NET  2007 = MOS6502_DIHOLD[4]
* NET  2008 = MOS6502_DIHOLD[3]
* NET  2009 = MOS6502_DIHOLD[2]
* NET  2010 = MOS6502_DIHOLD[1]
* NET  2011 = MOS6502_DIHOLD[0]
* NET  2012 = MOS6502_D
* NET  2013 = MOS6502_C
* NET  2014 = MOS6502_AXYS_3_7
* NET  2015 = MOS6502_AXYS_3_6
* NET  2016 = MOS6502_AXYS_3_5
* NET  2017 = MOS6502_AXYS_3_4
* NET  2018 = MOS6502_AXYS_3_3
* NET  2019 = MOS6502_AXYS_3_2
* NET  2020 = MOS6502_AXYS_3_1
* NET  2021 = MOS6502_AXYS_3_0
* NET  2022 = MOS6502_AXYS_2_7
* NET  2023 = MOS6502_AXYS_2_6
* NET  2024 = MOS6502_AXYS_2_5
* NET  2025 = MOS6502_AXYS_2_4
* NET  2026 = MOS6502_AXYS_2_3
* NET  2027 = MOS6502_AXYS_2_2
* NET  2028 = MOS6502_AXYS_2_1
* NET  2029 = MOS6502_AXYS_2_0
* NET  2030 = MOS6502_AXYS_1_7
* NET  2031 = MOS6502_AXYS_1_6
* NET  2032 = MOS6502_AXYS_1_5
* NET  2033 = MOS6502_AXYS_1_4
* NET  2034 = MOS6502_AXYS_1_3
* NET  2035 = MOS6502_AXYS_1_2
* NET  2036 = MOS6502_AXYS_1_1
* NET  2037 = MOS6502_AXYS_1_0
* NET  2038 = MOS6502_AXYS_0_7
* NET  2039 = MOS6502_AXYS_0_6
* NET  2040 = MOS6502_AXYS_0_5
* NET  2041 = MOS6502_AXYS_0_4
* NET  2042 = MOS6502_AXYS_0_3
* NET  2043 = MOS6502_AXYS_0_2
* NET  2044 = MOS6502_AXYS_0_1
* NET  2045 = MOS6502_AXYS_0_0
* NET  2046 = MOS6502_ALU_OUT[7]
* NET  2047 = MOS6502_ALU_OUT[6]
* NET  2048 = MOS6502_ALU_OUT[5]
* NET  2049 = MOS6502_ALU_OUT[4]
* NET  2050 = MOS6502_ALU_OUT[3]
* NET  2051 = MOS6502_ALU_OUT[2]
* NET  2052 = MOS6502_ALU_OUT[1]
* NET  2053 = MOS6502_ALU_OUT[0]
* NET  2054 = MOS6502_ALU_HC
* NET  2055 = MOS6502_ALU_CO
* NET  2056 = MOS6502_ALU_BI7
* NET  2057 = MOS6502_ALU_AI7
* NET  2058 = MOS6502_ABL[7]
* NET  2059 = MOS6502_ABL[6]
* NET  2060 = MOS6502_ABL[5]
* NET  2061 = MOS6502_ABL[4]
* NET  2062 = MOS6502_ABL[3]
* NET  2063 = MOS6502_ABL[2]
* NET  2064 = MOS6502_ABL[1]
* NET  2065 = MOS6502_ABL[0]
* NET  2066 = MOS6502_ABH[7]
* NET  2067 = MOS6502_ABH[6]
* NET  2068 = MOS6502_ABH[5]
* NET  2069 = MOS6502_ABH[4]
* NET  2070 = MOS6502_ABH[3]
* NET  2071 = MOS6502_ABH[2]
* NET  2072 = MOS6502_ABH[1]
* NET  2073 = MOS6502_ABH[0]
* NET  2074 = IRQ
* NET  2075 = DO[7]
* NET  2076 = DO[6]
* NET  2077 = DO[5]
* NET  2078 = DO[4]
* NET  2079 = DO[3]
* NET  2080 = DO[2]
* NET  2081 = DO[1]
* NET  2082 = DO[0]
* NET  2083 = DI[7]
* NET  2084 = DI[6]
* NET  2085 = DI[5]
* NET  2086 = DI[4]
* NET  2087 = DI[3]
* NET  2088 = DI[2]
* NET  2089 = DI[1]
* NET  2090 = DI[0]
* NET  2091 = A[9]
* NET  2092 = A[8]
* NET  2093 = A[7]
* NET  2094 = A[6]
* NET  2095 = A[5]
* NET  2096 = A[4]
* NET  2097 = A[3]
* NET  2098 = A[2]
* NET  2099 = A[15]
* NET  2100 = A[14]
* NET  2101 = A[13]
* NET  2102 = A[12]
* NET  2103 = A[11]
* NET  2104 = A[10]
* NET  2105 = A[1]
* NET  2106 = A[0]

xfeed_6739 0 1 decap_w0
xfeed_6738 0 1 decap_w0
xfeed_6737 0 1 decap_w0
xfeed_6736 0 1 decap_w0
xfeed_6735 0 1 decap_w0
xfeed_6734 0 1 tie
xfeed_6733 0 1 decap_w0
xfeed_6732 0 1 decap_w0
xfeed_6731 0 1 decap_w0
xfeed_409 0 1 decap_w0
xfeed_408 0 1 decap_w0
xfeed_407 0 1 decap_w0
xfeed_406 0 1 decap_w0
xfeed_405 0 1 decap_w0
xfeed_404 0 1 decap_w0
xfeed_403 0 1 decap_w0
xfeed_402 0 1 decap_w0
xfeed_401 0 1 decap_w0
xfeed_400 0 1 decap_w0
xsubckt_1035_nand2_x0 0 1 1500 1517 1501 nand2_x0
xsubckt_932_mux2_x1 0 1 1885 2025 1599 1578 mux2_x1
xsubckt_1653_and2_x1 0 1 941 944 942 and2_x1
xsubckt_1701_mux2_x1 0 1 893 1103 1105 897 mux2_x1
xspare_buffer_40 0 1 64 68 buf_x4
xspare_buffer_41 0 1 63 68 buf_x4
xspare_buffer_42 0 1 62 68 buf_x4
xspare_buffer_43 0 1 14 16 buf_x4
xspare_buffer_44 0 1 61 68 buf_x4
xfeed_13479 0 1 decap_w0
xfeed_13478 0 1 decap_w0
xfeed_13477 0 1 decap_w0
xfeed_13476 0 1 tie
xfeed_13475 0 1 decap_w0
xfeed_13474 0 1 decap_w0
xfeed_13473 0 1 decap_w0
xfeed_13472 0 1 decap_w0
xfeed_13471 0 1 decap_w0
xfeed_13470 0 1 decap_w0
xfeed_12949 0 1 decap_w0
xfeed_12948 0 1 decap_w0
xfeed_12947 0 1 decap_w0
xfeed_12946 0 1 decap_w0
xfeed_12945 0 1 decap_w0
xfeed_12944 0 1 tie
xfeed_12943 0 1 decap_w0
xfeed_12942 0 1 decap_w0
xfeed_12941 0 1 decap_w0
xfeed_12940 0 1 decap_w0
xfeed_7276 0 1 decap_w0
xfeed_7273 0 1 decap_w0
xfeed_7272 0 1 decap_w0
xfeed_7271 0 1 decap_w0
xfeed_7270 0 1 decap_w0
xfeed_2437 0 1 decap_w0
xfeed_2436 0 1 decap_w0
xfeed_2435 0 1 decap_w0
xfeed_2434 0 1 decap_w0
xfeed_2433 0 1 decap_w0
xfeed_2432 0 1 decap_w0
xfeed_2431 0 1 decap_w0
xfeed_2430 0 1 decap_w0
xsubckt_928_mux2_x1 0 1 1889 2029 1618 1578 mux2_x1
xsubckt_295_and4_x1 0 1 453 461 457 455 454 and4_x1
xsubckt_418_and21nor_x0 0 1 331 652 629 359 and21nor_x0
xsubckt_1283_and21nor_x0 0 1 1299 753 478 1317 and21nor_x0
xsubckt_1320_or2_x1 0 1 1265 1273 1266 or2_x1
xsubckt_1627_or21nand_x0 0 1 967 1656 1116 693 or21nand_x0
xspare_buffer_45 0 1 60 68 buf_x4
xspare_buffer_46 0 1 59 68 buf_x4
xspare_buffer_47 0 1 13 16 buf_x4
xspare_buffer_48 0 1 58 68 buf_x4
xspare_buffer_49 0 1 57 68 buf_x4
xfeed_7279 0 1 decap_w0
xfeed_7278 0 1 decap_w0
xfeed_7277 0 1 decap_w0
xfeed_6749 0 1 decap_w0
xfeed_6748 0 1 decap_w0
xfeed_6747 0 1 decap_w0
xfeed_6745 0 1 decap_w0
xfeed_6744 0 1 decap_w0
xfeed_6743 0 1 decap_w0
xfeed_6742 0 1 decap_w0
xfeed_6741 0 1 decap_w0
xfeed_6740 0 1 decap_w0
xfeed_2439 0 1 decap_w0
xfeed_2438 0 1 decap_w0
xfeed_1909 0 1 decap_w0
xfeed_1908 0 1 decap_w0
xfeed_1907 0 1 decap_w0
xfeed_1906 0 1 decap_w0
xfeed_1905 0 1 decap_w0
xfeed_1904 0 1 decap_w0
xfeed_1903 0 1 decap_w0
xfeed_1902 0 1 decap_w0
xfeed_1901 0 1 decap_w0
xfeed_1900 0 1 decap_w0
xfeed_419 0 1 decap_w0
xfeed_418 0 1 decap_w0
xfeed_417 0 1 decap_w0
xfeed_416 0 1 decap_w0
xfeed_415 0 1 decap_w0
xfeed_414 0 1 decap_w0
xfeed_413 0 1 decap_w0
xfeed_412 0 1 decap_w0
xfeed_411 0 1 decap_w0
xfeed_410 0 1 decap_w0
xsubckt_1079_and21nor_x0 0 1 1465 1522 1466 533 and21nor_x0
xsubckt_868_nand3_x0 0 1 1614 2052 1962 1617 nand3_x0
xsubckt_247_nand4_x0 0 1 504 712 1926 571 557 nand4_x0
xsubckt_557_or21nand_x0 0 1 198 447 610 616 or21nand_x0
xsubckt_1784_and21nor_x0 0 1 810 1037 1034 1031 and21nor_x0
xspare_buffer_50 0 1 56 68 buf_x4
xspare_buffer_51 0 1 12 16 buf_x4
xfeed_13489 0 1 tie
xfeed_13488 0 1 decap_w0
xfeed_13487 0 1 decap_w0
xfeed_13486 0 1 decap_w0
xfeed_13485 0 1 decap_w0
xfeed_13484 0 1 decap_w0
xfeed_13483 0 1 decap_w0
xfeed_13482 0 1 decap_w0
xfeed_13481 0 1 decap_w0
xfeed_13480 0 1 decap_w0
xfeed_12959 0 1 decap_w0
xfeed_12958 0 1 decap_w0
xfeed_12957 0 1 decap_w0
xfeed_12956 0 1 decap_w0
xfeed_12955 0 1 tie
xfeed_12954 0 1 decap_w0
xfeed_12953 0 1 decap_w0
xfeed_12952 0 1 decap_w0
xfeed_12951 0 1 decap_w0
xfeed_12950 0 1 decap_w0
xfeed_7283 0 1 decap_w0
xfeed_7282 0 1 decap_w0
xfeed_7281 0 1 decap_w0
xfeed_7280 0 1 decap_w0
xfeed_2444 0 1 decap_w0
xfeed_2443 0 1 decap_w0
xfeed_2442 0 1 decap_w0
xfeed_2441 0 1 decap_w0
xfeed_2440 0 1 decap_w0
xsubckt_1160_mux2_x1 0 1 1401 1402 695 484 mux2_x1
xsubckt_125_and4_x1 0 1 643 660 651 648 647 and4_x1
xsubckt_156_or21nand_x0 0 1 605 612 610 616 or21nand_x0
xsubckt_424_nand2_x0 0 1 325 610 460 nand2_x0
xsubckt_1725_nand2_x0 0 1 869 873 871 nand2_x0
xsubckt_1727_or21nand_x0 0 1 867 1105 874 872 or21nand_x0
xspare_buffer_52 0 1 54 55 buf_x4
xspare_buffer_53 0 1 53 55 buf_x4
xspare_buffer_54 0 1 52 55 buf_x4
xspare_buffer_55 0 1 10 11 buf_x4
xspare_buffer_56 0 1 51 55 buf_x4
xspare_buffer_57 0 1 50 55 buf_x4
xspare_buffer_58 0 1 49 55 buf_x4
xspare_buffer_59 0 1 9 11 buf_x4
xfeed_7289 0 1 decap_w0
xfeed_7288 0 1 decap_w0
xfeed_7287 0 1 decap_w0
xfeed_7286 0 1 tie
xfeed_7285 0 1 decap_w0
xfeed_7284 0 1 decap_w0
xfeed_6759 0 1 decap_w0
xfeed_6758 0 1 decap_w0
xfeed_6757 0 1 decap_w0
xfeed_6756 0 1 decap_w0
xfeed_6755 0 1 decap_w0
xfeed_6754 0 1 decap_w0
xfeed_6753 0 1 decap_w0
xfeed_6752 0 1 decap_w0
xfeed_6751 0 1 decap_w0
xfeed_6750 0 1 decap_w0
xfeed_2449 0 1 tie
xfeed_2448 0 1 decap_w0
xfeed_2447 0 1 decap_w0
xfeed_2446 0 1 decap_w0
xfeed_2445 0 1 decap_w0
xfeed_1919 0 1 decap_w0
xfeed_1918 0 1 decap_w0
xfeed_1917 0 1 decap_w0
xfeed_1916 0 1 decap_w0
xfeed_1915 0 1 decap_w0
xfeed_1914 0 1 decap_w0
xfeed_1913 0 1 decap_w0
xfeed_1912 0 1 decap_w0
xfeed_1911 0 1 decap_w0
xfeed_1910 0 1 decap_w0
xfeed_429 0 1 decap_w0
xfeed_428 0 1 decap_w0
xfeed_427 0 1 decap_w0
xfeed_426 0 1 decap_w0
xfeed_425 0 1 decap_w0
xfeed_424 0 1 decap_w0
xfeed_423 0 1 decap_w0
xfeed_422 0 1 decap_w0
xfeed_421 0 1 decap_w0
xfeed_420 0 1 decap_w0
xsubckt_1014_nand3_x0 0 1 1517 643 622 313 nand3_x0
xsubckt_851_nand3_x0 0 1 1628 2066 682 490 nand3_x0
xsubckt_334_nand2_x0 0 1 414 609 418 nand2_x0
xfeed_13499 0 1 tie
xfeed_13498 0 1 decap_w0
xfeed_13497 0 1 decap_w0
xfeed_13496 0 1 decap_w0
xfeed_13495 0 1 decap_w0
xfeed_13494 0 1 decap_w0
xfeed_13493 0 1 decap_w0
xfeed_13492 0 1 decap_w0
xfeed_13491 0 1 decap_w0
xfeed_13490 0 1 decap_w0
xfeed_12969 0 1 decap_w0
xfeed_12968 0 1 decap_w0
xfeed_12967 0 1 decap_w0
xfeed_12966 0 1 decap_w0
xfeed_12965 0 1 decap_w0
xfeed_12964 0 1 decap_w0
xfeed_12963 0 1 decap_w0
xfeed_12962 0 1 decap_w0
xfeed_12961 0 1 decap_w0
xfeed_12960 0 1 tie
xfeed_7290 0 1 decap_w0
xfeed_2451 0 1 decap_w0
xfeed_2450 0 1 decap_w0
xsubckt_1156_mux2_x1 0 1 1404 1996 2046 1408 mux2_x1
xsubckt_991_and4_x1 0 1 1537 638 632 525 520 and4_x1
xsubckt_696_and2_x1 0 1 1768 537 198 and2_x1
xsubckt_1679_mux2_x1 0 1 915 964 917 1142 mux2_x1
xspare_buffer_60 0 1 48 55 buf_x4
xspare_buffer_61 0 1 47 55 buf_x4
xspare_buffer_62 0 1 46 55 buf_x4
xspare_buffer_63 0 1 8 11 buf_x4
xspare_buffer_64 0 1 45 55 buf_x4
xspare_buffer_65 0 1 44 55 buf_x4
xspare_buffer_66 0 1 43 55 buf_x4
xspare_buffer_67 0 1 7 11 buf_x4
xspare_buffer_68 0 1 41 42 buf_x4
xspare_buffer_69 0 1 40 42 buf_x4
xfeed_7299 0 1 decap_w0
xfeed_7298 0 1 decap_w0
xfeed_7296 0 1 decap_w0
xfeed_7295 0 1 decap_w0
xfeed_7294 0 1 decap_w0
xfeed_7293 0 1 tie
xfeed_7292 0 1 decap_w0
xfeed_7291 0 1 decap_w0
xfeed_6769 0 1 decap_w0
xfeed_6768 0 1 decap_w0
xfeed_6767 0 1 decap_w0
xfeed_6766 0 1 decap_w0
xfeed_6765 0 1 decap_w0
xfeed_6764 0 1 decap_w0
xfeed_6763 0 1 decap_w0
xfeed_6762 0 1 decap_w0
xfeed_6761 0 1 decap_w0
xfeed_6760 0 1 decap_w0
xfeed_2459 0 1 decap_w0
xfeed_2458 0 1 decap_w0
xfeed_2457 0 1 decap_w0
xfeed_2456 0 1 decap_w0
xfeed_2455 0 1 decap_w0
xfeed_2454 0 1 decap_w0
xfeed_2453 0 1 decap_w0
xfeed_2452 0 1 decap_w0
xfeed_1929 0 1 decap_w0
xfeed_1928 0 1 decap_w0
xfeed_1927 0 1 decap_w0
xfeed_1926 0 1 decap_w0
xfeed_1925 0 1 tie
xfeed_1924 0 1 decap_w0
xfeed_1923 0 1 decap_w0
xfeed_1922 0 1 decap_w0
xfeed_1921 0 1 decap_w0
xfeed_1920 0 1 decap_w0
xfeed_439 0 1 decap_w0
xfeed_438 0 1 tie
xfeed_437 0 1 decap_w0
xfeed_436 0 1 decap_w0
xfeed_435 0 1 decap_w0
xfeed_434 0 1 decap_w0
xfeed_433 0 1 decap_w0
xfeed_432 0 1 decap_w0
xfeed_431 0 1 decap_w0
xfeed_430 0 1 decap_w0
xsubckt_757_or21nand_x0 0 1 1711 1766 116 119 or21nand_x0
xsubckt_169_and2_x1 0 1 589 1929 1924 and2_x1
xfeed_12979 0 1 decap_w0
xfeed_12978 0 1 decap_w0
xfeed_12977 0 1 decap_w0
xfeed_12976 0 1 decap_w0
xfeed_12975 0 1 decap_w0
xfeed_12974 0 1 decap_w0
xfeed_12973 0 1 decap_w0
xfeed_12972 0 1 decap_w0
xfeed_12971 0 1 decap_w0
xfeed_12970 0 1 decap_w0
xsubckt_1587_mux2_x1 0 1 1007 1008 1013 1020 mux2_x1
xspare_buffer_70 0 1 39 42 buf_x4
xspare_buffer_71 0 1 5 6 buf_x4
xspare_buffer_72 0 1 38 42 buf_x4
xspare_buffer_73 0 1 37 42 buf_x4
xspare_buffer_74 0 1 36 42 buf_x4
xspare_buffer_75 0 1 4 6 buf_x4
xspare_buffer_76 0 1 35 42 buf_x4
xspare_buffer_77 0 1 34 42 buf_x4
xspare_buffer_78 0 1 33 42 buf_x4
xspare_buffer_79 0 1 3 6 buf_x4
xcmpt_abc_11867_new_n431_hfns_0 0 1 666 664 buf_x4
xcmpt_abc_11867_new_n431_hfns_1 0 1 665 664 buf_x4
xcmpt_abc_11867_new_n431_hfns_2 0 1 664 667 buf_x4
xcmpt_abc_11867_new_n433_hfns_0 0 1 661 658 buf_x4
xcmpt_abc_11867_new_n433_hfns_1 0 1 660 658 buf_x4
xcmpt_abc_11867_new_n433_hfns_2 0 1 659 658 buf_x4
xcmpt_abc_11867_new_n433_hfns_3 0 1 658 662 buf_x4
xfeed_6779 0 1 decap_w0
xfeed_6778 0 1 decap_w0
xfeed_6777 0 1 decap_w0
xfeed_6776 0 1 decap_w0
xfeed_6775 0 1 decap_w0
xfeed_6774 0 1 tie
xfeed_6773 0 1 decap_w0
xfeed_6772 0 1 decap_w0
xfeed_6771 0 1 decap_w0
xfeed_6770 0 1 decap_w0
xfeed_2469 0 1 decap_w0
xfeed_2468 0 1 decap_w0
xfeed_2467 0 1 decap_w0
xfeed_2466 0 1 decap_w0
xfeed_2465 0 1 decap_w0
xfeed_2464 0 1 decap_w0
xfeed_2463 0 1 decap_w0
xfeed_2462 0 1 decap_w0
xfeed_2461 0 1 decap_w0
xfeed_2460 0 1 decap_w0
xfeed_1939 0 1 decap_w0
xfeed_1938 0 1 decap_w0
xfeed_1937 0 1 decap_w0
xfeed_1936 0 1 decap_w0
xfeed_1935 0 1 decap_w0
xfeed_1934 0 1 decap_w0
xfeed_1933 0 1 decap_w0
xfeed_1932 0 1 decap_w0
xfeed_1931 0 1 decap_w0
xfeed_1930 0 1 decap_w0
xfeed_449 0 1 decap_w0
xfeed_448 0 1 tie
xfeed_447 0 1 decap_w0
xfeed_446 0 1 decap_w0
xfeed_445 0 1 decap_w0
xfeed_444 0 1 decap_w0
xfeed_443 0 1 decap_w0
xfeed_442 0 1 decap_w0
xfeed_441 0 1 decap_w0
xfeed_440 0 1 decap_w0
xsubckt_577_nand4_x0 0 1 178 1932 195 194 189 nand4_x0
xsubckt_621_and21nor_x0 0 1 136 753 449 410 and21nor_x0
xfeed_12989 0 1 tie
xfeed_12988 0 1 decap_w0
xfeed_12987 0 1 decap_w0
xfeed_12986 0 1 decap_w0
xfeed_12985 0 1 decap_w0
xfeed_12984 0 1 decap_w0
xfeed_12983 0 1 decap_w0
xfeed_12982 0 1 decap_w0
xfeed_12981 0 1 decap_w0
xfeed_12980 0 1 decap_w0
xsubckt_1255_and3_x1 0 1 1325 284 1329 1326 and3_x1
xsubckt_760_or21nand_x0 0 1 1708 2061 1742 1740 or21nand_x0
xsubckt_754_nand2_x0 0 1 1713 1715 1714 nand2_x0
xsubckt_320_and3_x1 0 1 428 650 644 533 and3_x1
xsubckt_1921_dff_x1 0 1 2062 1827 35 dff_x1
xspare_buffer_80 0 1 32 42 buf_x4
xspare_buffer_81 0 1 31 42 buf_x4
xspare_buffer_82 0 1 30 42 buf_x4
xspare_buffer_83 0 1 2 6 buf_x4
xfeed_6789 0 1 decap_w0
xfeed_6788 0 1 tie
xfeed_6787 0 1 decap_w0
xfeed_6786 0 1 decap_w0
xfeed_6785 0 1 decap_w0
xfeed_6784 0 1 decap_w0
xfeed_6783 0 1 decap_w0
xfeed_6782 0 1 decap_w0
xfeed_6781 0 1 tie
xfeed_6780 0 1 decap_w0
xfeed_2479 0 1 decap_w0
xfeed_2478 0 1 decap_w0
xfeed_2477 0 1 decap_w0
xfeed_2476 0 1 decap_w0
xfeed_2475 0 1 decap_w0
xfeed_2474 0 1 decap_w0
xfeed_2473 0 1 decap_w0
xfeed_2472 0 1 tie
xfeed_2471 0 1 decap_w0
xfeed_2470 0 1 decap_w0
xfeed_1949 0 1 decap_w0
xfeed_1948 0 1 decap_w0
xfeed_1947 0 1 decap_w0
xfeed_1946 0 1 decap_w0
xfeed_1945 0 1 decap_w0
xfeed_1944 0 1 decap_w0
xfeed_1943 0 1 decap_w0
xfeed_1942 0 1 decap_w0
xfeed_1941 0 1 decap_w0
xfeed_1940 0 1 decap_w0
xfeed_459 0 1 decap_w0
xfeed_458 0 1 decap_w0
xfeed_457 0 1 decap_w0
xfeed_456 0 1 decap_w0
xfeed_455 0 1 decap_w0
xfeed_454 0 1 decap_w0
xfeed_453 0 1 tie
xfeed_452 0 1 decap_w0
xfeed_451 0 1 decap_w0
xfeed_450 0 1 decap_w0
xsubckt_280_and4_x1 0 1 468 1925 711 599 589 and4_x1
xsubckt_1923_dff_x1 0 1 2060 1825 38 dff_x1
xsubckt_1925_dff_x1 0 1 2058 1823 38 dff_x1
xsubckt_1927_dff_x1 0 1 2072 1821 61 dff_x1
xfeed_13609 0 1 decap_w0
xfeed_13608 0 1 decap_w0
xfeed_13607 0 1 decap_w0
xfeed_13606 0 1 decap_w0
xfeed_13605 0 1 decap_w0
xfeed_13604 0 1 decap_w0
xfeed_13603 0 1 decap_w0
xfeed_13602 0 1 decap_w0
xfeed_13601 0 1 decap_w0
xfeed_13600 0 1 decap_w0
xfeed_12999 0 1 decap_w0
xfeed_12998 0 1 decap_w0
xfeed_12997 0 1 decap_w0
xfeed_12996 0 1 decap_w0
xfeed_12995 0 1 decap_w0
xfeed_12994 0 1 decap_w0
xfeed_12993 0 1 decap_w0
xfeed_12992 0 1 decap_w0
xfeed_12991 0 1 decap_w0
xfeed_12990 0 1 decap_w0
xfeed_7409 0 1 decap_w0
xfeed_7408 0 1 decap_w0
xfeed_7407 0 1 decap_w0
xfeed_7406 0 1 decap_w0
xfeed_7405 0 1 decap_w0
xfeed_7404 0 1 decap_w0
xfeed_7403 0 1 decap_w0
xfeed_7402 0 1 decap_w0
xfeed_7401 0 1 decap_w0
xfeed_7400 0 1 decap_w0
xsubckt_913_mux2_x1 0 1 1902 1600 2042 1580 mux2_x1
xsubckt_839_and3_x1 0 1 1639 1976 1749 1739 and3_x1
xsubckt_725_and4_x1 0 1 1739 1767 1747 1743 1741 and4_x1
xsubckt_316_and3_x1 0 1 432 443 440 433 and3_x1
xsubckt_202_and4_x1 0 1 552 1925 711 673 669 and4_x1
xsubckt_394_nand2_x0 0 1 355 535 357 nand2_x0
xsubckt_1881_dff_x1 0 1 1963 1858 67 dff_x1
xsubckt_1883_dff_x1 0 1 1947 1856 77 dff_x1
xsubckt_1929_dff_x1 0 1 2070 1819 64 dff_x1
xfeed_6799 0 1 tie
xfeed_6798 0 1 decap_w0
xfeed_6797 0 1 decap_w0
xfeed_6796 0 1 decap_w0
xfeed_6795 0 1 decap_w0
xfeed_6794 0 1 decap_w0
xfeed_6793 0 1 decap_w0
xfeed_6791 0 1 decap_w0
xfeed_6790 0 1 decap_w0
xfeed_2489 0 1 decap_w0
xfeed_2488 0 1 decap_w0
xfeed_2487 0 1 decap_w0
xfeed_2486 0 1 decap_w0
xfeed_2485 0 1 decap_w0
xfeed_2484 0 1 decap_w0
xfeed_2483 0 1 decap_w0
xfeed_2482 0 1 decap_w0
xfeed_2481 0 1 decap_w0
xfeed_2480 0 1 decap_w0
xfeed_1959 0 1 tie
xfeed_1958 0 1 decap_w0
xfeed_1957 0 1 decap_w0
xfeed_1956 0 1 decap_w0
xfeed_1955 0 1 decap_w0
xfeed_1954 0 1 decap_w0
xfeed_1953 0 1 decap_w0
xfeed_1952 0 1 tie
xfeed_1951 0 1 decap_w0
xfeed_1950 0 1 decap_w0
xfeed_469 0 1 decap_w0
xfeed_468 0 1 decap_w0
xfeed_467 0 1 decap_w0
xfeed_466 0 1 decap_w0
xfeed_465 0 1 decap_w0
xfeed_464 0 1 decap_w0
xfeed_463 0 1 decap_w0
xfeed_462 0 1 decap_w0
xfeed_461 0 1 decap_w0
xfeed_460 0 1 decap_w0
xsubckt_1221_nor4_x0 0 1 1343 538 199 1753 1344 nor4_x0
xsubckt_1111_and2_x1 0 1 1438 771 1440 and2_x1
xsubckt_960_or21nand_x0 0 1 1873 1564 1562 1570 or21nand_x0
xsubckt_1594_and3_x1 0 1 1000 1070 1018 1016 and3_x1
xsubckt_1885_dff_x1 0 1 1921 1854 80 dff_x1
xsubckt_1887_dff_x1 0 1 1932 1852 67 dff_x1
xsubckt_1889_dff_x1 0 1 1951 1850 77 dff_x1
xfeed_13619 0 1 decap_w0
xfeed_13618 0 1 decap_w0
xfeed_13617 0 1 decap_w0
xfeed_13616 0 1 decap_w0
xfeed_13615 0 1 decap_w0
xfeed_13614 0 1 decap_w0
xfeed_13613 0 1 decap_w0
xfeed_13612 0 1 decap_w0
xfeed_13611 0 1 tie
xfeed_13610 0 1 decap_w0
xfeed_7416 0 1 decap_w0
xfeed_7415 0 1 tie
xfeed_7414 0 1 decap_w0
xfeed_7413 0 1 decap_w0
xfeed_7412 0 1 decap_w0
xfeed_7411 0 1 decap_w0
xfeed_7410 0 1 decap_w0
xfeed_3109 0 1 decap_w0
xfeed_3108 0 1 decap_w0
xfeed_3107 0 1 decap_w0
xfeed_3106 0 1 decap_w0
xfeed_3105 0 1 decap_w0
xfeed_3104 0 1 decap_w0
xfeed_3103 0 1 decap_w0
xfeed_3102 0 1 decap_w0
xfeed_3101 0 1 decap_w0
xfeed_3100 0 1 decap_w0
xsubckt_1233_mux2_x1 0 1 1828 2098 2063 1334 mux2_x1
xsubckt_1107_and2_x1 0 1 1441 1917 1442 and2_x1
xfeed_7419 0 1 decap_w0
xfeed_7418 0 1 decap_w0
xfeed_7417 0 1 decap_w0
xfeed_2499 0 1 decap_w0
xfeed_2498 0 1 decap_w0
xfeed_2497 0 1 decap_w0
xfeed_2496 0 1 decap_w0
xfeed_2495 0 1 decap_w0
xfeed_2494 0 1 decap_w0
xfeed_2493 0 1 decap_w0
xfeed_2492 0 1 decap_w0
xfeed_2491 0 1 decap_w0
xfeed_2490 0 1 decap_w0
xfeed_1969 0 1 decap_w0
xfeed_1968 0 1 decap_w0
xfeed_1967 0 1 decap_w0
xfeed_1966 0 1 decap_w0
xfeed_1965 0 1 decap_w0
xfeed_1964 0 1 tie
xfeed_1963 0 1 decap_w0
xfeed_1962 0 1 decap_w0
xfeed_1961 0 1 decap_w0
xfeed_1960 0 1 decap_w0
xfeed_479 0 1 decap_w0
xfeed_478 0 1 decap_w0
xfeed_477 0 1 decap_w0
xfeed_476 0 1 decap_w0
xfeed_475 0 1 decap_w0
xfeed_474 0 1 decap_w0
xfeed_473 0 1 tie
xfeed_472 0 1 decap_w0
xfeed_471 0 1 decap_w0
xfeed_470 0 1 decap_w0
xsubckt_1247_nand2_x0 0 1 1333 775 1982 nand2_x0
xsubckt_769_and2_x1 0 1 1700 1702 1701 and2_x1
xsubckt_629_and4_x1 0 1 129 133 132 131 130 and4_x1
xsubckt_1481_or2_x1 0 1 1115 689 1116 or2_x1
xfeed_13629 0 1 decap_w0
xfeed_13628 0 1 decap_w0
xfeed_13627 0 1 decap_w0
xfeed_13626 0 1 decap_w0
xfeed_13625 0 1 decap_w0
xfeed_13624 0 1 decap_w0
xfeed_13623 0 1 decap_w0
xfeed_13622 0 1 decap_w0
xfeed_13621 0 1 decap_w0
xfeed_13620 0 1 decap_w0
xfeed_7423 0 1 decap_w0
xfeed_7422 0 1 tie
xfeed_7421 0 1 decap_w0
xfeed_7420 0 1 decap_w0
xfeed_3119 0 1 decap_w0
xfeed_3118 0 1 decap_w0
xfeed_3117 0 1 decap_w0
xfeed_3116 0 1 decap_w0
xfeed_3115 0 1 decap_w0
xfeed_3114 0 1 decap_w0
xfeed_3113 0 1 decap_w0
xfeed_3112 0 1 decap_w0
xfeed_3111 0 1 decap_w0
xfeed_3110 0 1 decap_w0
xsubckt_1141_mux2_x1 0 1 1417 1418 2001 484 mux2_x1
xsubckt_980_nand4_x0 0 1 1547 637 633 622 520 nand4_x0
xsubckt_717_and21nor_x0 0 1 1747 570 460 617 and21nor_x0
xsubckt_681_and2_x1 0 1 1782 1784 1783 and2_x1
xsubckt_549_nand4_x0 0 1 205 716 1924 1926 599 nand4_x0
xsubckt_1779_and21nor_x0 0 1 815 1005 1002 999 and21nor_x0
xfeed_7429 0 1 decap_w0
xfeed_7428 0 1 decap_w0
xfeed_7427 0 1 tie
xfeed_7426 0 1 decap_w0
xfeed_7425 0 1 decap_w0
xfeed_7424 0 1 decap_w0
xfeed_1979 0 1 decap_w0
xfeed_1978 0 1 decap_w0
xfeed_1977 0 1 decap_w0
xfeed_1976 0 1 decap_w0
xfeed_1975 0 1 tie
xfeed_1974 0 1 decap_w0
xfeed_1973 0 1 decap_w0
xfeed_1972 0 1 decap_w0
xfeed_1971 0 1 tie
xfeed_1970 0 1 decap_w0
xfeed_489 0 1 decap_w0
xfeed_488 0 1 decap_w0
xfeed_487 0 1 tie
xfeed_486 0 1 decap_w0
xfeed_485 0 1 decap_w0
xfeed_484 0 1 decap_w0
xfeed_483 0 1 decap_w0
xfeed_482 0 1 decap_w0
xfeed_481 0 1 decap_w0
xfeed_480 0 1 tie
xsubckt_154_and2_x1 0 1 611 1925 711 and2_x1
xsubckt_537_and4_x1 0 1 216 507 463 219 217 and4_x1
xsubckt_1682_and21nor_x0 0 1 912 913 916 1076 and21nor_x0
xfeed_13639 0 1 decap_w0
xfeed_13638 0 1 decap_w0
xfeed_13637 0 1 decap_w0
xfeed_13636 0 1 decap_w0
xfeed_13635 0 1 decap_w0
xfeed_13634 0 1 decap_w0
xfeed_13633 0 1 decap_w0
xfeed_13632 0 1 decap_w0
xfeed_13631 0 1 decap_w0
xfeed_13630 0 1 decap_w0
xfeed_7430 0 1 decap_w0
xfeed_3129 0 1 decap_w0
xfeed_3128 0 1 decap_w0
xfeed_3127 0 1 decap_w0
xfeed_3126 0 1 decap_w0
xfeed_3125 0 1 decap_w0
xfeed_3124 0 1 decap_w0
xfeed_3123 0 1 decap_w0
xfeed_3122 0 1 decap_w0
xfeed_3121 0 1 decap_w0
xfeed_3120 0 1 decap_w0
xsubckt_0_inv_x0 0 1 786 1995 inv_x0
xsubckt_2_inv_x0 0 1 784 1939 inv_x0
xsubckt_4_inv_x0 0 1 782 1983 inv_x0
xsubckt_1316_nand3_x0 0 1 1269 2060 666 657 nand3_x0
xfeed_7439 0 1 decap_w0
xfeed_7438 0 1 decap_w0
xfeed_7436 0 1 decap_w0
xfeed_7435 0 1 decap_w0
xfeed_7434 0 1 tie
xfeed_7433 0 1 decap_w0
xfeed_7432 0 1 decap_w0
xfeed_7431 0 1 decap_w0
xfeed_6909 0 1 decap_w0
xfeed_6908 0 1 decap_w0
xfeed_6907 0 1 decap_w0
xfeed_6906 0 1 decap_w0
xfeed_6905 0 1 decap_w0
xfeed_6904 0 1 decap_w0
xfeed_6903 0 1 decap_w0
xfeed_6902 0 1 decap_w0
xfeed_6901 0 1 decap_w0
xfeed_6900 0 1 tie
xfeed_1989 0 1 decap_w0
xfeed_1988 0 1 decap_w0
xfeed_1987 0 1 tie
xfeed_1986 0 1 decap_w0
xfeed_1985 0 1 decap_w0
xfeed_1984 0 1 decap_w0
xfeed_1983 0 1 decap_w0
xfeed_1982 0 1 decap_w0
xfeed_1981 0 1 decap_w0
xfeed_1980 0 1 decap_w0
xfeed_499 0 1 decap_w0
xfeed_498 0 1 decap_w0
xfeed_497 0 1 decap_w0
xfeed_496 0 1 decap_w0
xfeed_495 0 1 decap_w0
xfeed_494 0 1 decap_w0
xfeed_493 0 1 decap_w0
xfeed_492 0 1 decap_w0
xfeed_491 0 1 decap_w0
xfeed_490 0 1 decap_w0
xsubckt_956_or21nand_x0 0 1 1874 1568 1565 1573 or21nand_x0
xsubckt_6_inv_x0 0 1 780 1940 inv_x0
xsubckt_8_inv_x0 0 1 778 1920 inv_x0
xsubckt_445_and4_x1 0 1 305 628 620 516 306 and4_x1
xsubckt_1782_and21nor_x0 0 1 812 997 816 814 and21nor_x0
xfeed_13649 0 1 decap_w0
xfeed_13648 0 1 decap_w0
xfeed_13647 0 1 decap_w0
xfeed_13646 0 1 decap_w0
xfeed_13645 0 1 decap_w0
xfeed_13644 0 1 decap_w0
xfeed_13643 0 1 decap_w0
xfeed_13642 0 1 decap_w0
xfeed_13641 0 1 decap_w0
xfeed_13640 0 1 decap_w0
xfeed_3137 0 1 decap_w0
xfeed_3136 0 1 decap_w0
xfeed_3135 0 1 decap_w0
xfeed_3134 0 1 decap_w0
xfeed_3133 0 1 decap_w0
xfeed_3132 0 1 decap_w0
xfeed_3131 0 1 decap_w0
xfeed_3130 0 1 decap_w0
xfeed_7449 0 1 decap_w0
xfeed_7448 0 1 decap_w0
xfeed_7447 0 1 decap_w0
xfeed_7446 0 1 decap_w0
xfeed_7445 0 1 decap_w0
xfeed_7444 0 1 decap_w0
xfeed_7443 0 1 decap_w0
xfeed_7442 0 1 decap_w0
xfeed_7441 0 1 tie
xfeed_7440 0 1 decap_w0
xfeed_6919 0 1 decap_w0
xfeed_6918 0 1 decap_w0
xfeed_6917 0 1 decap_w0
xfeed_6916 0 1 decap_w0
xfeed_6915 0 1 decap_w0
xfeed_6914 0 1 decap_w0
xfeed_6913 0 1 decap_w0
xfeed_6912 0 1 decap_w0
xfeed_6911 0 1 decap_w0
xfeed_6910 0 1 decap_w0
xfeed_3139 0 1 decap_w0
xfeed_3138 0 1 decap_w0
xfeed_2609 0 1 decap_w0
xfeed_2608 0 1 decap_w0
xfeed_2607 0 1 tie
xfeed_2606 0 1 decap_w0
xfeed_2605 0 1 decap_w0
xfeed_2604 0 1 decap_w0
xfeed_2603 0 1 decap_w0
xfeed_2602 0 1 decap_w0
xfeed_2601 0 1 decap_w0
xfeed_2600 0 1 tie
xfeed_1999 0 1 decap_w0
xfeed_1998 0 1 decap_w0
xfeed_1997 0 1 decap_w0
xfeed_1996 0 1 tie
xfeed_1995 0 1 decap_w0
xfeed_1994 0 1 decap_w0
xfeed_1993 0 1 decap_w0
xfeed_1992 0 1 decap_w0
xfeed_1991 0 1 decap_w0
xfeed_1990 0 1 decap_w0
xsubckt_820_and21nor_x0 0 1 1655 744 600 1745 and21nor_x0
xsubckt_1487_nand2_x0 0 1 1109 1119 1112 nand2_x0
xfeed_13659 0 1 decap_w0
xfeed_13658 0 1 decap_w0
xfeed_13657 0 1 decap_w0
xfeed_13656 0 1 decap_w0
xfeed_13655 0 1 decap_w0
xfeed_13654 0 1 decap_w0
xfeed_13653 0 1 decap_w0
xfeed_13652 0 1 decap_w0
xfeed_13651 0 1 decap_w0
xfeed_13650 0 1 decap_w0
xfeed_3144 0 1 decap_w0
xfeed_3143 0 1 decap_w0
xfeed_3142 0 1 decap_w0
xfeed_3141 0 1 decap_w0
xfeed_3140 0 1 decap_w0
xfeed_7459 0 1 decap_w0
xfeed_7458 0 1 decap_w0
xfeed_7457 0 1 decap_w0
xfeed_7456 0 1 tie
xfeed_7455 0 1 decap_w0
xfeed_7454 0 1 decap_w0
xfeed_7453 0 1 decap_w0
xfeed_7452 0 1 decap_w0
xfeed_7451 0 1 decap_w0
xfeed_7450 0 1 decap_w0
xfeed_6929 0 1 decap_w0
xfeed_6928 0 1 decap_w0
xfeed_6927 0 1 decap_w0
xfeed_6926 0 1 decap_w0
xfeed_6925 0 1 decap_w0
xfeed_6924 0 1 tie
xfeed_6923 0 1 decap_w0
xfeed_6922 0 1 decap_w0
xfeed_6921 0 1 decap_w0
xfeed_6920 0 1 decap_w0
xfeed_3149 0 1 decap_w0
xfeed_3148 0 1 decap_w0
xfeed_3147 0 1 decap_w0
xfeed_3146 0 1 decap_w0
xfeed_3145 0 1 decap_w0
xfeed_2619 0 1 decap_w0
xfeed_2618 0 1 decap_w0
xfeed_2617 0 1 tie
xfeed_2616 0 1 decap_w0
xfeed_2615 0 1 decap_w0
xfeed_2614 0 1 decap_w0
xfeed_2613 0 1 decap_w0
xfeed_2612 0 1 decap_w0
xfeed_2611 0 1 decap_w0
xfeed_2610 0 1 decap_w0
xsubckt_1277_and21nor_x0 0 1 1304 1305 1321 2052 and21nor_x0
xsubckt_1025_nand4_x0 0 1 1509 1916 1927 679 674 nand4_x0
xsubckt_966_nand2_x0 0 1 1558 1935 1575 nand2_x0
xsubckt_830_or2_x1 0 1 2102 1653 1647 or2_x1
xsubckt_1434_nor2_x0 0 1 1160 1165 1161 nor2_x0
xfeed_13669 0 1 decap_w0
xfeed_13668 0 1 decap_w0
xfeed_13667 0 1 decap_w0
xfeed_13666 0 1 decap_w0
xfeed_13665 0 1 decap_w0
xfeed_13664 0 1 decap_w0
xfeed_13663 0 1 decap_w0
xfeed_13662 0 1 decap_w0
xfeed_13661 0 1 decap_w0
xfeed_13660 0 1 decap_w0
xfeed_3151 0 1 decap_w0
xfeed_3150 0 1 decap_w0
xsubckt_1581_and21nor_x0 0 1 1013 1104 1018 1016 and21nor_x0
xfeed_7469 0 1 decap_w0
xfeed_7468 0 1 decap_w0
xfeed_7467 0 1 decap_w0
xfeed_7466 0 1 decap_w0
xfeed_7465 0 1 decap_w0
xfeed_7464 0 1 decap_w0
xfeed_7463 0 1 decap_w0
xfeed_7462 0 1 decap_w0
xfeed_7461 0 1 decap_w0
xfeed_7460 0 1 tie
xfeed_6939 0 1 decap_w0
xfeed_6938 0 1 decap_w0
xfeed_6937 0 1 decap_w0
xfeed_6936 0 1 decap_w0
xfeed_6935 0 1 decap_w0
xfeed_6934 0 1 decap_w0
xfeed_6933 0 1 decap_w0
xfeed_6932 0 1 tie
xfeed_6931 0 1 decap_w0
xfeed_6930 0 1 decap_w0
xfeed_3159 0 1 decap_w0
xfeed_3158 0 1 decap_w0
xfeed_3157 0 1 decap_w0
xfeed_3156 0 1 decap_w0
xfeed_3155 0 1 tie
xfeed_3154 0 1 decap_w0
xfeed_3153 0 1 decap_w0
xfeed_3152 0 1 decap_w0
xfeed_2629 0 1 tie
xfeed_2628 0 1 decap_w0
xfeed_2627 0 1 decap_w0
xfeed_2626 0 1 decap_w0
xfeed_2625 0 1 decap_w0
xfeed_2624 0 1 decap_w0
xfeed_2623 0 1 decap_w0
xfeed_2622 0 1 decap_w0
xfeed_2621 0 1 decap_w0
xfeed_2620 0 1 decap_w0
xfeed_609 0 1 decap_w0
xfeed_608 0 1 decap_w0
xfeed_607 0 1 decap_w0
xfeed_606 0 1 decap_w0
xfeed_605 0 1 decap_w0
xfeed_604 0 1 decap_w0
xfeed_603 0 1 decap_w0
xfeed_602 0 1 decap_w0
xfeed_601 0 1 decap_w0
xfeed_600 0 1 decap_w0
xsubckt_838_or2_x1 0 1 2101 1646 1640 or2_x1
xsubckt_786_nand2_x0 0 1 1685 1687 1686 nand2_x0
xsubckt_283_and3_x1 0 1 465 1920 1917 771 and3_x1
xsubckt_231_and2_x1 0 1 520 661 521 and2_x1
xsubckt_1466_nand3_x0 0 1 1130 1929 610 452 nand3_x0
xsubckt_1575_and3_x1 0 1 1019 1971 679 594 and3_x1
xsubckt_1689_and2_x1 0 1 905 1670 906 and2_x1
xfeed_13679 0 1 decap_w0
xfeed_13678 0 1 decap_w0
xfeed_13677 0 1 decap_w0
xfeed_13676 0 1 decap_w0
xfeed_13675 0 1 decap_w0
xfeed_13674 0 1 decap_w0
xfeed_13673 0 1 decap_w0
xfeed_13672 0 1 decap_w0
xfeed_13671 0 1 decap_w0
xfeed_13670 0 1 decap_w0
xsubckt_816_and21nor_x0 0 1 1659 693 1755 1754 and21nor_x0
xsubckt_798_or2_x1 0 1 2092 1683 1675 or2_x1
xsubckt_279_and3_x1 0 1 469 507 496 470 and3_x1
xsubckt_165_and4_x1 0 1 596 716 1924 714 1928 and4_x1
xsubckt_14_inv_x0 0 1 768 2052 inv_x0
xsubckt_12_inv_x0 0 1 770 1958 inv_x0
xsubckt_10_inv_x0 0 1 776 1917 inv_x0
xsubckt_428_nand2_x0 0 1 321 323 322 nand2_x0
xsubckt_1286_nand3_x0 0 1 1296 679 447 1297 nand3_x0
xsubckt_1523_and2_x1 0 1 1073 1081 1077 and2_x1
xfeed_7478 0 1 decap_w0
xfeed_7477 0 1 decap_w0
xfeed_7476 0 1 decap_w0
xfeed_7475 0 1 decap_w0
xfeed_7474 0 1 decap_w0
xfeed_7473 0 1 decap_w0
xfeed_7472 0 1 decap_w0
xfeed_7471 0 1 decap_w0
xfeed_7470 0 1 decap_w0
xfeed_6949 0 1 decap_w0
xfeed_6948 0 1 decap_w0
xfeed_6947 0 1 tie
xfeed_6946 0 1 decap_w0
xfeed_6945 0 1 decap_w0
xfeed_6944 0 1 decap_w0
xfeed_6943 0 1 decap_w0
xfeed_6942 0 1 decap_w0
xfeed_6941 0 1 decap_w0
xfeed_6940 0 1 decap_w0
xfeed_3169 0 1 decap_w0
xfeed_3168 0 1 decap_w0
xfeed_3167 0 1 decap_w0
xfeed_3166 0 1 decap_w0
xfeed_3165 0 1 decap_w0
xfeed_3164 0 1 decap_w0
xfeed_3163 0 1 decap_w0
xfeed_3162 0 1 decap_w0
xfeed_3161 0 1 decap_w0
xfeed_3160 0 1 decap_w0
xfeed_2639 0 1 decap_w0
xfeed_2638 0 1 tie
xfeed_2637 0 1 decap_w0
xfeed_2636 0 1 decap_w0
xfeed_2635 0 1 decap_w0
xfeed_2634 0 1 decap_w0
xfeed_2633 0 1 decap_w0
xfeed_2632 0 1 decap_w0
xfeed_2631 0 1 decap_w0
xfeed_2630 0 1 decap_w0
xfeed_619 0 1 decap_w0
xfeed_618 0 1 decap_w0
xfeed_617 0 1 decap_w0
xfeed_616 0 1 decap_w0
xfeed_615 0 1 decap_w0
xfeed_614 0 1 decap_w0
xfeed_613 0 1 decap_w0
xfeed_612 0 1 decap_w0
xfeed_611 0 1 decap_w0
xfeed_610 0 1 decap_w0
xsubckt_1074_and2_x1 0 1 1469 1471 1470 and2_x1
xsubckt_18_inv_x0 0 1 764 2050 inv_x0
xsubckt_16_inv_x0 0 1 766 2054 inv_x0
xsubckt_338_nand2_x0 0 1 410 682 421 nand2_x0
xsubckt_522_and4_x1 0 1 230 504 502 492 486 and4_x1
xsubckt_636_and3_x1 0 1 122 127 126 123 and3_x1
xsubckt_1645_mux2_x1 0 1 949 955 952 964 mux2_x1
xsubckt_1688_or2_x1 0 1 906 695 1116 or2_x1
xfeed_13689 0 1 decap_w0
xfeed_13688 0 1 decap_w0
xfeed_13687 0 1 decap_w0
xfeed_13686 0 1 decap_w0
xfeed_13685 0 1 decap_w0
xfeed_13684 0 1 tie
xfeed_13683 0 1 decap_w0
xfeed_13682 0 1 decap_w0
xfeed_13681 0 1 decap_w0
xfeed_13680 0 1 decap_w0
xsubckt_248_nand2_x0 0 1 503 617 603 nand2_x0
xsubckt_1802_nand2_x0 0 1 1797 1061 793 nand2_x0
xfeed_7489 0 1 decap_w0
xfeed_7488 0 1 decap_w0
xfeed_7487 0 1 decap_w0
xfeed_7486 0 1 decap_w0
xfeed_7485 0 1 decap_w0
xfeed_7484 0 1 decap_w0
xfeed_7483 0 1 decap_w0
xfeed_7482 0 1 decap_w0
xfeed_7481 0 1 decap_w0
xfeed_7480 0 1 tie
xfeed_6959 0 1 decap_w0
xfeed_6958 0 1 decap_w0
xfeed_6957 0 1 decap_w0
xfeed_6956 0 1 decap_w0
xfeed_6955 0 1 decap_w0
xfeed_6954 0 1 decap_w0
xfeed_6953 0 1 decap_w0
xfeed_6952 0 1 tie
xfeed_6951 0 1 decap_w0
xfeed_6950 0 1 decap_w0
xfeed_3179 0 1 decap_w0
xfeed_3178 0 1 decap_w0
xfeed_3177 0 1 decap_w0
xfeed_3176 0 1 decap_w0
xfeed_3175 0 1 decap_w0
xfeed_3174 0 1 decap_w0
xfeed_3173 0 1 decap_w0
xfeed_3172 0 1 decap_w0
xfeed_3171 0 1 decap_w0
xfeed_3170 0 1 decap_w0
xfeed_2649 0 1 decap_w0
xfeed_2648 0 1 decap_w0
xfeed_2647 0 1 decap_w0
xfeed_2646 0 1 decap_w0
xfeed_2645 0 1 decap_w0
xfeed_2644 0 1 decap_w0
xfeed_2643 0 1 decap_w0
xfeed_2642 0 1 decap_w0
xfeed_2641 0 1 decap_w0
xfeed_2640 0 1 decap_w0
xfeed_629 0 1 decap_w0
xfeed_628 0 1 decap_w0
xfeed_627 0 1 decap_w0
xfeed_626 0 1 decap_w0
xfeed_625 0 1 decap_w0
xfeed_624 0 1 decap_w0
xfeed_623 0 1 decap_w0
xfeed_622 0 1 decap_w0
xfeed_621 0 1 decap_w0
xfeed_620 0 1 decap_w0
xsubckt_1118_mux2_x1 0 1 1839 1997 1988 1438 mux2_x1
xsubckt_135_and2_x1 0 1 633 661 634 and2_x1
xsubckt_570_and2_x1 0 1 185 191 186 and2_x1
xsubckt_1722_and4_x1 0 1 872 2003 1128 1098 1097 and4_x1
xfeed_13699 0 1 decap_w0
xfeed_13698 0 1 decap_w0
xfeed_13697 0 1 tie
xfeed_13696 0 1 decap_w0
xfeed_13695 0 1 decap_w0
xfeed_13694 0 1 decap_w0
xfeed_13693 0 1 decap_w0
xfeed_13692 0 1 decap_w0
xfeed_13691 0 1 decap_w0
xfeed_13690 0 1 decap_w0
xfeed_8109 0 1 decap_w0
xfeed_8108 0 1 decap_w0
xfeed_8107 0 1 decap_w0
xfeed_8106 0 1 decap_w0
xfeed_8105 0 1 decap_w0
xfeed_8104 0 1 decap_w0
xfeed_8103 0 1 decap_w0
xfeed_8102 0 1 decap_w0
xfeed_8101 0 1 decap_w0
xfeed_8100 0 1 decap_w0
xsubckt_869_nexor2_x0 0 1 1613 768 1616 nexor2_x0
xsubckt_407_nand3_x0 0 1 342 608 558 489 nand3_x0
xsubckt_585_nand3_x0 0 1 170 2021 184 177 nand3_x0
xsubckt_1480_and21nor_x0 0 1 1116 468 595 681 and21nor_x0
xfeed_7499 0 1 decap_w0
xfeed_7498 0 1 decap_w0
xfeed_7497 0 1 decap_w0
xfeed_7496 0 1 decap_w0
xfeed_7495 0 1 decap_w0
xfeed_7494 0 1 decap_w0
xfeed_7493 0 1 decap_w0
xfeed_7492 0 1 decap_w0
xfeed_7491 0 1 decap_w0
xfeed_7490 0 1 tie
xfeed_6969 0 1 decap_w0
xfeed_6968 0 1 decap_w0
xfeed_6967 0 1 decap_w0
xfeed_6966 0 1 decap_w0
xfeed_6965 0 1 decap_w0
xfeed_6964 0 1 decap_w0
xfeed_6963 0 1 decap_w0
xfeed_6962 0 1 decap_w0
xfeed_6961 0 1 decap_w0
xfeed_6960 0 1 decap_w0
xfeed_3189 0 1 decap_w0
xfeed_3188 0 1 decap_w0
xfeed_3187 0 1 decap_w0
xfeed_3186 0 1 decap_w0
xfeed_3185 0 1 decap_w0
xfeed_3184 0 1 decap_w0
xfeed_3183 0 1 decap_w0
xfeed_3182 0 1 decap_w0
xfeed_3181 0 1 decap_w0
xfeed_3180 0 1 decap_w0
xfeed_2659 0 1 decap_w0
xfeed_2658 0 1 decap_w0
xfeed_2657 0 1 decap_w0
xfeed_2656 0 1 decap_w0
xfeed_2655 0 1 decap_w0
xfeed_2654 0 1 decap_w0
xfeed_2653 0 1 decap_w0
xfeed_2652 0 1 decap_w0
xfeed_2651 0 1 decap_w0
xfeed_2650 0 1 decap_w0
xfeed_639 0 1 decap_w0
xfeed_638 0 1 decap_w0
xfeed_637 0 1 decap_w0
xfeed_636 0 1 decap_w0
xfeed_635 0 1 decap_w0
xfeed_634 0 1 decap_w0
xfeed_633 0 1 decap_w0
xfeed_632 0 1 decap_w0
xfeed_631 0 1 decap_w0
xfeed_630 0 1 decap_w0
xsubckt_400_and2_x1 0 1 349 351 350 and2_x1
xsubckt_566_and2_x1 0 1 189 663 191 and2_x1
xsubckt_1442_nand2_x0 0 1 1153 2046 479 nand2_x0
xfeed_10009 0 1 decap_w0
xfeed_10008 0 1 decap_w0
xfeed_10007 0 1 decap_w0
xfeed_10006 0 1 decap_w0
xfeed_10005 0 1 decap_w0
xfeed_10004 0 1 decap_w0
xfeed_10003 0 1 decap_w0
xfeed_10002 0 1 decap_w0
xfeed_10001 0 1 decap_w0
xfeed_10000 0 1 decap_w0
xfeed_8116 0 1 decap_w0
xfeed_8115 0 1 decap_w0
xfeed_8114 0 1 tie
xfeed_8113 0 1 decap_w0
xfeed_8112 0 1 decap_w0
xfeed_8111 0 1 decap_w0
xsubckt_1262_nand2_x0 0 1 1318 435 1320 nand2_x0
xsubckt_997_and2_x1 0 1 1532 524 1563 and2_x1
xfeed_8119 0 1 decap_w0
xfeed_8118 0 1 decap_w0
xfeed_8117 0 1 decap_w0
xfeed_6979 0 1 decap_w0
xfeed_6978 0 1 decap_w0
xfeed_6977 0 1 decap_w0
xfeed_6976 0 1 decap_w0
xfeed_6975 0 1 decap_w0
xfeed_6974 0 1 decap_w0
xfeed_6973 0 1 decap_w0
xfeed_6972 0 1 decap_w0
xfeed_6971 0 1 decap_w0
xfeed_6970 0 1 decap_w0
xfeed_3199 0 1 decap_w0
xfeed_3198 0 1 decap_w0
xfeed_3197 0 1 decap_w0
xfeed_3196 0 1 decap_w0
xfeed_3195 0 1 decap_w0
xfeed_3194 0 1 decap_w0
xfeed_3193 0 1 decap_w0
xfeed_3192 0 1 decap_w0
xfeed_3191 0 1 decap_w0
xfeed_3190 0 1 decap_w0
xfeed_2669 0 1 tie
xfeed_2668 0 1 decap_w0
xfeed_2667 0 1 decap_w0
xfeed_2666 0 1 decap_w0
xfeed_2665 0 1 decap_w0
xfeed_2664 0 1 decap_w0
xfeed_2663 0 1 decap_w0
xfeed_2662 0 1 decap_w0
xfeed_2661 0 1 decap_w0
xfeed_2660 0 1 decap_w0
xfeed_646 0 1 decap_w0
xfeed_645 0 1 decap_w0
xfeed_644 0 1 decap_w0
xfeed_643 0 1 decap_w0
xfeed_642 0 1 decap_w0
xfeed_641 0 1 decap_w0
xfeed_640 0 1 decap_w0
xsubckt_300_nand3_x0 0 1 448 616 556 451 nand3_x0
xsubckt_578_nand2_x0 0 1 177 181 178 nand2_x0
xsubckt_1777_and21nor_x0 0 1 817 971 820 819 and21nor_x0
xsubckt_1814_mux2_x1 0 1 1791 2048 800 773 mux2_x1
xsubckt_1930_dff_x1 0 1 2069 1818 67 dff_x1
xsubckt_1932_dff_x1 0 1 2067 1816 58 dff_x1
xsubckt_1934_dff_x1 0 1 1982 1814 51 dff_x1
xfeed_10019 0 1 decap_w0
xfeed_10018 0 1 decap_w0
xfeed_10017 0 1 decap_w0
xfeed_10016 0 1 decap_w0
xfeed_10015 0 1 decap_w0
xfeed_10014 0 1 decap_w0
xfeed_10013 0 1 decap_w0
xfeed_10012 0 1 decap_w0
xfeed_10011 0 1 decap_w0
xfeed_10010 0 1 decap_w0
xfeed_8123 0 1 decap_w0
xfeed_8122 0 1 decap_w0
xfeed_8121 0 1 decap_w0
xfeed_8120 0 1 decap_w0
xfeed_649 0 1 decap_w0
xfeed_648 0 1 decap_w0
xfeed_647 0 1 decap_w0
xsubckt_1122_or21nand_x0 0 1 1435 663 606 494 or21nand_x0
xsubckt_741_nand2_x0 0 1 1725 140 1766 nand2_x0
xsubckt_646_nor2_x0 0 1 113 1983 2074 nor2_x0
xsubckt_1511_nand3_x0 0 1 1085 1141 1087 1086 nand3_x0
xsubckt_1680_and21nor_x0 0 1 914 1070 925 1073 and21nor_x0
xsubckt_1890_dff_x1 0 1 1950 1849 77 dff_x1
xsubckt_1936_dff_x1 0 1 1974 1812 41 dff_x1
xsubckt_1938_dff_x1 0 1 1972 1810 41 dff_x1
xfeed_8129 0 1 tie
xfeed_8128 0 1 decap_w0
xfeed_8127 0 1 decap_w0
xfeed_8126 0 1 decap_w0
xfeed_8125 0 1 decap_w0
xfeed_8124 0 1 decap_w0
xfeed_6989 0 1 decap_w0
xfeed_6988 0 1 decap_w0
xfeed_6987 0 1 decap_w0
xfeed_6986 0 1 tie
xfeed_6985 0 1 decap_w0
xfeed_6984 0 1 decap_w0
xfeed_6983 0 1 decap_w0
xfeed_6982 0 1 tie
xfeed_6981 0 1 decap_w0
xfeed_6980 0 1 decap_w0
xfeed_2679 0 1 decap_w0
xfeed_2678 0 1 decap_w0
xfeed_2677 0 1 decap_w0
xfeed_2676 0 1 decap_w0
xfeed_2675 0 1 decap_w0
xfeed_2674 0 1 tie
xfeed_2673 0 1 decap_w0
xfeed_2672 0 1 decap_w0
xfeed_2671 0 1 decap_w0
xfeed_2670 0 1 decap_w0
xfeed_653 0 1 decap_w0
xfeed_652 0 1 decap_w0
xfeed_651 0 1 decap_w0
xfeed_650 0 1 decap_w0
xsubckt_1270_or3_x1 0 1 1310 774 1312 1311 or3_x1
xsubckt_1011_and4_x1 0 1 1518 1576 1550 1547 1542 and4_x1
xsubckt_827_nand3_x0 0 1 1649 2069 681 490 nand3_x0
xsubckt_294_nand4_x0 0 1 454 680 599 589 558 nand4_x0
xsubckt_251_or2_x1 0 1 500 684 501 or2_x1
xsubckt_1331_nand3_x0 0 1 1255 1273 1266 1257 nand3_x0
xsubckt_1476_and21nor_x0 0 1 1120 1122 1778 1782 and21nor_x0
xsubckt_1674_and2_x1 0 1 920 1101 921 and2_x1
xsubckt_1892_dff_x1 0 1 2011 2003 64 dff_x1
xsubckt_1894_dff_x1 0 1 2009 2001 64 dff_x1
xsubckt_1896_dff_x1 0 1 2007 1999 64 dff_x1
xfeed_13809 0 1 decap_w0
xfeed_13808 0 1 decap_w0
xfeed_13807 0 1 decap_w0
xfeed_13806 0 1 decap_w0
xfeed_13805 0 1 decap_w0
xfeed_13804 0 1 decap_w0
xfeed_13803 0 1 decap_w0
xfeed_13802 0 1 decap_w0
xfeed_13801 0 1 decap_w0
xfeed_13800 0 1 decap_w0
xfeed_10028 0 1 decap_w0
xfeed_10027 0 1 decap_w0
xfeed_10026 0 1 decap_w0
xfeed_10025 0 1 decap_w0
xfeed_10024 0 1 tie
xfeed_10023 0 1 decap_w0
xfeed_10022 0 1 decap_w0
xfeed_10021 0 1 decap_w0
xfeed_10020 0 1 decap_w0
xfeed_8130 0 1 decap_w0
xfeed_659 0 1 decap_w0
xfeed_658 0 1 decap_w0
xfeed_657 0 1 decap_w0
xfeed_656 0 1 decap_w0
xfeed_655 0 1 tie
xfeed_654 0 1 decap_w0
xsubckt_1075_and21nor_x0 0 1 1851 1477 1469 1480 and21nor_x0
xsubckt_647_nand3_x0 0 1 112 678 447 113 nand3_x0
xsubckt_471_nand2_x0 0 1 279 558 544 nand2_x0
xsubckt_1898_dff_x1 0 1 2005 1997 38 dff_x1
xfeed_8139 0 1 decap_w0
xfeed_8138 0 1 tie
xfeed_8137 0 1 decap_w0
xfeed_8136 0 1 decap_w0
xfeed_8135 0 1 decap_w0
xfeed_8134 0 1 decap_w0
xfeed_8132 0 1 decap_w0
xfeed_8131 0 1 decap_w0
xfeed_7609 0 1 decap_w0
xfeed_7608 0 1 decap_w0
xfeed_7607 0 1 decap_w0
xfeed_7606 0 1 decap_w0
xfeed_7605 0 1 decap_w0
xfeed_7604 0 1 decap_w0
xfeed_7603 0 1 decap_w0
xfeed_7602 0 1 decap_w0
xfeed_7601 0 1 decap_w0
xfeed_7600 0 1 decap_w0
xfeed_6999 0 1 decap_w0
xfeed_6998 0 1 decap_w0
xfeed_6997 0 1 decap_w0
xfeed_6996 0 1 decap_w0
xfeed_6995 0 1 decap_w0
xfeed_6994 0 1 decap_w0
xfeed_6993 0 1 decap_w0
xfeed_6992 0 1 decap_w0
xfeed_6991 0 1 decap_w0
xfeed_6990 0 1 decap_w0
xfeed_2689 0 1 decap_w0
xfeed_2688 0 1 decap_w0
xfeed_2687 0 1 decap_w0
xfeed_2686 0 1 decap_w0
xfeed_2685 0 1 decap_w0
xfeed_2684 0 1 decap_w0
xfeed_2683 0 1 decap_w0
xfeed_2682 0 1 decap_w0
xfeed_2681 0 1 decap_w0
xfeed_2680 0 1 decap_w0
xfeed_660 0 1 decap_w0
xsubckt_735_and2_x1 0 1 1730 2052 1748 and2_x1
xsubckt_1536_or2_x1 0 1 1058 690 1116 or2_x1
xfeed_13819 0 1 decap_w0
xfeed_13818 0 1 decap_w0
xfeed_13817 0 1 decap_w0
xfeed_13816 0 1 decap_w0
xfeed_13815 0 1 decap_w0
xfeed_13814 0 1 decap_w0
xfeed_13813 0 1 decap_w0
xfeed_13812 0 1 decap_w0
xfeed_13811 0 1 tie
xfeed_13810 0 1 decap_w0
xfeed_10039 0 1 decap_w0
xfeed_10038 0 1 decap_w0
xfeed_10037 0 1 decap_w0
xfeed_10036 0 1 tie
xfeed_10035 0 1 decap_w0
xfeed_10034 0 1 decap_w0
xfeed_10033 0 1 decap_w0
xfeed_10032 0 1 decap_w0
xfeed_10031 0 1 tie
xfeed_10030 0 1 decap_w0
xfeed_669 0 1 decap_w0
xfeed_668 0 1 decap_w0
xfeed_667 0 1 decap_w0
xfeed_666 0 1 decap_w0
xfeed_665 0 1 tie
xfeed_664 0 1 decap_w0
xfeed_663 0 1 decap_w0
xfeed_662 0 1 decap_w0
xfeed_661 0 1 decap_w0
xsubckt_113_nand2_x0 0 1 655 785 1999 nand2_x0
xsubckt_1414_nand2_x0 0 1 1179 774 1977 nand2_x0
xfeed_8149 0 1 decap_w0
xfeed_8148 0 1 decap_w0
xfeed_8147 0 1 decap_w0
xfeed_8146 0 1 decap_w0
xfeed_8145 0 1 tie
xfeed_8144 0 1 decap_w0
xfeed_8143 0 1 decap_w0
xfeed_8142 0 1 decap_w0
xfeed_8141 0 1 decap_w0
xfeed_8140 0 1 decap_w0
xfeed_7619 0 1 decap_w0
xfeed_7618 0 1 decap_w0
xfeed_7617 0 1 decap_w0
xfeed_7616 0 1 decap_w0
xfeed_7615 0 1 tie
xfeed_7614 0 1 tie
xfeed_7613 0 1 decap_w0
xfeed_7612 0 1 decap_w0
xfeed_7611 0 1 decap_w0
xfeed_7610 0 1 decap_w0
xfeed_3309 0 1 decap_w0
xfeed_3308 0 1 decap_w0
xfeed_3307 0 1 decap_w0
xfeed_3306 0 1 decap_w0
xfeed_3305 0 1 decap_w0
xfeed_3304 0 1 decap_w0
xfeed_3303 0 1 decap_w0
xfeed_3302 0 1 decap_w0
xfeed_3301 0 1 decap_w0
xfeed_3300 0 1 decap_w0
xfeed_2699 0 1 decap_w0
xfeed_2698 0 1 decap_w0
xfeed_2697 0 1 decap_w0
xfeed_2696 0 1 decap_w0
xfeed_2695 0 1 tie
xfeed_2694 0 1 decap_w0
xfeed_2693 0 1 decap_w0
xfeed_2692 0 1 decap_w0
xfeed_2691 0 1 tie
xfeed_2690 0 1 decap_w0
xsubckt_168_and3_x1 0 1 590 605 600 591 and3_x1
xsubckt_109_nand3_x0 0 1 663 679 674 670 nand3_x0
xsubckt_1324_nand2_x0 0 1 1262 774 1970 nand2_x0
xfeed_13829 0 1 decap_w0
xfeed_13828 0 1 decap_w0
xfeed_13827 0 1 decap_w0
xfeed_13826 0 1 decap_w0
xfeed_13825 0 1 decap_w0
xfeed_13824 0 1 decap_w0
xfeed_13823 0 1 decap_w0
xfeed_13822 0 1 decap_w0
xfeed_13821 0 1 decap_w0
xfeed_13820 0 1 decap_w0
xfeed_10049 0 1 decap_w0
xfeed_10048 0 1 decap_w0
xfeed_10047 0 1 decap_w0
xfeed_10046 0 1 tie
xfeed_10045 0 1 decap_w0
xfeed_10044 0 1 decap_w0
xfeed_10043 0 1 decap_w0
xfeed_10042 0 1 decap_w0
xfeed_10040 0 1 decap_w0
xfeed_679 0 1 decap_w0
xfeed_678 0 1 decap_w0
xfeed_677 0 1 decap_w0
xfeed_676 0 1 decap_w0
xfeed_675 0 1 decap_w0
xfeed_674 0 1 decap_w0
xfeed_673 0 1 decap_w0
xfeed_672 0 1 decap_w0
xfeed_671 0 1 decap_w0
xfeed_670 0 1 tie
xsubckt_197_nand3_x0 0 1 561 590 577 562 nand3_x0
xsubckt_1486_and2_x1 0 1 1110 1119 1112 and2_x1
xfeed_8159 0 1 decap_w0
xfeed_8158 0 1 decap_w0
xfeed_8157 0 1 decap_w0
xfeed_8156 0 1 decap_w0
xfeed_8155 0 1 decap_w0
xfeed_8154 0 1 decap_w0
xfeed_8153 0 1 decap_w0
xfeed_8152 0 1 tie
xfeed_8151 0 1 decap_w0
xfeed_8150 0 1 decap_w0
xfeed_7629 0 1 decap_w0
xfeed_7628 0 1 decap_w0
xfeed_7627 0 1 tie
xfeed_7626 0 1 decap_w0
xfeed_7625 0 1 decap_w0
xfeed_7624 0 1 decap_w0
xfeed_7623 0 1 decap_w0
xfeed_7622 0 1 decap_w0
xfeed_7621 0 1 decap_w0
xfeed_7620 0 1 decap_w0
xfeed_3319 0 1 tie
xfeed_3318 0 1 decap_w0
xfeed_3317 0 1 decap_w0
xfeed_3316 0 1 decap_w0
xfeed_3315 0 1 tie
xfeed_3314 0 1 decap_w0
xfeed_3313 0 1 decap_w0
xfeed_3312 0 1 decap_w0
xfeed_3311 0 1 decap_w0
xfeed_3310 0 1 decap_w0
xsubckt_1054_nand2_x0 0 1 1487 1503 1488 nand2_x0
xfeed_13839 0 1 tie
xfeed_13838 0 1 decap_w0
xfeed_13837 0 1 decap_w0
xfeed_13836 0 1 decap_w0
xfeed_13835 0 1 decap_w0
xfeed_13834 0 1 decap_w0
xfeed_13833 0 1 decap_w0
xfeed_13832 0 1 decap_w0
xfeed_13831 0 1 decap_w0
xfeed_13830 0 1 decap_w0
xfeed_10059 0 1 decap_w0
xfeed_10058 0 1 decap_w0
xfeed_10057 0 1 decap_w0
xfeed_10056 0 1 decap_w0
xfeed_10055 0 1 decap_w0
xfeed_10054 0 1 decap_w0
xfeed_10053 0 1 decap_w0
xfeed_10052 0 1 decap_w0
xfeed_10051 0 1 decap_w0
xfeed_10050 0 1 tie
xfeed_689 0 1 tie
xfeed_688 0 1 decap_w0
xfeed_687 0 1 decap_w0
xfeed_686 0 1 decap_w0
xfeed_685 0 1 decap_w0
xfeed_684 0 1 decap_w0
xfeed_683 0 1 decap_w0
xfeed_682 0 1 tie
xfeed_681 0 1 decap_w0
xfeed_680 0 1 decap_w0
xsubckt_180_nand3_x0 0 1 578 617 586 581 nand3_x0
xsubckt_101_inv_x0 0 1 1996 689 inv_x0
xsubckt_452_or21nand_x0 0 1 298 299 302 358 or21nand_x0
xsubckt_547_and2_x1 0 1 207 600 209 and2_x1
xsubckt_1394_and2_x1 0 1 1197 1203 1198 and2_x1
xfeed_8169 0 1 decap_w0
xfeed_8168 0 1 decap_w0
xfeed_8167 0 1 decap_w0
xfeed_8166 0 1 tie
xfeed_8165 0 1 decap_w0
xfeed_8164 0 1 decap_w0
xfeed_8163 0 1 decap_w0
xfeed_8162 0 1 decap_w0
xfeed_8161 0 1 decap_w0
xfeed_8160 0 1 decap_w0
xfeed_7639 0 1 decap_w0
xfeed_7638 0 1 decap_w0
xfeed_7637 0 1 decap_w0
xfeed_7636 0 1 decap_w0
xfeed_7635 0 1 decap_w0
xfeed_7634 0 1 tie
xfeed_7633 0 1 decap_w0
xfeed_7632 0 1 decap_w0
xfeed_7631 0 1 decap_w0
xfeed_7630 0 1 decap_w0
xfeed_3329 0 1 decap_w0
xfeed_3328 0 1 decap_w0
xfeed_3327 0 1 decap_w0
xfeed_3326 0 1 decap_w0
xfeed_3325 0 1 decap_w0
xfeed_3324 0 1 decap_w0
xfeed_3322 0 1 decap_w0
xfeed_3321 0 1 decap_w0
xfeed_3320 0 1 decap_w0
xsubckt_1127_xor2_x0 0 1 1430 2056 2057 xor2_x0
xsubckt_176_nand4_x0 0 1 582 681 599 589 584 nand4_x0
xsubckt_1318_or21nand_x0 0 1 1267 1268 1322 762 or21nand_x0
xsubckt_1391_nand3_x0 0 1 1200 2070 666 657 nand3_x0
xfeed_13849 0 1 decap_w0
xfeed_13848 0 1 decap_w0
xfeed_13847 0 1 decap_w0
xfeed_13846 0 1 decap_w0
xfeed_13845 0 1 decap_w0
xfeed_13844 0 1 decap_w0
xfeed_13843 0 1 decap_w0
xfeed_13842 0 1 decap_w0
xfeed_13841 0 1 decap_w0
xfeed_13840 0 1 decap_w0
xfeed_10069 0 1 decap_w0
xfeed_10068 0 1 decap_w0
xfeed_10067 0 1 decap_w0
xfeed_10066 0 1 decap_w0
xfeed_10065 0 1 decap_w0
xfeed_10064 0 1 tie
xfeed_10063 0 1 decap_w0
xfeed_10062 0 1 decap_w0
xfeed_10061 0 1 decap_w0
xfeed_10060 0 1 tie
xfeed_699 0 1 tie
xfeed_698 0 1 decap_w0
xfeed_697 0 1 decap_w0
xfeed_696 0 1 decap_w0
xfeed_695 0 1 decap_w0
xfeed_694 0 1 tie
xfeed_693 0 1 decap_w0
xfeed_692 0 1 decap_w0
xfeed_691 0 1 decap_w0
xfeed_690 0 1 decap_w0
xfeed_8179 0 1 decap_w0
xfeed_8178 0 1 decap_w0
xfeed_8177 0 1 decap_w0
xfeed_8176 0 1 decap_w0
xfeed_8175 0 1 decap_w0
xfeed_8174 0 1 decap_w0
xfeed_8173 0 1 decap_w0
xfeed_8172 0 1 decap_w0
xfeed_8171 0 1 decap_w0
xfeed_8170 0 1 decap_w0
xfeed_7649 0 1 decap_w0
xfeed_7648 0 1 tie
xfeed_7647 0 1 decap_w0
xfeed_7646 0 1 decap_w0
xfeed_7645 0 1 decap_w0
xfeed_7644 0 1 decap_w0
xfeed_7643 0 1 decap_w0
xfeed_7642 0 1 decap_w0
xfeed_7641 0 1 tie
xfeed_7640 0 1 decap_w0
xfeed_3339 0 1 decap_w0
xfeed_3338 0 1 decap_w0
xfeed_3337 0 1 decap_w0
xfeed_3336 0 1 decap_w0
xfeed_3335 0 1 decap_w0
xfeed_3334 0 1 decap_w0
xfeed_3333 0 1 decap_w0
xfeed_3332 0 1 decap_w0
xfeed_3331 0 1 decap_w0
xfeed_3330 0 1 decap_w0
xfeed_2809 0 1 decap_w0
xfeed_2808 0 1 decap_w0
xfeed_2807 0 1 decap_w0
xfeed_2806 0 1 decap_w0
xfeed_2804 0 1 decap_w0
xfeed_2803 0 1 decap_w0
xfeed_2802 0 1 decap_w0
xfeed_2801 0 1 decap_w0
xfeed_2800 0 1 decap_w0
xsubckt_1033_nand3_x0 0 1 1502 645 637 633 nand3_x0
xsubckt_104_nor2_x0 0 1 683 1925 1926 nor2_x0
xsubckt_349_nand3_x0 0 1 399 712 1926 405 nand3_x0
xfeed_13859 0 1 decap_w0
xfeed_13858 0 1 decap_w0
xfeed_13857 0 1 decap_w0
xfeed_13856 0 1 decap_w0
xfeed_13855 0 1 decap_w0
xfeed_13854 0 1 decap_w0
xfeed_13853 0 1 decap_w0
xfeed_13852 0 1 decap_w0
xfeed_13851 0 1 decap_w0
xfeed_13850 0 1 decap_w0
xfeed_10079 0 1 tie
xfeed_10078 0 1 decap_w0
xfeed_10077 0 1 decap_w0
xfeed_10076 0 1 decap_w0
xfeed_10075 0 1 decap_w0
xfeed_10074 0 1 decap_w0
xfeed_10073 0 1 decap_w0
xfeed_10071 0 1 decap_w0
xfeed_10070 0 1 decap_w0
xsubckt_934_mux2_x1 0 1 1883 2023 1586 1578 mux2_x1
xsubckt_259_nand3_x0 0 1 492 617 557 495 nand3_x0
xsubckt_105_or2_x1 0 1 676 1925 1926 or2_x1
xsubckt_1519_or3_x1 0 1 1077 208 1080 1079 or3_x1
xfeed_8189 0 1 decap_w0
xfeed_8188 0 1 decap_w0
xfeed_8187 0 1 tie
xfeed_8186 0 1 decap_w0
xfeed_8185 0 1 decap_w0
xfeed_8184 0 1 decap_w0
xfeed_8183 0 1 decap_w0
xfeed_8182 0 1 decap_w0
xfeed_8181 0 1 decap_w0
xfeed_8180 0 1 decap_w0
xfeed_7659 0 1 decap_w0
xfeed_7658 0 1 decap_w0
xfeed_7657 0 1 decap_w0
xfeed_7656 0 1 decap_w0
xfeed_7655 0 1 tie
xfeed_7654 0 1 decap_w0
xfeed_7653 0 1 decap_w0
xfeed_7652 0 1 decap_w0
xfeed_7651 0 1 decap_w0
xfeed_7650 0 1 decap_w0
xfeed_3349 0 1 decap_w0
xfeed_3348 0 1 decap_w0
xfeed_3347 0 1 decap_w0
xfeed_3346 0 1 decap_w0
xfeed_3345 0 1 decap_w0
xfeed_3344 0 1 decap_w0
xfeed_3343 0 1 decap_w0
xfeed_3342 0 1 decap_w0
xfeed_3341 0 1 decap_w0
xfeed_3340 0 1 decap_w0
xfeed_2819 0 1 decap_w0
xfeed_2818 0 1 decap_w0
xfeed_2817 0 1 decap_w0
xfeed_2816 0 1 decap_w0
xfeed_2815 0 1 decap_w0
xfeed_2814 0 1 decap_w0
xfeed_2813 0 1 tie
xfeed_2812 0 1 decap_w0
xfeed_2811 0 1 decap_w0
xfeed_2810 0 1 decap_w0
xsubckt_1206_nand2_x0 0 1 1358 712 405 nand2_x0
xsubckt_794_and2_x1 0 1 1678 1681 1679 and2_x1
xsubckt_245_and3_x1 0 1 506 712 1926 571 and3_x1
xsubckt_1340_or2_x1 0 1 1247 1252 1249 or2_x1
xfeed_13869 0 1 decap_w0
xfeed_13868 0 1 decap_w0
xfeed_13867 0 1 decap_w0
xfeed_13866 0 1 decap_w0
xfeed_13865 0 1 decap_w0
xfeed_13864 0 1 decap_w0
xfeed_13863 0 1 decap_w0
xfeed_13862 0 1 decap_w0
xfeed_13861 0 1 decap_w0
xfeed_13860 0 1 decap_w0
xfeed_10089 0 1 decap_w0
xfeed_10088 0 1 decap_w0
xfeed_10087 0 1 tie
xfeed_10086 0 1 decap_w0
xfeed_10085 0 1 decap_w0
xfeed_10084 0 1 decap_w0
xfeed_10083 0 1 decap_w0
xfeed_10082 0 1 decap_w0
xfeed_10081 0 1 decap_w0
xfeed_10080 0 1 decap_w0
xsubckt_1026_nand2_x0 0 1 1508 1964 1509 nand2_x0
xsubckt_752_or21nand_x0 0 1 1715 2062 1742 1740 or21nand_x0
xsubckt_21_inv_x0 0 1 761 2055 inv_x0
xsubckt_332_nand3_x0 0 1 416 686 617 418 nand3_x0
xsubckt_1348_or2_x1 0 1 1240 696 1323 or2_x1
xsubckt_1633_nand3_x0 0 1 961 1973 682 595 nand3_x0
xfeed_8199 0 1 decap_w0
xfeed_8198 0 1 decap_w0
xfeed_8197 0 1 decap_w0
xfeed_8196 0 1 decap_w0
xfeed_8195 0 1 decap_w0
xfeed_8194 0 1 decap_w0
xfeed_8193 0 1 decap_w0
xfeed_8192 0 1 decap_w0
xfeed_8191 0 1 decap_w0
xfeed_8190 0 1 decap_w0
xfeed_7669 0 1 decap_w0
xfeed_7668 0 1 decap_w0
xfeed_7667 0 1 decap_w0
xfeed_7666 0 1 tie
xfeed_7665 0 1 decap_w0
xfeed_7664 0 1 decap_w0
xfeed_7663 0 1 decap_w0
xfeed_7662 0 1 tie
xfeed_7661 0 1 decap_w0
xfeed_7660 0 1 decap_w0
xfeed_3359 0 1 decap_w0
xfeed_3358 0 1 tie
xfeed_3357 0 1 decap_w0
xfeed_3356 0 1 decap_w0
xfeed_3355 0 1 decap_w0
xfeed_3354 0 1 decap_w0
xfeed_3353 0 1 decap_w0
xfeed_3352 0 1 decap_w0
xfeed_3351 0 1 decap_w0
xfeed_3350 0 1 decap_w0
xfeed_2829 0 1 decap_w0
xfeed_2828 0 1 decap_w0
xfeed_2827 0 1 decap_w0
xfeed_2826 0 1 decap_w0
xfeed_2825 0 1 decap_w0
xfeed_2824 0 1 decap_w0
xfeed_2823 0 1 tie
xfeed_2822 0 1 decap_w0
xfeed_2821 0 1 decap_w0
xfeed_2820 0 1 decap_w0
xfeed_800 0 1 decap_w0
xsubckt_23_inv_x0 0 1 759 2046 inv_x0
xsubckt_25_inv_x0 0 1 757 1954 inv_x0
xsubckt_153_and3_x1 0 1 612 716 1924 670 and3_x1
xsubckt_328_nand4_x0 0 1 420 716 1924 1927 713 nand4_x0
xsubckt_1419_and4_x1 0 1 1174 435 1642 1176 1175 and4_x1
xfeed_13879 0 1 tie
xfeed_13876 0 1 tie
xfeed_13875 0 1 tie
xfeed_13874 0 1 tie
xfeed_13873 0 1 decap_w0
xfeed_13872 0 1 decap_w0
xfeed_13871 0 1 decap_w0
xfeed_13870 0 1 decap_w0
xfeed_10099 0 1 decap_w0
xfeed_10098 0 1 decap_w0
xfeed_10097 0 1 decap_w0
xfeed_10096 0 1 decap_w0
xfeed_10095 0 1 decap_w0
xfeed_10094 0 1 decap_w0
xfeed_10093 0 1 decap_w0
xfeed_10092 0 1 decap_w0
xfeed_10091 0 1 decap_w0
xfeed_10090 0 1 decap_w0
xfeed_809 0 1 decap_w0
xfeed_808 0 1 decap_w0
xfeed_807 0 1 decap_w0
xfeed_806 0 1 decap_w0
xfeed_805 0 1 tie
xfeed_804 0 1 decap_w0
xfeed_803 0 1 decap_w0
xfeed_802 0 1 decap_w0
xfeed_801 0 1 decap_w0
xsubckt_1172_nor3_x0 0 1 1390 1959 1940 1937 nor3_x0
xsubckt_683_nand2_x0 0 1 1780 2030 175 nand2_x0
xsubckt_238_nand4_x0 0 1 513 687 616 585 581 nand4_x0
xsubckt_27_inv_x0 0 1 755 1938 inv_x0
xsubckt_29_inv_x0 0 1 753 1974 inv_x0
xsubckt_147_or21nand_x0 0 1 621 661 646 639 or21nand_x0
xsubckt_1363_nand3_x0 0 1 1226 2072 666 657 nand3_x0
xsubckt_1718_or21nand_x0 0 1 876 877 1118 769 or21nand_x0
xsubckt_1806_nand2_x0 0 1 1796 792 790 nand2_x0
xfeed_7679 0 1 decap_w0
xfeed_7678 0 1 tie
xfeed_7677 0 1 decap_w0
xfeed_7676 0 1 decap_w0
xfeed_7675 0 1 decap_w0
xfeed_7674 0 1 decap_w0
xfeed_7673 0 1 decap_w0
xfeed_7672 0 1 decap_w0
xfeed_7671 0 1 decap_w0
xfeed_7670 0 1 decap_w0
xfeed_3369 0 1 decap_w0
xfeed_3368 0 1 decap_w0
xfeed_3367 0 1 decap_w0
xfeed_3366 0 1 decap_w0
xfeed_3365 0 1 decap_w0
xfeed_3364 0 1 decap_w0
xfeed_3363 0 1 decap_w0
xfeed_3362 0 1 decap_w0
xfeed_3361 0 1 decap_w0
xfeed_3360 0 1 decap_w0
xfeed_2839 0 1 decap_w0
xfeed_2838 0 1 decap_w0
xfeed_2837 0 1 decap_w0
xfeed_2836 0 1 decap_w0
xfeed_2835 0 1 decap_w0
xfeed_2834 0 1 decap_w0
xfeed_2833 0 1 decap_w0
xfeed_2832 0 1 decap_w0
xfeed_2831 0 1 decap_w0
xfeed_2830 0 1 tie
xsubckt_679_nand3_x0 0 1 1784 2022 184 176 nand3_x0
xfeed_13889 0 1 tie
xfeed_13887 0 1 tie
xfeed_13886 0 1 tie
xfeed_13884 0 1 tie
xfeed_13883 0 1 tie
xfeed_13881 0 1 tie
xfeed_13880 0 1 tie
xfeed_819 0 1 decap_w0
xfeed_818 0 1 decap_w0
xfeed_817 0 1 decap_w0
xfeed_816 0 1 decap_w0
xfeed_815 0 1 decap_w0
xfeed_814 0 1 decap_w0
xfeed_813 0 1 decap_w0
xfeed_812 0 1 decap_w0
xfeed_811 0 1 decap_w0
xfeed_810 0 1 decap_w0
xsubckt_589_nand3_x0 0 1 166 1941 608 460 nand3_x0
xfeed_7689 0 1 decap_w0
xfeed_7688 0 1 decap_w0
xfeed_7687 0 1 decap_w0
xfeed_7686 0 1 decap_w0
xfeed_7685 0 1 tie
xfeed_7684 0 1 decap_w0
xfeed_7683 0 1 decap_w0
xfeed_7682 0 1 decap_w0
xfeed_7681 0 1 decap_w0
xfeed_7680 0 1 decap_w0
xfeed_3379 0 1 tie
xfeed_3378 0 1 decap_w0
xfeed_3377 0 1 decap_w0
xfeed_3376 0 1 decap_w0
xfeed_3375 0 1 tie
xfeed_3374 0 1 decap_w0
xfeed_3373 0 1 decap_w0
xfeed_3372 0 1 decap_w0
xfeed_3371 0 1 decap_w0
xfeed_3370 0 1 decap_w0
xfeed_2849 0 1 decap_w0
xfeed_2848 0 1 decap_w0
xfeed_2847 0 1 decap_w0
xfeed_2846 0 1 decap_w0
xfeed_2845 0 1 decap_w0
xfeed_2844 0 1 decap_w0
xfeed_2843 0 1 decap_w0
xfeed_2842 0 1 decap_w0
xfeed_2841 0 1 decap_w0
xfeed_2840 0 1 decap_w0
xsubckt_704_nor2_x0 0 1 1760 506 1761 nor2_x0
xsubckt_528_and2_x1 0 1 224 370 225 and2_x1
xsubckt_1589_mux2_x1 0 1 1005 1052 1007 1142 mux2_x1
xfeed_13898 0 1 tie
xfeed_13897 0 1 tie
xfeed_13896 0 1 tie
xfeed_13895 0 1 tie
xfeed_13894 0 1 tie
xfeed_13893 0 1 tie
xfeed_13892 0 1 tie
xfeed_13891 0 1 tie
xfeed_829 0 1 decap_w0
xfeed_828 0 1 decap_w0
xfeed_827 0 1 decap_w0
xfeed_826 0 1 decap_w0
xfeed_825 0 1 decap_w0
xfeed_824 0 1 decap_w0
xfeed_823 0 1 decap_w0
xfeed_822 0 1 decap_w0
xfeed_821 0 1 decap_w0
xfeed_820 0 1 decap_w0
xsubckt_897_and4_x1 0 1 1590 1962 1964 2055 2047 and4_x1
xsubckt_690_nor2_x0 0 1 1773 726 212 nor2_x0
xsubckt_488_and3_x1 0 1 262 510 336 263 and3_x1
xfeed_8309 0 1 decap_w0
xfeed_8308 0 1 decap_w0
xfeed_8307 0 1 decap_w0
xfeed_8306 0 1 decap_w0
xfeed_8305 0 1 decap_w0
xfeed_8303 0 1 decap_w0
xfeed_8302 0 1 decap_w0
xfeed_8301 0 1 tie
xfeed_8300 0 1 decap_w0
xfeed_7699 0 1 tie
xfeed_7698 0 1 decap_w0
xfeed_7697 0 1 decap_w0
xfeed_7696 0 1 decap_w0
xfeed_7695 0 1 decap_w0
xfeed_7694 0 1 decap_w0
xfeed_7693 0 1 decap_w0
xfeed_7692 0 1 tie
xfeed_7691 0 1 decap_w0
xfeed_7690 0 1 decap_w0
xfeed_3389 0 1 decap_w0
xfeed_3388 0 1 decap_w0
xfeed_3387 0 1 decap_w0
xfeed_3386 0 1 decap_w0
xfeed_3385 0 1 decap_w0
xfeed_3384 0 1 decap_w0
xfeed_3383 0 1 decap_w0
xfeed_3382 0 1 decap_w0
xfeed_3381 0 1 decap_w0
xfeed_3380 0 1 decap_w0
xfeed_2859 0 1 decap_w0
xfeed_2858 0 1 decap_w0
xfeed_2857 0 1 decap_w0
xfeed_2856 0 1 decap_w0
xfeed_2855 0 1 decap_w0
xfeed_2854 0 1 decap_w0
xfeed_2853 0 1 decap_w0
xfeed_2852 0 1 decap_w0
xfeed_2851 0 1 decap_w0
xfeed_2850 0 1 decap_w0
xsubckt_1257_and3_x1 0 1 1323 605 493 1756 and3_x1
xsubckt_304_nand3_x0 0 1 444 686 617 447 nand3_x0
xsubckt_568_nand4_x0 0 1 187 1931 195 194 189 nand4_x0
xsubckt_1605_nand3_x0 0 1 989 1972 680 594 nand3_x0
xsubckt_1941_dff_x1 0 1 1969 1807 38 dff_x1
xfeed_10209 0 1 decap_w0
xfeed_10208 0 1 tie
xfeed_10207 0 1 decap_w0
xfeed_10206 0 1 decap_w0
xfeed_10205 0 1 decap_w0
xfeed_10204 0 1 decap_w0
xfeed_10203 0 1 tie
xfeed_10202 0 1 decap_w0
xfeed_10201 0 1 decap_w0
xfeed_10200 0 1 decap_w0
xfeed_839 0 1 decap_w0
xfeed_838 0 1 decap_w0
xfeed_837 0 1 decap_w0
xfeed_836 0 1 decap_w0
xfeed_835 0 1 decap_w0
xfeed_834 0 1 decap_w0
xfeed_833 0 1 decap_w0
xfeed_832 0 1 decap_w0
xfeed_831 0 1 decap_w0
xfeed_830 0 1 decap_w0
xsubckt_1500_and4_x1 0 1 1096 1996 1128 1098 1097 and4_x1
xsubckt_1943_dff_x1 0 1 1967 1805 38 dff_x1
xsubckt_1945_dff_x1 0 1 1979 1803 58 dff_x1
xsubckt_1947_dff_x1 0 1 1977 1801 58 dff_x1
xfeed_8319 0 1 decap_w0
xfeed_8318 0 1 decap_w0
xfeed_8317 0 1 decap_w0
xfeed_8316 0 1 decap_w0
xfeed_8315 0 1 decap_w0
xfeed_8314 0 1 decap_w0
xfeed_8313 0 1 decap_w0
xfeed_8312 0 1 decap_w0
xfeed_8311 0 1 tie
xfeed_8310 0 1 decap_w0
xfeed_4009 0 1 decap_w0
xfeed_4008 0 1 decap_w0
xfeed_4007 0 1 decap_w0
xfeed_4006 0 1 decap_w0
xfeed_4005 0 1 decap_w0
xfeed_4004 0 1 decap_w0
xfeed_4003 0 1 decap_w0
xfeed_4002 0 1 decap_w0
xfeed_4001 0 1 decap_w0
xfeed_4000 0 1 decap_w0
xfeed_3399 0 1 decap_w0
xfeed_3398 0 1 decap_w0
xfeed_3397 0 1 decap_w0
xfeed_3396 0 1 decap_w0
xfeed_3395 0 1 decap_w0
xfeed_3394 0 1 decap_w0
xfeed_3393 0 1 decap_w0
xfeed_3392 0 1 decap_w0
xfeed_3391 0 1 decap_w0
xfeed_3390 0 1 decap_w0
xfeed_2869 0 1 decap_w0
xfeed_2868 0 1 tie
xfeed_2867 0 1 decap_w0
xfeed_2866 0 1 decap_w0
xfeed_2865 0 1 decap_w0
xfeed_2864 0 1 decap_w0
xfeed_2863 0 1 decap_w0
xfeed_2862 0 1 decap_w0
xfeed_2861 0 1 decap_w0
xfeed_2860 0 1 decap_w0
xsubckt_1279_and2_x1 0 1 1302 1311 1303 and2_x1
xsubckt_1216_or21nand_x0 0 1 1348 451 610 617 or21nand_x0
xsubckt_915_mux2_x1 0 1 1900 1593 2040 1580 mux2_x1
xsubckt_745_nand2_x0 0 1 1721 2001 1746 nand2_x0
xsubckt_655_nand2_x0 0 1 2078 115 105 nand2_x0
xsubckt_1636_and2_x1 0 1 958 961 959 and2_x1
xsubckt_1949_dff_x1 0 1 1975 1799 58 dff_x1
xfeed_10219 0 1 decap_w0
xfeed_10218 0 1 decap_w0
xfeed_10217 0 1 decap_w0
xfeed_10216 0 1 decap_w0
xfeed_10215 0 1 decap_w0
xfeed_10214 0 1 decap_w0
xfeed_10213 0 1 decap_w0
xfeed_10212 0 1 decap_w0
xfeed_10211 0 1 decap_w0
xfeed_10210 0 1 decap_w0
xfeed_849 0 1 decap_w0
xfeed_848 0 1 decap_w0
xfeed_847 0 1 decap_w0
xfeed_846 0 1 decap_w0
xfeed_845 0 1 decap_w0
xfeed_844 0 1 decap_w0
xfeed_843 0 1 decap_w0
xfeed_842 0 1 decap_w0
xfeed_841 0 1 decap_w0
xfeed_840 0 1 decap_w0
xsubckt_989_mux2_x1 0 1 1867 1539 1945 1576 mux2_x1
xsubckt_1522_and3_x1 0 1 1074 1125 1085 1076 and3_x1
xfeed_8329 0 1 decap_w0
xfeed_8328 0 1 decap_w0
xfeed_8327 0 1 decap_w0
xfeed_8326 0 1 decap_w0
xfeed_8325 0 1 decap_w0
xfeed_8324 0 1 decap_w0
xfeed_8323 0 1 tie
xfeed_8322 0 1 decap_w0
xfeed_8321 0 1 decap_w0
xfeed_8320 0 1 decap_w0
xfeed_4019 0 1 decap_w0
xfeed_4018 0 1 decap_w0
xfeed_4017 0 1 decap_w0
xfeed_4016 0 1 decap_w0
xfeed_4015 0 1 decap_w0
xfeed_4014 0 1 decap_w0
xfeed_4013 0 1 decap_w0
xfeed_4012 0 1 decap_w0
xfeed_4011 0 1 decap_w0
xfeed_4010 0 1 decap_w0
xfeed_2879 0 1 decap_w0
xfeed_2878 0 1 decap_w0
xfeed_2877 0 1 decap_w0
xfeed_2876 0 1 decap_w0
xfeed_2875 0 1 decap_w0
xfeed_2874 0 1 decap_w0
xfeed_2873 0 1 decap_w0
xfeed_2872 0 1 tie
xfeed_2871 0 1 decap_w0
xfeed_2870 0 1 decap_w0
xsubckt_1235_mux2_x1 0 1 1826 2096 2061 1334 mux2_x1
xsubckt_1187_and2_x1 0 1 1377 551 1379 and2_x1
xsubckt_812_and21nor_x0 0 1 1662 745 600 1745 and21nor_x0
xsubckt_252_and2_x1 0 1 499 679 571 and2_x1
xsubckt_385_nand2_x0 0 1 364 687 468 nand2_x0
xfeed_10229 0 1 decap_w0
xfeed_10228 0 1 decap_w0
xfeed_10227 0 1 decap_w0
xfeed_10225 0 1 decap_w0
xfeed_10224 0 1 decap_w0
xfeed_10223 0 1 decap_w0
xfeed_10222 0 1 decap_w0
xfeed_10221 0 1 decap_w0
xfeed_10220 0 1 decap_w0
xfeed_859 0 1 decap_w0
xfeed_858 0 1 decap_w0
xfeed_857 0 1 decap_w0
xfeed_856 0 1 decap_w0
xfeed_855 0 1 decap_w0
xfeed_854 0 1 decap_w0
xfeed_853 0 1 decap_w0
xfeed_852 0 1 decap_w0
xfeed_851 0 1 decap_w0
xfeed_850 0 1 decap_w0
xsubckt_988_nand4_x0 0 1 1539 525 1549 1546 1543 nand4_x0
xsubckt_951_or21nand_x0 0 1 1875 1571 1569 1573 or21nand_x0
xsubckt_724_nand3_x0 0 1 1740 592 574 478 nand3_x0
xsubckt_281_nand4_x0 0 1 467 1925 711 599 589 nand4_x0
xsubckt_411_and21nor_x0 0 1 338 339 343 344 and21nor_x0
xsubckt_1508_nand2_x0 0 1 1088 1101 1089 nand2_x0
xsubckt_1620_or21nand_x0 0 1 974 975 976 1075 or21nand_x0
xfeed_8339 0 1 decap_w0
xfeed_8337 0 1 decap_w0
xfeed_8336 0 1 decap_w0
xfeed_8335 0 1 tie
xfeed_8334 0 1 decap_w0
xfeed_8333 0 1 decap_w0
xfeed_8332 0 1 decap_w0
xfeed_8331 0 1 decap_w0
xfeed_8330 0 1 decap_w0
xfeed_7809 0 1 decap_w0
xfeed_7808 0 1 decap_w0
xfeed_7807 0 1 decap_w0
xfeed_7806 0 1 decap_w0
xfeed_7804 0 1 decap_w0
xfeed_7803 0 1 decap_w0
xfeed_7802 0 1 decap_w0
xfeed_7801 0 1 decap_w0
xfeed_7800 0 1 decap_w0
xfeed_4029 0 1 decap_w0
xfeed_4028 0 1 decap_w0
xfeed_4027 0 1 decap_w0
xfeed_4026 0 1 decap_w0
xfeed_4025 0 1 decap_w0
xfeed_4024 0 1 decap_w0
xfeed_4023 0 1 decap_w0
xfeed_4022 0 1 decap_w0
xfeed_4021 0 1 decap_w0
xfeed_4020 0 1 decap_w0
xfeed_2889 0 1 decap_w0
xfeed_2888 0 1 decap_w0
xfeed_2887 0 1 decap_w0
xfeed_2886 0 1 decap_w0
xfeed_2885 0 1 decap_w0
xfeed_2884 0 1 decap_w0
xfeed_2883 0 1 decap_w0
xfeed_2882 0 1 decap_w0
xfeed_2881 0 1 decap_w0
xfeed_2880 0 1 decap_w0
xsubckt_1072_and21nor_x0 0 1 1471 1472 1474 1555 and21nor_x0
xsubckt_160_and2_x1 0 1 601 610 603 and2_x1
xsubckt_608_and21nor_x0 0 1 148 754 449 410 and21nor_x0
xfeed_10239 0 1 decap_w0
xfeed_10238 0 1 decap_w0
xfeed_10237 0 1 decap_w0
xfeed_10236 0 1 decap_w0
xfeed_10235 0 1 decap_w0
xfeed_10234 0 1 tie
xfeed_10233 0 1 decap_w0
xfeed_10232 0 1 decap_w0
xfeed_10231 0 1 decap_w0
xfeed_10230 0 1 decap_w0
xfeed_869 0 1 decap_w0
xfeed_868 0 1 decap_w0
xfeed_867 0 1 decap_w0
xfeed_866 0 1 decap_w0
xfeed_865 0 1 decap_w0
xfeed_864 0 1 decap_w0
xfeed_863 0 1 decap_w0
xfeed_862 0 1 decap_w0
xfeed_861 0 1 decap_w0
xfeed_860 0 1 decap_w0
xsubckt_1269_and21nor_x0 0 1 1311 1324 1315 1313 and21nor_x0
xsubckt_650_or21nand_x0 0 1 109 608 603 460 or21nand_x0
xsubckt_110_and21nor_x0 0 1 662 1983 2074 786 and21nor_x0
xfeed_8349 0 1 tie
xfeed_8348 0 1 decap_w0
xfeed_8347 0 1 decap_w0
xfeed_8346 0 1 decap_w0
xfeed_8345 0 1 decap_w0
xfeed_8344 0 1 decap_w0
xfeed_8343 0 1 decap_w0
xfeed_8341 0 1 decap_w0
xfeed_8340 0 1 decap_w0
xfeed_7819 0 1 decap_w0
xfeed_7818 0 1 decap_w0
xfeed_7817 0 1 decap_w0
xfeed_7816 0 1 decap_w0
xfeed_7815 0 1 decap_w0
xfeed_7814 0 1 decap_w0
xfeed_7813 0 1 decap_w0
xfeed_7812 0 1 decap_w0
xfeed_7811 0 1 decap_w0
xfeed_7810 0 1 decap_w0
xfeed_4039 0 1 decap_w0
xfeed_4038 0 1 decap_w0
xfeed_4037 0 1 decap_w0
xfeed_4036 0 1 tie
xfeed_4035 0 1 decap_w0
xfeed_4034 0 1 decap_w0
xfeed_4033 0 1 decap_w0
xfeed_4032 0 1 decap_w0
xfeed_4031 0 1 tie
xfeed_4030 0 1 decap_w0
xfeed_3509 0 1 decap_w0
xfeed_3508 0 1 decap_w0
xfeed_3507 0 1 decap_w0
xfeed_3506 0 1 decap_w0
xfeed_3505 0 1 decap_w0
xfeed_3504 0 1 decap_w0
xfeed_3503 0 1 decap_w0
xfeed_3502 0 1 tie
xfeed_3501 0 1 decap_w0
xfeed_3500 0 1 decap_w0
xfeed_2899 0 1 decap_w0
xfeed_2898 0 1 decap_w0
xfeed_2897 0 1 decap_w0
xfeed_2896 0 1 decap_w0
xfeed_2895 0 1 tie
xfeed_2894 0 1 decap_w0
xfeed_2892 0 1 decap_w0
xfeed_2891 0 1 decap_w0
xfeed_2890 0 1 decap_w0
xsubckt_1401_nand2_x0 0 1 1191 1978 1316 nand2_x0
xfeed_10249 0 1 tie
xfeed_10248 0 1 decap_w0
xfeed_10247 0 1 decap_w0
xfeed_10246 0 1 decap_w0
xfeed_10245 0 1 decap_w0
xfeed_10244 0 1 decap_w0
xfeed_10243 0 1 decap_w0
xfeed_10242 0 1 decap_w0
xfeed_10241 0 1 decap_w0
xfeed_10240 0 1 decap_w0
xfeed_879 0 1 decap_w0
xfeed_878 0 1 decap_w0
xfeed_877 0 1 decap_w0
xfeed_876 0 1 decap_w0
xfeed_875 0 1 tie
xfeed_874 0 1 decap_w0
xfeed_873 0 1 decap_w0
xfeed_872 0 1 decap_w0
xfeed_871 0 1 decap_w0
xfeed_870 0 1 decap_w0
xsubckt_808_and21nor_x0 0 1 1666 694 1755 1754 and21nor_x0
xsubckt_447_and4_x1 0 1 303 660 656 655 624 and4_x1
xsubckt_627_nand2_x0 0 1 131 2034 175 nand2_x0
xfeed_8359 0 1 decap_w0
xfeed_8358 0 1 decap_w0
xfeed_8357 0 1 decap_w0
xfeed_8356 0 1 decap_w0
xfeed_8354 0 1 decap_w0
xfeed_8353 0 1 decap_w0
xfeed_8352 0 1 decap_w0
xfeed_8351 0 1 decap_w0
xfeed_8350 0 1 decap_w0
xfeed_7829 0 1 decap_w0
xfeed_7828 0 1 decap_w0
xfeed_7827 0 1 decap_w0
xfeed_7826 0 1 decap_w0
xfeed_7825 0 1 decap_w0
xfeed_7824 0 1 decap_w0
xfeed_7823 0 1 decap_w0
xfeed_7822 0 1 decap_w0
xfeed_7821 0 1 decap_w0
xfeed_7820 0 1 decap_w0
xfeed_4049 0 1 decap_w0
xfeed_4048 0 1 decap_w0
xfeed_4047 0 1 decap_w0
xfeed_4046 0 1 decap_w0
xfeed_4045 0 1 decap_w0
xfeed_4044 0 1 decap_w0
xfeed_4043 0 1 decap_w0
xfeed_4042 0 1 decap_w0
xfeed_4041 0 1 decap_w0
xfeed_4040 0 1 decap_w0
xfeed_3519 0 1 decap_w0
xfeed_3518 0 1 decap_w0
xfeed_3517 0 1 decap_w0
xfeed_3516 0 1 decap_w0
xfeed_3514 0 1 decap_w0
xfeed_3513 0 1 decap_w0
xfeed_3512 0 1 decap_w0
xfeed_3511 0 1 decap_w0
xfeed_3510 0 1 decap_w0
xsubckt_947_or21nand_x0 0 1 1876 1572 1573 295 or21nand_x0
xsubckt_805_or4_x1 0 1 1668 1673 1672 1671 1669 or4_x1
xsubckt_421_and2_x1 0 1 328 330 329 and2_x1
xsubckt_1713_and2_x1 0 1 881 884 882 and2_x1
xfeed_10259 0 1 decap_w0
xfeed_10258 0 1 decap_w0
xfeed_10257 0 1 decap_w0
xfeed_10256 0 1 tie
xfeed_10255 0 1 decap_w0
xfeed_10254 0 1 decap_w0
xfeed_10253 0 1 decap_w0
xfeed_10252 0 1 decap_w0
xfeed_10251 0 1 decap_w0
xfeed_10250 0 1 decap_w0
xfeed_889 0 1 decap_w0
xfeed_888 0 1 decap_w0
xfeed_887 0 1 decap_w0
xfeed_886 0 1 decap_w0
xfeed_885 0 1 decap_w0
xfeed_884 0 1 decap_w0
xfeed_883 0 1 decap_w0
xfeed_882 0 1 decap_w0
xfeed_881 0 1 decap_w0
xfeed_880 0 1 decap_w0
xsubckt_495_and2_x1 0 1 256 258 257 and2_x1
xsubckt_1773_and21nor_x0 0 1 821 822 825 833 and21nor_x0
xfeed_8369 0 1 decap_w0
xfeed_8368 0 1 decap_w0
xfeed_8367 0 1 decap_w0
xfeed_8366 0 1 decap_w0
xfeed_8365 0 1 decap_w0
xfeed_8364 0 1 decap_w0
xfeed_8363 0 1 decap_w0
xfeed_8362 0 1 decap_w0
xfeed_8361 0 1 decap_w0
xfeed_8360 0 1 tie
xfeed_7839 0 1 tie
xfeed_7838 0 1 decap_w0
xfeed_7837 0 1 decap_w0
xfeed_7836 0 1 decap_w0
xfeed_7835 0 1 decap_w0
xfeed_7834 0 1 decap_w0
xfeed_7833 0 1 decap_w0
xfeed_7832 0 1 tie
xfeed_7831 0 1 decap_w0
xfeed_7830 0 1 decap_w0
xfeed_4059 0 1 decap_w0
xfeed_4058 0 1 decap_w0
xfeed_4057 0 1 decap_w0
xfeed_4056 0 1 decap_w0
xfeed_4055 0 1 decap_w0
xfeed_4054 0 1 decap_w0
xfeed_4053 0 1 decap_w0
xfeed_4052 0 1 decap_w0
xfeed_4051 0 1 decap_w0
xfeed_4050 0 1 decap_w0
xfeed_3529 0 1 decap_w0
xfeed_3528 0 1 decap_w0
xfeed_3527 0 1 decap_w0
xfeed_3526 0 1 decap_w0
xfeed_3525 0 1 decap_w0
xfeed_3524 0 1 decap_w0
xfeed_3523 0 1 decap_w0
xfeed_3522 0 1 tie
xfeed_3521 0 1 decap_w0
xfeed_3520 0 1 decap_w0
xsubckt_826_and3_x1 0 1 1650 2069 681 490 and3_x1
xsubckt_417_and2_x1 0 1 332 335 333 and2_x1
xfeed_10269 0 1 decap_w0
xfeed_10268 0 1 decap_w0
xfeed_10267 0 1 decap_w0
xfeed_10266 0 1 decap_w0
xfeed_10265 0 1 decap_w0
xfeed_10263 0 1 decap_w0
xfeed_10262 0 1 decap_w0
xfeed_10261 0 1 tie
xfeed_10260 0 1 decap_w0
xfeed_899 0 1 tie
xfeed_898 0 1 decap_w0
xfeed_897 0 1 decap_w0
xfeed_896 0 1 decap_w0
xfeed_895 0 1 decap_w0
xfeed_894 0 1 tie
xfeed_893 0 1 decap_w0
xfeed_892 0 1 decap_w0
xfeed_891 0 1 decap_w0
xfeed_890 0 1 tie
xsubckt_377_and3_x1 0 1 372 617 603 557 and3_x1
xfeed_8379 0 1 decap_w0
xfeed_8378 0 1 decap_w0
xfeed_8377 0 1 decap_w0
xfeed_8376 0 1 decap_w0
xfeed_8375 0 1 decap_w0
xfeed_8374 0 1 decap_w0
xfeed_8373 0 1 decap_w0
xfeed_8372 0 1 decap_w0
xfeed_8371 0 1 decap_w0
xfeed_8370 0 1 decap_w0
xfeed_7849 0 1 decap_w0
xfeed_7848 0 1 decap_w0
xfeed_7847 0 1 decap_w0
xfeed_7845 0 1 decap_w0
xfeed_7844 0 1 decap_w0
xfeed_7843 0 1 decap_w0
xfeed_7842 0 1 decap_w0
xfeed_7841 0 1 decap_w0
xfeed_7840 0 1 decap_w0
xfeed_4069 0 1 tie
xfeed_4068 0 1 decap_w0
xfeed_4067 0 1 decap_w0
xfeed_4066 0 1 decap_w0
xfeed_4065 0 1 decap_w0
xfeed_4064 0 1 decap_w0
xfeed_4063 0 1 decap_w0
xfeed_4062 0 1 tie
xfeed_4061 0 1 decap_w0
xfeed_4060 0 1 decap_w0
xfeed_3539 0 1 decap_w0
xfeed_3538 0 1 decap_w0
xfeed_3537 0 1 decap_w0
xfeed_3536 0 1 decap_w0
xfeed_3535 0 1 decap_w0
xfeed_3534 0 1 decap_w0
xfeed_3533 0 1 decap_w0
xfeed_3532 0 1 decap_w0
xfeed_3531 0 1 decap_w0
xfeed_3530 0 1 decap_w0
xsubckt_854_or2_x1 0 1 2099 1632 1626 or2_x1
xsubckt_734_and3_x1 0 1 1731 1981 1749 1739 and3_x1
xsubckt_1388_nand2_x0 0 1 1203 1979 1316 nand2_x0
xsubckt_1641_nand2_x0 0 1 953 955 954 nand2_x0
xfeed_10279 0 1 decap_w0
xfeed_10278 0 1 decap_w0
xfeed_10277 0 1 decap_w0
xfeed_10276 0 1 decap_w0
xfeed_10275 0 1 decap_w0
xfeed_10274 0 1 tie
xfeed_10273 0 1 decap_w0
xfeed_10272 0 1 decap_w0
xfeed_10271 0 1 decap_w0
xfeed_10270 0 1 decap_w0
xsubckt_957_nand2_x0 0 1 1564 1958 1575 nand2_x0
xsubckt_616_and4_x1 0 1 141 145 144 143 142 and4_x1
xfeed_8389 0 1 decap_w0
xfeed_8388 0 1 tie
xfeed_8387 0 1 decap_w0
xfeed_8385 0 1 decap_w0
xfeed_8384 0 1 decap_w0
xfeed_8383 0 1 tie
xfeed_8382 0 1 decap_w0
xfeed_8381 0 1 decap_w0
xfeed_8380 0 1 decap_w0
xfeed_7859 0 1 decap_w0
xfeed_7858 0 1 tie
xfeed_7857 0 1 decap_w0
xfeed_7856 0 1 decap_w0
xfeed_7855 0 1 decap_w0
xfeed_7854 0 1 decap_w0
xfeed_7853 0 1 decap_w0
xfeed_7852 0 1 decap_w0
xfeed_7851 0 1 decap_w0
xfeed_7850 0 1 decap_w0
xfeed_4079 0 1 decap_w0
xfeed_4078 0 1 decap_w0
xfeed_4077 0 1 decap_w0
xfeed_4076 0 1 decap_w0
xfeed_4075 0 1 decap_w0
xfeed_4074 0 1 tie
xfeed_4073 0 1 decap_w0
xfeed_4072 0 1 decap_w0
xfeed_4071 0 1 decap_w0
xfeed_4070 0 1 decap_w0
xfeed_3549 0 1 decap_w0
xfeed_3548 0 1 decap_w0
xfeed_3547 0 1 decap_w0
xfeed_3546 0 1 decap_w0
xfeed_3545 0 1 decap_w0
xfeed_3544 0 1 decap_w0
xfeed_3543 0 1 decap_w0
xfeed_3542 0 1 decap_w0
xfeed_3541 0 1 decap_w0
xfeed_3540 0 1 decap_w0
xsubckt_246_nand3_x0 0 1 505 712 1926 571 nand3_x0
xsubckt_30_inv_x0 0 1 752 1973 inv_x0
xsubckt_32_inv_x0 0 1 750 1971 inv_x0
xsubckt_343_nor4_x0 0 1 405 1929 1924 1927 1928 nor4_x0
xsubckt_1371_nand2_x0 0 1 1218 1917 1221 nand2_x0
xsubckt_1461_nand2_x0 0 1 1135 779 1949 nand2_x0
xsubckt_1515_or21nand_x0 0 1 1081 1942 548 1744 or21nand_x0
xsubckt_1769_and21nor_x0 0 1 825 830 828 826 and21nor_x0
xfeed_10289 0 1 decap_w0
xfeed_10288 0 1 decap_w0
xfeed_10287 0 1 decap_w0
xfeed_10285 0 1 decap_w0
xfeed_10284 0 1 decap_w0
xfeed_10283 0 1 decap_w0
xfeed_10282 0 1 decap_w0
xfeed_10281 0 1 decap_w0
xfeed_10280 0 1 decap_w0
xsubckt_878_mux2_x1 0 1 1605 1606 2001 445 mux2_x1
xsubckt_664_and2_x1 0 1 96 99 97 and2_x1
xsubckt_34_inv_x0 0 1 748 1969 inv_x0
xsubckt_36_inv_x0 0 1 746 2072 inv_x0
xsubckt_38_inv_x0 0 1 744 2070 inv_x0
xsubckt_1647_mux2_x1 0 1 947 992 949 1142 mux2_x1
xfeed_9009 0 1 decap_w0
xfeed_9008 0 1 decap_w0
xfeed_9007 0 1 decap_w0
xfeed_9006 0 1 decap_w0
xfeed_9005 0 1 tie
xfeed_9004 0 1 decap_w0
xfeed_9003 0 1 decap_w0
xfeed_9002 0 1 decap_w0
xfeed_9001 0 1 decap_w0
xfeed_9000 0 1 decap_w0
xfeed_8399 0 1 decap_w0
xfeed_8398 0 1 decap_w0
xfeed_8397 0 1 decap_w0
xfeed_8396 0 1 decap_w0
xfeed_8395 0 1 decap_w0
xfeed_8394 0 1 decap_w0
xfeed_8393 0 1 decap_w0
xfeed_8392 0 1 decap_w0
xfeed_8391 0 1 decap_w0
xfeed_8390 0 1 decap_w0
xfeed_7869 0 1 decap_w0
xfeed_7868 0 1 decap_w0
xfeed_7867 0 1 decap_w0
xfeed_7866 0 1 decap_w0
xfeed_7865 0 1 decap_w0
xfeed_7864 0 1 decap_w0
xfeed_7863 0 1 decap_w0
xfeed_7862 0 1 decap_w0
xfeed_7861 0 1 decap_w0
xfeed_7860 0 1 decap_w0
xfeed_4089 0 1 decap_w0
xfeed_4088 0 1 decap_w0
xfeed_4087 0 1 decap_w0
xfeed_4086 0 1 decap_w0
xfeed_4085 0 1 decap_w0
xfeed_4084 0 1 decap_w0
xfeed_4083 0 1 decap_w0
xfeed_4082 0 1 decap_w0
xfeed_4081 0 1 decap_w0
xfeed_4080 0 1 decap_w0
xfeed_3558 0 1 tie
xfeed_3557 0 1 decap_w0
xfeed_3556 0 1 decap_w0
xfeed_3555 0 1 decap_w0
xfeed_3554 0 1 decap_w0
xfeed_3553 0 1 decap_w0
xfeed_3551 0 1 decap_w0
xfeed_3550 0 1 decap_w0
xfeed_10299 0 1 decap_w0
xfeed_10298 0 1 decap_w0
xfeed_10297 0 1 decap_w0
xfeed_10296 0 1 decap_w0
xfeed_10295 0 1 decap_w0
xfeed_10294 0 1 decap_w0
xfeed_10293 0 1 decap_w0
xfeed_10292 0 1 tie
xfeed_10291 0 1 decap_w0
xfeed_10290 0 1 decap_w0
xsubckt_1429_and2_x1 0 1 1165 1976 1316 and2_x1
xsubckt_1530_nand3_x0 0 1 1063 1099 1095 1070 nand3_x0
xsubckt_1555_mux2_x1 0 1 1039 1040 1045 1052 mux2_x1
xfeed_9019 0 1 decap_w0
xfeed_9018 0 1 decap_w0
xfeed_9015 0 1 decap_w0
xfeed_9014 0 1 decap_w0
xfeed_9013 0 1 decap_w0
xfeed_9012 0 1 decap_w0
xfeed_9011 0 1 decap_w0
xfeed_9010 0 1 tie
xfeed_7879 0 1 decap_w0
xfeed_7878 0 1 decap_w0
xfeed_7877 0 1 decap_w0
xfeed_7876 0 1 decap_w0
xfeed_7875 0 1 decap_w0
xfeed_7874 0 1 decap_w0
xfeed_7873 0 1 decap_w0
xfeed_7872 0 1 decap_w0
xfeed_7871 0 1 decap_w0
xfeed_7870 0 1 decap_w0
xfeed_4099 0 1 decap_w0
xfeed_4098 0 1 decap_w0
xfeed_4097 0 1 decap_w0
xfeed_4096 0 1 decap_w0
xfeed_4095 0 1 decap_w0
xfeed_4094 0 1 decap_w0
xfeed_4093 0 1 decap_w0
xfeed_4092 0 1 decap_w0
xfeed_4091 0 1 decap_w0
xfeed_4090 0 1 decap_w0
xfeed_3569 0 1 decap_w0
xfeed_3568 0 1 tie
xfeed_3567 0 1 decap_w0
xfeed_3566 0 1 decap_w0
xfeed_3565 0 1 decap_w0
xfeed_3564 0 1 decap_w0
xfeed_3563 0 1 decap_w0
xfeed_3562 0 1 decap_w0
xfeed_3561 0 1 decap_w0
xfeed_3560 0 1 decap_w0
xsubckt_670_nand2_x0 0 1 91 2039 172 nand2_x0
xsubckt_1341_and2_x1 0 1 1246 1255 1248 and2_x1
xsubckt_1350_nand3_x0 0 1 1238 2073 666 657 nand3_x0
xsubckt_1223_and3_x1 0 1 1341 462 438 284 and3_x1
xsubckt_340_and4_x1 0 1 408 1927 713 682 674 and4_x1
xsubckt_490_nand2_x0 0 1 261 535 298 nand2_x0
xsubckt_1337_and2_x1 0 1 1250 435 1251 and2_x1
xsubckt_1703_nand2_x0 0 1 891 1101 893 nand2_x0
xfeed_9029 0 1 tie
xfeed_9028 0 1 decap_w0
xfeed_9027 0 1 decap_w0
xfeed_9026 0 1 decap_w0
xfeed_9025 0 1 decap_w0
xfeed_9024 0 1 decap_w0
xfeed_9023 0 1 decap_w0
xfeed_9022 0 1 tie
xfeed_9021 0 1 decap_w0
xfeed_9020 0 1 decap_w0
xfeed_7889 0 1 decap_w0
xfeed_7888 0 1 decap_w0
xfeed_7887 0 1 decap_w0
xfeed_7886 0 1 tie
xfeed_7885 0 1 decap_w0
xfeed_7884 0 1 decap_w0
xfeed_7883 0 1 decap_w0
xfeed_7882 0 1 decap_w0
xfeed_7881 0 1 decap_w0
xfeed_7880 0 1 decap_w0
xfeed_3579 0 1 decap_w0
xfeed_3578 0 1 decap_w0
xfeed_3577 0 1 decap_w0
xfeed_3576 0 1 decap_w0
xfeed_3575 0 1 decap_w0
xfeed_3574 0 1 decap_w0
xfeed_3573 0 1 decap_w0
xfeed_3572 0 1 decap_w0
xfeed_3571 0 1 decap_w0
xfeed_3570 0 1 decap_w0
xsubckt_1080_nand3_x0 0 1 1464 643 313 1483 nand3_x0
xsubckt_222_nand2_x0 0 1 529 1986 1989 nand2_x0
xsubckt_1267_and21nor_x0 0 1 1313 1314 1321 2053 and21nor_x0
xsubckt_833_and2_x1 0 1 1644 2048 1740 and2_x1
xsubckt_807_and3_x1 0 1 1667 1980 1749 1739 and3_x1
xsubckt_132_nand2_x0 0 1 636 1986 1993 nand2_x0
xsubckt_362_and3_x1 0 1 387 616 556 447 and3_x1
xsubckt_1654_and3_x1 0 1 940 948 944 942 and3_x1
xsubckt_1816_mux2_x1 0 1 1789 2046 801 775 mux2_x1
xsubckt_1950_dff_x1 0 1 2056 1798 45 dff_x1
xsubckt_1952_dff_x1 0 1 2053 1796 45 dff_x1
xsubckt_1954_dff_x1 0 1 2051 1794 45 dff_x1
xfeed_9039 0 1 tie
xfeed_9038 0 1 decap_w0
xfeed_9037 0 1 decap_w0
xfeed_9036 0 1 decap_w0
xfeed_9035 0 1 decap_w0
xfeed_9034 0 1 decap_w0
xfeed_9032 0 1 decap_w0
xfeed_9031 0 1 decap_w0
xfeed_9030 0 1 decap_w0
xfeed_8509 0 1 decap_w0
xfeed_8508 0 1 decap_w0
xfeed_8507 0 1 decap_w0
xfeed_8506 0 1 decap_w0
xfeed_8505 0 1 decap_w0
xfeed_8504 0 1 decap_w0
xfeed_8503 0 1 decap_w0
xfeed_8502 0 1 decap_w0
xfeed_8501 0 1 decap_w0
xfeed_8500 0 1 decap_w0
xfeed_7899 0 1 decap_w0
xfeed_7898 0 1 decap_w0
xfeed_7897 0 1 decap_w0
xfeed_7896 0 1 decap_w0
xfeed_7895 0 1 decap_w0
xfeed_7894 0 1 decap_w0
xfeed_7893 0 1 tie
xfeed_7892 0 1 decap_w0
xfeed_7891 0 1 decap_w0
xfeed_7890 0 1 decap_w0
xfeed_3589 0 1 decap_w0
xfeed_3588 0 1 decap_w0
xfeed_3587 0 1 decap_w0
xfeed_3586 0 1 decap_w0
xfeed_3585 0 1 decap_w0
xfeed_3584 0 1 decap_w0
xfeed_3583 0 1 decap_w0
xfeed_3582 0 1 decap_w0
xfeed_3581 0 1 decap_w0
xfeed_3580 0 1 decap_w0
xsubckt_1201_or2_x1 0 1 1363 1374 1364 or2_x1
xsubckt_1091_and4_x1 0 1 1456 637 623 526 519 and4_x1
xsubckt_749_nand2_x0 0 1 1718 128 1766 nand2_x0
xsubckt_659_nand2_x0 0 1 101 2040 172 nand2_x0
xsubckt_358_and3_x1 0 1 390 424 423 391 and3_x1
xsubckt_1571_and21nor_x0 0 1 1023 1024 1117 2048 and21nor_x0
xsubckt_1602_and2_x1 0 1 992 995 993 and2_x1
xsubckt_1956_dff_x1 0 1 2049 1792 45 dff_x1
xsubckt_1958_dff_x1 0 1 2047 1790 45 dff_x1
xfeed_10408 0 1 tie
xfeed_10407 0 1 decap_w0
xfeed_10406 0 1 decap_w0
xfeed_10405 0 1 decap_w0
xfeed_10404 0 1 decap_w0
xfeed_10403 0 1 decap_w0
xfeed_10402 0 1 decap_w0
xfeed_10401 0 1 tie
xfeed_10400 0 1 decap_w0
xsubckt_715_and3_x1 0 1 1749 476 1759 1750 and3_x1
xsubckt_199_nor2_x0 0 1 559 1917 20 nor2_x0
xsubckt_1562_and3_x1 0 1 1032 1070 1050 1048 and3_x1
xsubckt_1671_and21nor_x0 0 1 923 1104 927 926 and21nor_x0
xfeed_9049 0 1 decap_w0
xfeed_9048 0 1 decap_w0
xfeed_9047 0 1 decap_w0
xfeed_9046 0 1 decap_w0
xfeed_9045 0 1 decap_w0
xfeed_9044 0 1 decap_w0
xfeed_9043 0 1 decap_w0
xfeed_9041 0 1 decap_w0
xfeed_9040 0 1 decap_w0
xfeed_8519 0 1 decap_w0
xfeed_8518 0 1 decap_w0
xfeed_8517 0 1 decap_w0
xfeed_8516 0 1 decap_w0
xfeed_8515 0 1 decap_w0
xfeed_8514 0 1 decap_w0
xfeed_8513 0 1 decap_w0
xfeed_8512 0 1 decap_w0
xfeed_8511 0 1 decap_w0
xfeed_8510 0 1 decap_w0
xfeed_4209 0 1 decap_w0
xfeed_4208 0 1 decap_w0
xfeed_4207 0 1 decap_w0
xfeed_4206 0 1 decap_w0
xfeed_4205 0 1 decap_w0
xfeed_4204 0 1 decap_w0
xfeed_4203 0 1 decap_w0
xfeed_4202 0 1 decap_w0
xfeed_4201 0 1 decap_w0
xfeed_4200 0 1 decap_w0
xfeed_3599 0 1 decap_w0
xfeed_3598 0 1 decap_w0
xfeed_3597 0 1 decap_w0
xfeed_3596 0 1 decap_w0
xfeed_3595 0 1 tie
xfeed_3594 0 1 decap_w0
xfeed_3593 0 1 decap_w0
xfeed_3592 0 1 decap_w0
xfeed_3591 0 1 decap_w0
xfeed_3590 0 1 decap_w0
xsubckt_863_mux2_x1 0 1 1618 2003 2053 446 mux2_x1
xsubckt_789_and3_x1 0 1 1683 1968 1749 1739 and3_x1
xsubckt_732_nand2_x0 0 1 2106 1765 1733 nand2_x0
xsubckt_201_nand3_x0 0 1 553 612 609 557 nand3_x0
xsubckt_1687_or3_x1 0 1 907 915 912 911 or3_x1
xfeed_10419 0 1 decap_w0
xfeed_10418 0 1 decap_w0
xfeed_10417 0 1 decap_w0
xfeed_10416 0 1 decap_w0
xfeed_10415 0 1 tie
xfeed_10414 0 1 decap_w0
xfeed_10413 0 1 decap_w0
xfeed_10412 0 1 decap_w0
xfeed_10411 0 1 decap_w0
xfeed_10410 0 1 decap_w0
xsubckt_1061_and2_x1 0 1 1481 1521 1482 and2_x1
xsubckt_945_or21nand_x0 0 1 1877 1574 1573 381 or21nand_x0
xsubckt_642_nand2_x0 0 1 117 2041 172 nand2_x0
xsubckt_299_nand2_x0 0 1 449 616 451 nand2_x0
xsubckt_214_and2_x1 0 1 540 549 541 and2_x1
xsubckt_623_and3_x1 0 1 134 139 138 135 and3_x1
xsubckt_1322_nand3_x0 0 1 1263 1916 1265 1264 nand3_x0
xsubckt_1444_and4_x1 0 1 1151 435 1628 1153 1152 and4_x1
xsubckt_1470_and3_x1 0 1 1126 1133 1131 1127 and3_x1
xsubckt_1771_and21nor_x0 0 1 823 940 937 834 and21nor_x0
xfeed_9059 0 1 decap_w0
xfeed_9058 0 1 decap_w0
xfeed_9057 0 1 decap_w0
xfeed_9056 0 1 decap_w0
xfeed_9055 0 1 decap_w0
xfeed_9054 0 1 decap_w0
xfeed_9053 0 1 decap_w0
xfeed_9052 0 1 decap_w0
xfeed_9051 0 1 decap_w0
xfeed_9050 0 1 decap_w0
xfeed_8529 0 1 decap_w0
xfeed_8528 0 1 decap_w0
xfeed_8527 0 1 decap_w0
xfeed_8526 0 1 decap_w0
xfeed_8525 0 1 decap_w0
xfeed_8524 0 1 decap_w0
xfeed_8521 0 1 decap_w0
xfeed_8520 0 1 decap_w0
xfeed_4219 0 1 decap_w0
xfeed_4218 0 1 decap_w0
xfeed_4217 0 1 decap_w0
xfeed_4216 0 1 decap_w0
xfeed_4215 0 1 tie
xfeed_4214 0 1 decap_w0
xfeed_4213 0 1 decap_w0
xfeed_4212 0 1 decap_w0
xfeed_4211 0 1 tie
xfeed_4210 0 1 decap_w0
xsubckt_1183_mux2_x1 0 1 1831 2083 1961 1916 mux2_x1
xsubckt_697_and3_x1 0 1 1767 537 198 1769 and3_x1
xsubckt_583_and4_x1 0 1 172 187 185 181 178 and4_x1
xsubckt_638_nand3_x0 0 1 121 2025 184 176 nand3_x0
xsubckt_1797_nexor2_x0 0 1 797 811 808 nexor2_x0
xfeed_10429 0 1 decap_w0
xfeed_10428 0 1 decap_w0
xfeed_10427 0 1 decap_w0
xfeed_10426 0 1 decap_w0
xfeed_10425 0 1 decap_w0
xfeed_10424 0 1 decap_w0
xfeed_10423 0 1 decap_w0
xfeed_10422 0 1 decap_w0
xfeed_10421 0 1 decap_w0
xfeed_10420 0 1 decap_w0
xsubckt_644_or21nand_x0 0 1 115 207 119 116 or21nand_x0
xsubckt_531_and3_x1 0 1 222 401 326 324 and3_x1
xsubckt_1313_or21nand_x0 0 1 1810 1281 1274 1272 or21nand_x0
xfeed_10 0 1 decap_w0
xfeed_11 0 1 decap_w0
xfeed_12 0 1 decap_w0
xfeed_14 0 1 tie
xfeed_15 0 1 decap_w0
xfeed_16 0 1 decap_w0
xfeed_17 0 1 decap_w0
xfeed_18 0 1 decap_w0
xfeed_19 0 1 decap_w0
xfeed_9069 0 1 decap_w0
xfeed_9068 0 1 decap_w0
xfeed_9067 0 1 decap_w0
xfeed_9066 0 1 decap_w0
xfeed_9065 0 1 decap_w0
xfeed_9064 0 1 decap_w0
xfeed_9063 0 1 decap_w0
xfeed_9062 0 1 decap_w0
xfeed_9061 0 1 decap_w0
xfeed_9060 0 1 decap_w0
xfeed_8539 0 1 decap_w0
xfeed_8538 0 1 decap_w0
xfeed_8536 0 1 decap_w0
xfeed_8535 0 1 decap_w0
xfeed_8534 0 1 decap_w0
xfeed_8533 0 1 decap_w0
xfeed_8532 0 1 decap_w0
xfeed_8531 0 1 decap_w0
xfeed_8530 0 1 decap_w0
xfeed_4229 0 1 decap_w0
xfeed_4228 0 1 decap_w0
xfeed_4227 0 1 decap_w0
xfeed_4226 0 1 decap_w0
xfeed_4225 0 1 decap_w0
xfeed_4224 0 1 decap_w0
xfeed_4223 0 1 decap_w0
xfeed_4222 0 1 decap_w0
xfeed_4221 0 1 decap_w0
xfeed_4220 0 1 decap_w0
xsubckt_1179_mux2_x1 0 1 1383 1384 2055 1391 mux2_x1
xsubckt_1166_and21nor_x0 0 1 1395 1396 1401 600 and21nor_x0
xsubckt_1048_nand4_x0 0 1 1492 660 646 641 640 nand4_x0
xsubckt_282_nand2_x0 0 1 466 558 468 nand2_x0
xsubckt_118_and2_x1 0 1 650 659 651 and2_x1
xsubckt_368_nand3_x0 0 1 381 652 526 383 nand3_x0
xsubckt_413_and4_x1 0 1 336 361 355 349 337 and4_x1
xfeed_10439 0 1 decap_w0
xfeed_10438 0 1 decap_w0
xfeed_10437 0 1 decap_w0
xfeed_10436 0 1 decap_w0
xfeed_10435 0 1 decap_w0
xfeed_10434 0 1 decap_w0
xfeed_10433 0 1 decap_w0
xfeed_10432 0 1 tie
xfeed_10431 0 1 decap_w0
xfeed_10430 0 1 decap_w0
xsubckt_1013_mux2_x1 0 1 1864 1540 1942 1576 mux2_x1
xsubckt_744_or21nand_x0 0 1 1722 2063 1742 1740 or21nand_x0
xsubckt_707_nand4_x0 0 1 1757 716 1923 712 599 nand4_x0
xsubckt_1413_or21nand_x0 0 1 1802 1192 1182 1180 or21nand_x0
xfeed_20 0 1 decap_w0
xfeed_21 0 1 decap_w0
xfeed_22 0 1 decap_w0
xfeed_23 0 1 decap_w0
xfeed_24 0 1 decap_w0
xfeed_25 0 1 decap_w0
xfeed_26 0 1 decap_w0
xfeed_27 0 1 decap_w0
xfeed_28 0 1 decap_w0
xfeed_29 0 1 tie
xfeed_9079 0 1 decap_w0
xfeed_9078 0 1 decap_w0
xfeed_9077 0 1 decap_w0
xfeed_9076 0 1 decap_w0
xfeed_9075 0 1 decap_w0
xfeed_9074 0 1 decap_w0
xfeed_9073 0 1 decap_w0
xfeed_9072 0 1 decap_w0
xfeed_9071 0 1 decap_w0
xfeed_9070 0 1 decap_w0
xfeed_8549 0 1 decap_w0
xfeed_8548 0 1 decap_w0
xfeed_8547 0 1 tie
xfeed_8546 0 1 decap_w0
xfeed_8545 0 1 decap_w0
xfeed_8544 0 1 decap_w0
xfeed_8543 0 1 decap_w0
xfeed_8542 0 1 decap_w0
xfeed_8541 0 1 decap_w0
xfeed_8540 0 1 tie
xfeed_4239 0 1 decap_w0
xfeed_4238 0 1 decap_w0
xfeed_4237 0 1 decap_w0
xfeed_4236 0 1 decap_w0
xfeed_4235 0 1 decap_w0
xfeed_4234 0 1 decap_w0
xfeed_4233 0 1 decap_w0
xfeed_4232 0 1 decap_w0
xfeed_4231 0 1 decap_w0
xfeed_4230 0 1 decap_w0
xfeed_3709 0 1 decap_w0
xfeed_3708 0 1 decap_w0
xfeed_3707 0 1 decap_w0
xfeed_3706 0 1 decap_w0
xfeed_3704 0 1 decap_w0
xfeed_3703 0 1 decap_w0
xfeed_3702 0 1 decap_w0
xfeed_3701 0 1 decap_w0
xfeed_3700 0 1 decap_w0
xsubckt_1209_or21nand_x0 0 1 1355 1361 1356 1375 or21nand_x0
xsubckt_958_and3_x1 0 1 1563 659 624 521 and3_x1
xsubckt_321_and4_x1 0 1 427 643 622 533 524 and4_x1
xsubckt_617_nand4_x0 0 1 140 145 144 143 142 nand4_x0
xfeed_10448 0 1 tie
xfeed_10447 0 1 decap_w0
xfeed_10446 0 1 decap_w0
xfeed_10445 0 1 decap_w0
xfeed_10444 0 1 decap_w0
xfeed_10443 0 1 decap_w0
xfeed_10442 0 1 decap_w0
xfeed_10441 0 1 decap_w0
xfeed_10440 0 1 decap_w0
xsubckt_1045_nand2_x0 0 1 1494 1920 1575 nand2_x0
xsubckt_351_nand3_x0 0 1 397 616 598 558 nand3_x0
xsubckt_395_and4_x1 0 1 354 686 605 600 591 and4_x1
xsubckt_1652_nand3_x0 0 1 942 1070 961 959 nand3_x0
xfeed_30 0 1 decap_w0
xfeed_31 0 1 decap_w0
xfeed_32 0 1 decap_w0
xfeed_33 0 1 tie
xfeed_34 0 1 decap_w0
xfeed_35 0 1 decap_w0
xfeed_36 0 1 decap_w0
xfeed_37 0 1 decap_w0
xfeed_38 0 1 decap_w0
xfeed_39 0 1 decap_w0
xfeed_9089 0 1 decap_w0
xfeed_9088 0 1 decap_w0
xfeed_9087 0 1 decap_w0
xfeed_9086 0 1 decap_w0
xfeed_9085 0 1 tie
xfeed_9084 0 1 decap_w0
xfeed_9083 0 1 decap_w0
xfeed_9082 0 1 decap_w0
xfeed_9081 0 1 decap_w0
xfeed_9080 0 1 decap_w0
xfeed_8559 0 1 decap_w0
xfeed_8558 0 1 decap_w0
xfeed_8557 0 1 tie
xfeed_8556 0 1 decap_w0
xfeed_8555 0 1 decap_w0
xfeed_8554 0 1 decap_w0
xfeed_8553 0 1 decap_w0
xfeed_8552 0 1 decap_w0
xfeed_8551 0 1 decap_w0
xfeed_8550 0 1 decap_w0
xfeed_4249 0 1 decap_w0
xfeed_4248 0 1 decap_w0
xfeed_4247 0 1 decap_w0
xfeed_4245 0 1 tie
xfeed_4244 0 1 decap_w0
xfeed_4243 0 1 decap_w0
xfeed_4242 0 1 decap_w0
xfeed_4241 0 1 decap_w0
xfeed_4240 0 1 decap_w0
xfeed_3719 0 1 decap_w0
xfeed_3718 0 1 decap_w0
xfeed_3717 0 1 decap_w0
xfeed_3716 0 1 decap_w0
xfeed_3715 0 1 decap_w0
xfeed_3714 0 1 tie
xfeed_3713 0 1 decap_w0
xfeed_3712 0 1 decap_w0
xfeed_3710 0 1 decap_w0
xsubckt_1226_and2_x1 0 1 1338 1340 1339 and2_x1
xsubckt_940_mux2_x1 0 1 1878 1952 623 774 mux2_x1
xsubckt_171_nand3_x0 0 1 587 680 599 589 nand3_x0
xsubckt_614_nand2_x0 0 1 143 2035 175 nand2_x0
xsubckt_633_nor2_x0 0 1 125 731 212 nor2_x0
xfeed_10459 0 1 tie
xfeed_10458 0 1 decap_w0
xfeed_10456 0 1 decap_w0
xfeed_10455 0 1 tie
xfeed_10454 0 1 decap_w0
xfeed_10453 0 1 decap_w0
xfeed_10452 0 1 decap_w0
xfeed_10451 0 1 decap_w0
xfeed_10450 0 1 decap_w0
xsubckt_106_nor2_x0 0 1 675 1929 1924 nor2_x0
xsubckt_1661_and2_x1 0 1 933 1663 934 and2_x1
xfeed_40 0 1 tie
xfeed_41 0 1 decap_w0
xfeed_43 0 1 decap_w0
xfeed_44 0 1 decap_w0
xfeed_45 0 1 decap_w0
xfeed_46 0 1 decap_w0
xfeed_9099 0 1 decap_w0
xfeed_9098 0 1 decap_w0
xfeed_9097 0 1 decap_w0
xfeed_9096 0 1 decap_w0
xfeed_9095 0 1 tie
xfeed_9094 0 1 decap_w0
xfeed_9093 0 1 decap_w0
xfeed_9092 0 1 decap_w0
xfeed_9091 0 1 decap_w0
xfeed_9090 0 1 decap_w0
xfeed_8569 0 1 decap_w0
xfeed_8568 0 1 tie
xfeed_8567 0 1 decap_w0
xfeed_8565 0 1 decap_w0
xfeed_8564 0 1 tie
xfeed_8563 0 1 decap_w0
xfeed_8562 0 1 decap_w0
xfeed_8561 0 1 decap_w0
xfeed_8560 0 1 decap_w0
xfeed_4259 0 1 decap_w0
xfeed_4258 0 1 decap_w0
xfeed_4257 0 1 tie
xfeed_4256 0 1 decap_w0
xfeed_4255 0 1 decap_w0
xfeed_4254 0 1 decap_w0
xfeed_4253 0 1 decap_w0
xfeed_4252 0 1 decap_w0
xfeed_4251 0 1 decap_w0
xfeed_4250 0 1 tie
xfeed_3729 0 1 decap_w0
xfeed_3728 0 1 decap_w0
xfeed_3727 0 1 decap_w0
xfeed_3726 0 1 decap_w0
xfeed_3725 0 1 decap_w0
xfeed_3724 0 1 decap_w0
xfeed_3723 0 1 decap_w0
xfeed_3722 0 1 decap_w0
xfeed_3721 0 1 decap_w0
xfeed_3720 0 1 decap_w0
xsubckt_698_nand3_x0 0 1 1766 537 198 1769 nand3_x0
xsubckt_660_and4_x1 0 1 100 104 103 102 101 and4_x1
xsubckt_1402_or2_x1 0 1 1190 692 1323 or2_x1
xsubckt_1409_or21nand_x0 0 1 1183 1185 1197 1206 or21nand_x0
xsubckt_1543_and3_x1 0 1 1051 1970 679 595 and3_x1
xfeed_47 0 1 decap_w0
xfeed_48 0 1 decap_w0
xfeed_49 0 1 decap_w0
xfeed_10469 0 1 tie
xfeed_10468 0 1 decap_w0
xfeed_10467 0 1 decap_w0
xfeed_10465 0 1 decap_w0
xfeed_10464 0 1 decap_w0
xfeed_10463 0 1 decap_w0
xfeed_10462 0 1 decap_w0
xfeed_10461 0 1 decap_w0
xfeed_10460 0 1 decap_w0
xsubckt_1705_mux2_x1 0 1 889 894 892 901 mux2_x1
xfeed_50 0 1 tie
xfeed_51 0 1 decap_w0
xfeed_52 0 1 decap_w0
xfeed_53 0 1 decap_w0
xfeed_8579 0 1 decap_w0
xfeed_8578 0 1 decap_w0
xfeed_8577 0 1 decap_w0
xfeed_8576 0 1 decap_w0
xfeed_8575 0 1 decap_w0
xfeed_8574 0 1 decap_w0
xfeed_8573 0 1 tie
xfeed_8572 0 1 decap_w0
xfeed_8571 0 1 decap_w0
xfeed_8570 0 1 decap_w0
xfeed_4269 0 1 decap_w0
xfeed_4268 0 1 decap_w0
xfeed_4267 0 1 decap_w0
xfeed_4266 0 1 decap_w0
xfeed_4265 0 1 decap_w0
xfeed_4264 0 1 tie
xfeed_4263 0 1 decap_w0
xfeed_4262 0 1 decap_w0
xfeed_4261 0 1 decap_w0
xfeed_4260 0 1 decap_w0
xfeed_3739 0 1 decap_w0
xfeed_3738 0 1 decap_w0
xfeed_3737 0 1 decap_w0
xfeed_3736 0 1 decap_w0
xfeed_3735 0 1 decap_w0
xfeed_3734 0 1 decap_w0
xfeed_3733 0 1 decap_w0
xfeed_3732 0 1 decap_w0
xfeed_3731 0 1 decap_w0
xfeed_3730 0 1 decap_w0
xsubckt_1165_and21nor_x0 0 1 1396 1397 1400 600 and21nor_x0
xsubckt_1016_and3_x1 0 1 1515 661 646 527 and3_x1
xsubckt_857_nand4_x0 0 1 1624 780 682 674 670 nand4_x0
xsubckt_1465_nand2_x0 0 1 1131 2055 1132 nand2_x0
xsubckt_1813_or21nand_x0 0 1 1792 789 788 787 or21nand_x0
xfeed_54 0 1 decap_w0
xfeed_55 0 1 decap_w0
xfeed_56 0 1 decap_w0
xfeed_57 0 1 tie
xfeed_59 0 1 decap_w0
xfeed_10476 0 1 tie
xfeed_10475 0 1 decap_w0
xfeed_10474 0 1 decap_w0
xfeed_10473 0 1 decap_w0
xfeed_10472 0 1 decap_w0
xfeed_10471 0 1 decap_w0
xsubckt_181_and2_x1 0 1 577 582 578 and2_x1
xsubckt_45_inv_x0 0 1 737 1943 inv_x0
xsubckt_43_inv_x0 0 1 739 1945 inv_x0
xsubckt_41_inv_x0 0 1 741 2067 inv_x0
xsubckt_564_and4_x1 0 1 191 501 462 456 403 and4_x1
xsubckt_1285_nand2_x0 0 1 1297 784 1983 nand2_x0
xsubckt_1499_and4_x1 0 1 1097 467 198 1769 1368 and4_x1
xfeed_60 0 1 decap_w0
xfeed_10479 0 1 decap_w0
xfeed_10478 0 1 decap_w0
xfeed_10477 0 1 decap_w0
xfeed_8589 0 1 decap_w0
xfeed_8588 0 1 decap_w0
xfeed_8587 0 1 decap_w0
xfeed_8586 0 1 decap_w0
xfeed_8585 0 1 decap_w0
xfeed_8584 0 1 decap_w0
xfeed_8583 0 1 decap_w0
xfeed_8582 0 1 decap_w0
xfeed_8581 0 1 decap_w0
xfeed_8580 0 1 decap_w0
xfeed_4279 0 1 decap_w0
xfeed_4278 0 1 decap_w0
xfeed_4277 0 1 decap_w0
xfeed_4276 0 1 decap_w0
xfeed_4275 0 1 decap_w0
xfeed_4274 0 1 decap_w0
xfeed_4273 0 1 decap_w0
xfeed_4272 0 1 decap_w0
xfeed_4271 0 1 tie
xfeed_4270 0 1 decap_w0
xfeed_3749 0 1 decap_w0
xfeed_3748 0 1 decap_w0
xfeed_3747 0 1 decap_w0
xfeed_3746 0 1 decap_w0
xfeed_3745 0 1 decap_w0
xfeed_3744 0 1 decap_w0
xfeed_3743 0 1 decap_w0
xfeed_3742 0 1 decap_w0
xfeed_3741 0 1 decap_w0
xfeed_3740 0 1 decap_w0
xsubckt_1195_nand2_x0 0 1 1369 1373 1372 nand2_x0
xsubckt_49_inv_x0 0 1 733 1967 inv_x0
xsubckt_47_inv_x0 0 1 735 1941 inv_x0
xsubckt_587_nand4_x0 0 1 168 174 173 171 170 nand4_x0
xsubckt_1473_and2_x1 0 1 1123 1380 1139 and2_x1
xsubckt_1624_nand3_x0 0 1 970 977 974 973 nand3_x0
xfeed_62 0 1 decap_w0
xfeed_63 0 1 decap_w0
xfeed_64 0 1 tie
xfeed_65 0 1 decap_w0
xfeed_66 0 1 decap_w0
xfeed_67 0 1 decap_w0
xfeed_68 0 1 tie
xfeed_69 0 1 decap_w0
xfeed_10483 0 1 decap_w0
xfeed_10482 0 1 decap_w0
xfeed_10481 0 1 decap_w0
xfeed_10480 0 1 decap_w0
xsubckt_764_nand2_x0 0 1 2096 1711 1705 nand2_x0
xsubckt_1469_and2_x1 0 1 1127 1129 1128 and2_x1
xfeed_10489 0 1 decap_w0
xfeed_10488 0 1 decap_w0
xfeed_10487 0 1 decap_w0
xfeed_10486 0 1 decap_w0
xfeed_10485 0 1 decap_w0
xfeed_10484 0 1 decap_w0
xfeed_9209 0 1 decap_w0
xfeed_9208 0 1 decap_w0
xfeed_9207 0 1 decap_w0
xfeed_9206 0 1 decap_w0
xfeed_9205 0 1 decap_w0
xfeed_9204 0 1 decap_w0
xfeed_9203 0 1 tie
xfeed_9202 0 1 decap_w0
xfeed_9201 0 1 decap_w0
xfeed_9200 0 1 decap_w0
xfeed_8599 0 1 decap_w0
xfeed_8598 0 1 tie
xfeed_8597 0 1 decap_w0
xfeed_8596 0 1 decap_w0
xfeed_8595 0 1 decap_w0
xfeed_8594 0 1 decap_w0
xfeed_8593 0 1 decap_w0
xfeed_8592 0 1 decap_w0
xfeed_8591 0 1 decap_w0
xfeed_8590 0 1 tie
xfeed_4289 0 1 decap_w0
xfeed_4288 0 1 tie
xfeed_4287 0 1 decap_w0
xfeed_4286 0 1 decap_w0
xfeed_4285 0 1 decap_w0
xfeed_4284 0 1 decap_w0
xfeed_4283 0 1 decap_w0
xfeed_4282 0 1 decap_w0
xfeed_4281 0 1 tie
xfeed_4280 0 1 decap_w0
xfeed_3759 0 1 decap_w0
xfeed_3758 0 1 decap_w0
xfeed_3757 0 1 decap_w0
xfeed_3756 0 1 decap_w0
xfeed_3755 0 1 decap_w0
xfeed_3754 0 1 decap_w0
xfeed_3753 0 1 decap_w0
xfeed_3752 0 1 tie
xfeed_3751 0 1 decap_w0
xfeed_3750 0 1 decap_w0
xsubckt_804_and21nor_x0 0 1 1669 746 600 1745 and21nor_x0
xsubckt_139_nand4_x0 0 1 629 650 644 638 632 nand4_x0
xsubckt_1709_or21nand_x0 0 1 885 1067 896 1072 or21nand_x0
xfeed_70 0 1 decap_w0
xfeed_71 0 1 decap_w0
xfeed_72 0 1 decap_w0
xfeed_73 0 1 decap_w0
xfeed_74 0 1 decap_w0
xfeed_76 0 1 decap_w0
xfeed_77 0 1 decap_w0
xfeed_78 0 1 decap_w0
xfeed_79 0 1 decap_w0
xfeed_11109 0 1 decap_w0
xfeed_11108 0 1 decap_w0
xfeed_11107 0 1 decap_w0
xfeed_11106 0 1 decap_w0
xfeed_11105 0 1 decap_w0
xfeed_11104 0 1 decap_w0
xfeed_11103 0 1 decap_w0
xfeed_11102 0 1 decap_w0
xfeed_11101 0 1 decap_w0
xfeed_11100 0 1 decap_w0
xfeed_10490 0 1 decap_w0
xsubckt_1000_nand2_x0 0 1 1529 630 1530 nand2_x0
xsubckt_584_nand2_x0 0 1 171 2045 172 nand2_x0
xcmpt_abc_11867_new_n473_hfns_0 0 1 617 615 buf_x4
xcmpt_abc_11867_new_n473_hfns_1 0 1 616 615 buf_x4
xcmpt_abc_11867_new_n473_hfns_2 0 1 615 618 buf_x4
xfeed_10499 0 1 decap_w0
xfeed_10498 0 1 decap_w0
xfeed_10497 0 1 decap_w0
xfeed_10496 0 1 decap_w0
xfeed_10495 0 1 decap_w0
xfeed_10494 0 1 tie
xfeed_10493 0 1 decap_w0
xfeed_10492 0 1 decap_w0
xfeed_10491 0 1 decap_w0
xfeed_9219 0 1 decap_w0
xfeed_9218 0 1 decap_w0
xfeed_9217 0 1 decap_w0
xfeed_9216 0 1 decap_w0
xfeed_9215 0 1 decap_w0
xfeed_9214 0 1 decap_w0
xfeed_9213 0 1 decap_w0
xfeed_9212 0 1 decap_w0
xfeed_9211 0 1 decap_w0
xfeed_9210 0 1 tie
xfeed_4299 0 1 decap_w0
xfeed_4298 0 1 decap_w0
xfeed_4297 0 1 decap_w0
xfeed_4296 0 1 decap_w0
xfeed_4295 0 1 tie
xfeed_4294 0 1 decap_w0
xfeed_4293 0 1 decap_w0
xfeed_4292 0 1 decap_w0
xfeed_4291 0 1 decap_w0
xfeed_4290 0 1 decap_w0
xfeed_3768 0 1 decap_w0
xfeed_3767 0 1 decap_w0
xfeed_3766 0 1 decap_w0
xfeed_3765 0 1 decap_w0
xfeed_3764 0 1 decap_w0
xfeed_3763 0 1 decap_w0
xfeed_3762 0 1 decap_w0
xfeed_3761 0 1 decap_w0
xfeed_3760 0 1 decap_w0
xsubckt_1211_and2_x1 0 1 1353 1756 1354 and2_x1
xsubckt_1084_nand3_x0 0 1 1461 643 533 1473 nand3_x0
xsubckt_692_nor2_x0 0 1 1771 1773 1772 nor2_x0
xsubckt_226_nand2_x0 0 1 525 661 527 nand2_x0
xsubckt_141_or21nand_x0 0 1 627 661 654 651 or21nand_x0
xcmpt_abc_11867_new_n477_hfns_0 0 1 610 607 buf_x4
xcmpt_abc_11867_new_n477_hfns_1 0 1 609 607 buf_x4
xcmpt_abc_11867_new_n477_hfns_2 0 1 608 607 buf_x4
xcmpt_abc_11867_new_n477_hfns_3 0 1 607 611 buf_x4
xfeed_80 0 1 decap_w0
xfeed_81 0 1 decap_w0
xfeed_82 0 1 decap_w0
xfeed_83 0 1 tie
xfeed_84 0 1 decap_w0
xfeed_85 0 1 decap_w0
xfeed_86 0 1 decap_w0
xfeed_87 0 1 decap_w0
xfeed_88 0 1 decap_w0
xfeed_89 0 1 decap_w0
xfeed_11119 0 1 decap_w0
xfeed_11118 0 1 decap_w0
xfeed_11117 0 1 decap_w0
xfeed_11116 0 1 decap_w0
xfeed_11115 0 1 decap_w0
xfeed_11114 0 1 decap_w0
xfeed_11113 0 1 decap_w0
xfeed_11112 0 1 decap_w0
xfeed_11111 0 1 decap_w0
xfeed_11110 0 1 decap_w0
xsubckt_847_and3_x1 0 1 1632 1975 1749 1739 and3_x1
xsubckt_129_mux2_x1 0 1 639 1994 2003 1986 mux2_x1
xsubckt_136_nand2_x0 0 1 632 661 634 nand2_x0
xsubckt_1961_dff_x1 0 1 2057 1787 45 dff_x1
xfeed_9229 0 1 decap_w0
xfeed_9228 0 1 decap_w0
xfeed_9227 0 1 decap_w0
xfeed_9226 0 1 decap_w0
xfeed_9225 0 1 decap_w0
xfeed_9224 0 1 decap_w0
xfeed_9223 0 1 decap_w0
xfeed_9222 0 1 decap_w0
xfeed_9221 0 1 decap_w0
xfeed_9220 0 1 decap_w0
xfeed_3775 0 1 decap_w0
xfeed_3774 0 1 decap_w0
xfeed_3772 0 1 decap_w0
xfeed_3771 0 1 decap_w0
xfeed_3770 0 1 decap_w0
xsubckt_921_mux2_x1 0 1 1895 1605 2035 1579 mux2_x1
xsubckt_210_and4_x1 0 1 544 712 1926 674 670 and4_x1
xsubckt_1347_nand2_x0 0 1 1241 1968 1316 nand2_x0
xfeed_90 0 1 tie
xfeed_91 0 1 decap_w0
xfeed_92 0 1 decap_w0
xfeed_93 0 1 decap_w0
xfeed_94 0 1 decap_w0
xfeed_95 0 1 decap_w0
xfeed_96 0 1 decap_w0
xfeed_97 0 1 decap_w0
xfeed_98 0 1 decap_w0
xfeed_99 0 1 decap_w0
xfeed_11129 0 1 decap_w0
xfeed_11128 0 1 decap_w0
xfeed_11127 0 1 decap_w0
xfeed_11126 0 1 decap_w0
xfeed_11125 0 1 decap_w0
xfeed_11124 0 1 decap_w0
xfeed_11123 0 1 decap_w0
xfeed_11122 0 1 decap_w0
xfeed_11121 0 1 decap_w0
xfeed_11120 0 1 decap_w0
xfeed_3779 0 1 decap_w0
xfeed_3778 0 1 decap_w0
xfeed_3777 0 1 tie
xfeed_3776 0 1 decap_w0
xsubckt_1241_mux2_x1 0 1 1820 2104 2071 1334 mux2_x1
xsubckt_917_mux2_x1 0 1 1898 1581 2038 1580 mux2_x1
xsubckt_206_and4_x1 0 1 548 716 1924 682 670 and4_x1
xsubckt_473_nand3_x0 0 1 277 686 608 451 nand3_x0
xsubckt_559_nand4_x0 0 1 196 1927 713 711 673 nand4_x0
xsubckt_1665_and21nor_x0 0 1 929 930 1121 140 and21nor_x0
xsubckt_1812_or21nand_x0 0 1 787 1917 821 818 or21nand_x0
xfeed_9239 0 1 decap_w0
xfeed_9238 0 1 decap_w0
xfeed_9237 0 1 decap_w0
xfeed_9236 0 1 decap_w0
xfeed_9235 0 1 decap_w0
xfeed_9234 0 1 decap_w0
xfeed_9233 0 1 decap_w0
xfeed_9232 0 1 decap_w0
xfeed_9231 0 1 decap_w0
xfeed_9230 0 1 decap_w0
xfeed_8709 0 1 decap_w0
xfeed_8708 0 1 decap_w0
xfeed_8707 0 1 decap_w0
xfeed_8705 0 1 decap_w0
xfeed_8704 0 1 tie
xfeed_8703 0 1 decap_w0
xfeed_8702 0 1 decap_w0
xfeed_8701 0 1 decap_w0
xfeed_8700 0 1 decap_w0
xfeed_3782 0 1 decap_w0
xfeed_3781 0 1 decap_w0
xfeed_3780 0 1 decap_w0
xsubckt_1077_nand2_x0 0 1 1467 652 644 nand2_x0
xsubckt_1506_nand3_x0 0 1 1090 1103 1099 1095 nand3_x0
xsubckt_1684_nand3_x0 0 1 910 1070 927 926 nand3_x0
xfeed_11139 0 1 decap_w0
xfeed_11138 0 1 decap_w0
xfeed_11137 0 1 decap_w0
xfeed_11136 0 1 tie
xfeed_11135 0 1 decap_w0
xfeed_11133 0 1 decap_w0
xfeed_11132 0 1 decap_w0
xfeed_11131 0 1 decap_w0
xfeed_11130 0 1 decap_w0
xfeed_10609 0 1 decap_w0
xfeed_10608 0 1 decap_w0
xfeed_10607 0 1 decap_w0
xfeed_10606 0 1 tie
xfeed_10605 0 1 decap_w0
xfeed_10604 0 1 decap_w0
xfeed_10603 0 1 decap_w0
xfeed_10602 0 1 decap_w0
xfeed_10601 0 1 tie
xfeed_10600 0 1 decap_w0
xfeed_3789 0 1 decap_w0
xfeed_3788 0 1 decap_w0
xfeed_3787 0 1 decap_w0
xfeed_3786 0 1 decap_w0
xfeed_3785 0 1 decap_w0
xfeed_3784 0 1 decap_w0
xfeed_3783 0 1 decap_w0
xsubckt_1237_mux2_x1 0 1 1824 2094 2059 1334 mux2_x1
xsubckt_777_and2_x1 0 1 1693 1695 1694 and2_x1
xsubckt_1326_nand3_x0 0 1 1260 2059 666 657 nand3_x0
xfeed_9249 0 1 decap_w0
xfeed_9248 0 1 decap_w0
xfeed_9247 0 1 decap_w0
xfeed_9246 0 1 decap_w0
xfeed_9245 0 1 decap_w0
xfeed_9244 0 1 decap_w0
xfeed_9243 0 1 tie
xfeed_9242 0 1 decap_w0
xfeed_9241 0 1 decap_w0
xfeed_9240 0 1 decap_w0
xfeed_8719 0 1 decap_w0
xfeed_8718 0 1 tie
xfeed_8717 0 1 decap_w0
xfeed_8716 0 1 decap_w0
xfeed_8715 0 1 decap_w0
xfeed_8714 0 1 decap_w0
xfeed_8713 0 1 decap_w0
xfeed_8712 0 1 decap_w0
xfeed_8711 0 1 tie
xfeed_8710 0 1 decap_w0
xfeed_4409 0 1 decap_w0
xfeed_4408 0 1 decap_w0
xfeed_4407 0 1 decap_w0
xfeed_4406 0 1 decap_w0
xfeed_4405 0 1 decap_w0
xfeed_4404 0 1 decap_w0
xfeed_4403 0 1 tie
xfeed_4402 0 1 decap_w0
xfeed_4401 0 1 decap_w0
xfeed_4400 0 1 decap_w0
xsubckt_695_and21nor_x0 0 1 1769 408 460 609 and21nor_x0
xsubckt_556_nand2_x0 0 1 199 505 438 nand2_x0
xfeed_11149 0 1 decap_w0
xfeed_11148 0 1 decap_w0
xfeed_11147 0 1 decap_w0
xfeed_11146 0 1 decap_w0
xfeed_11145 0 1 decap_w0
xfeed_11144 0 1 decap_w0
xfeed_11143 0 1 decap_w0
xfeed_11142 0 1 decap_w0
xfeed_11141 0 1 decap_w0
xfeed_11140 0 1 decap_w0
xfeed_10616 0 1 decap_w0
xfeed_10615 0 1 decap_w0
xfeed_10613 0 1 decap_w0
xfeed_10612 0 1 decap_w0
xfeed_10611 0 1 decap_w0
xfeed_10610 0 1 decap_w0
xfeed_3799 0 1 decap_w0
xfeed_3798 0 1 decap_w0
xfeed_3797 0 1 decap_w0
xfeed_3796 0 1 decap_w0
xfeed_3795 0 1 decap_w0
xfeed_3794 0 1 decap_w0
xfeed_3792 0 1 decap_w0
xfeed_3791 0 1 decap_w0
xfeed_3790 0 1 decap_w0
xsubckt_983_nand3_x0 0 1 1544 660 527 521 nand3_x0
xsubckt_685_and2_x1 0 1 1778 1780 1779 and2_x1
xsubckt_545_and4_x1 0 1 209 449 410 325 210 and4_x1
xsubckt_1307_or21nand_x0 0 1 1277 1278 1322 763 or21nand_x0
xsubckt_1392_and4_x1 0 1 1199 435 1656 1201 1200 and4_x1
xfeed_10619 0 1 decap_w0
xfeed_10618 0 1 decap_w0
xfeed_10617 0 1 decap_w0
xfeed_9259 0 1 decap_w0
xfeed_9258 0 1 decap_w0
xfeed_9257 0 1 decap_w0
xfeed_9256 0 1 decap_w0
xfeed_9255 0 1 tie
xfeed_9254 0 1 decap_w0
xfeed_9253 0 1 decap_w0
xfeed_9252 0 1 decap_w0
xfeed_9251 0 1 decap_w0
xfeed_9250 0 1 decap_w0
xfeed_8729 0 1 decap_w0
xfeed_8728 0 1 tie
xfeed_8727 0 1 decap_w0
xfeed_8726 0 1 decap_w0
xfeed_8725 0 1 decap_w0
xfeed_8724 0 1 decap_w0
xfeed_8723 0 1 decap_w0
xfeed_8722 0 1 decap_w0
xfeed_8721 0 1 decap_w0
xfeed_8720 0 1 decap_w0
xfeed_4419 0 1 decap_w0
xfeed_4418 0 1 decap_w0
xfeed_4417 0 1 decap_w0
xfeed_4416 0 1 decap_w0
xfeed_4415 0 1 tie
xfeed_4414 0 1 decap_w0
xfeed_4413 0 1 decap_w0
xfeed_4412 0 1 decap_w0
xfeed_4411 0 1 decap_w0
xfeed_4410 0 1 tie
xsubckt_1210_or21nand_x0 0 1 1354 681 594 421 or21nand_x0
xsubckt_903_and21nor_x0 0 1 1585 1590 1589 1596 and21nor_x0
xsubckt_882_nexor2_x0 0 1 1602 764 1603 nexor2_x0
xsubckt_795_and21nor_x0 0 1 1677 696 1755 1754 and21nor_x0
xsubckt_1811_and2_x1 0 1 788 821 818 and2_x1
xfeed_11159 0 1 decap_w0
xfeed_11158 0 1 decap_w0
xfeed_11157 0 1 decap_w0
xfeed_11156 0 1 decap_w0
xfeed_11155 0 1 decap_w0
xfeed_11154 0 1 decap_w0
xfeed_11153 0 1 decap_w0
xfeed_11152 0 1 decap_w0
xfeed_11151 0 1 decap_w0
xfeed_11150 0 1 decap_w0
xfeed_10623 0 1 decap_w0
xfeed_10622 0 1 decap_w0
xfeed_10621 0 1 tie
xfeed_10620 0 1 decap_w0
xsubckt_453_and4_x1 0 1 297 533 518 384 360 and4_x1
xsubckt_625_nand3_x0 0 1 133 2026 184 176 nand3_x0
xfeed_10629 0 1 decap_w0
xfeed_10628 0 1 decap_w0
xfeed_10627 0 1 decap_w0
xfeed_10626 0 1 decap_w0
xfeed_10625 0 1 decap_w0
xfeed_10624 0 1 decap_w0
xfeed_9269 0 1 decap_w0
xfeed_9268 0 1 decap_w0
xfeed_9267 0 1 decap_w0
xfeed_9266 0 1 decap_w0
xfeed_9265 0 1 decap_w0
xfeed_9264 0 1 decap_w0
xfeed_9263 0 1 decap_w0
xfeed_9262 0 1 decap_w0
xfeed_9261 0 1 decap_w0
xfeed_9260 0 1 decap_w0
xfeed_8739 0 1 decap_w0
xfeed_8738 0 1 decap_w0
xfeed_8737 0 1 decap_w0
xfeed_8736 0 1 decap_w0
xfeed_8735 0 1 decap_w0
xfeed_8734 0 1 decap_w0
xfeed_8733 0 1 decap_w0
xfeed_8732 0 1 decap_w0
xfeed_8731 0 1 decap_w0
xfeed_8730 0 1 decap_w0
xfeed_4429 0 1 decap_w0
xfeed_4428 0 1 decap_w0
xfeed_4427 0 1 decap_w0
xfeed_4426 0 1 decap_w0
xfeed_4425 0 1 decap_w0
xfeed_4424 0 1 decap_w0
xfeed_4423 0 1 decap_w0
xfeed_4422 0 1 tie
xfeed_4421 0 1 decap_w0
xfeed_4420 0 1 decap_w0
xsubckt_1049_mux2_x1 0 1 1491 633 644 638 mux2_x1
xsubckt_739_nor3_x0 0 1 1726 1731 1730 1727 nor3_x0
xsubckt_1534_nor2_x0 0 1 1060 1083 1062 nor2_x0
xfeed_11169 0 1 tie
xfeed_11168 0 1 decap_w0
xfeed_11167 0 1 decap_w0
xfeed_11166 0 1 decap_w0
xfeed_11165 0 1 decap_w0
xfeed_11164 0 1 decap_w0
xfeed_11163 0 1 decap_w0
xfeed_11162 0 1 decap_w0
xfeed_11161 0 1 decap_w0
xfeed_11160 0 1 decap_w0
xfeed_10630 0 1 decap_w0
xsubckt_976_nand2_x0 0 1 1550 382 1552 nand2_x0
xsubckt_821_or4_x1 0 1 1654 1659 1658 1657 1655 or4_x1
xsubckt_114_mux2_x1 0 1 654 1990 1999 1986 mux2_x1
xsubckt_355_nand3_x0 0 1 393 680 598 558 nand3_x0
xfeed_10639 0 1 decap_w0
xfeed_10638 0 1 decap_w0
xfeed_10637 0 1 decap_w0
xfeed_10636 0 1 decap_w0
xfeed_10635 0 1 decap_w0
xfeed_10634 0 1 decap_w0
xfeed_10633 0 1 decap_w0
xfeed_10632 0 1 decap_w0
xfeed_10631 0 1 decap_w0
xfeed_9279 0 1 decap_w0
xfeed_9278 0 1 decap_w0
xfeed_9277 0 1 decap_w0
xfeed_9276 0 1 decap_w0
xfeed_9275 0 1 decap_w0
xfeed_9274 0 1 decap_w0
xfeed_9273 0 1 decap_w0
xfeed_9272 0 1 decap_w0
xfeed_9271 0 1 decap_w0
xfeed_9270 0 1 decap_w0
xfeed_8747 0 1 decap_w0
xfeed_8746 0 1 decap_w0
xfeed_8745 0 1 decap_w0
xfeed_8744 0 1 decap_w0
xfeed_8743 0 1 decap_w0
xfeed_8742 0 1 decap_w0
xfeed_8741 0 1 decap_w0
xfeed_8740 0 1 decap_w0
xfeed_4439 0 1 decap_w0
xfeed_4438 0 1 decap_w0
xfeed_4437 0 1 decap_w0
xfeed_4436 0 1 decap_w0
xfeed_4435 0 1 decap_w0
xfeed_4434 0 1 decap_w0
xfeed_4433 0 1 decap_w0
xfeed_4432 0 1 decap_w0
xfeed_4431 0 1 decap_w0
xfeed_4430 0 1 decap_w0
xfeed_3906 0 1 decap_w0
xfeed_3905 0 1 decap_w0
xfeed_3904 0 1 decap_w0
xfeed_3903 0 1 decap_w0
xfeed_3902 0 1 decap_w0
xfeed_3901 0 1 decap_w0
xfeed_3900 0 1 tie
xsubckt_1263_and21nor_x0 0 1 1317 1331 1322 1319 and21nor_x0
xsubckt_1212_nand2_x0 0 1 1352 1363 1355 nand2_x0
xsubckt_829_or4_x1 0 1 1647 1652 1651 1650 1648 or4_x1
xsubckt_265_nand3_x0 0 1 483 609 557 495 nand3_x0
xsubckt_357_and4_x1 0 1 391 412 406 396 392 and4_x1
xsubckt_604_nand4_x0 0 1 152 157 156 155 154 nand4_x0
xsubckt_1390_nand2_x0 0 1 1201 2050 479 nand2_x0
xsubckt_1566_nand3_x0 0 1 1028 1037 1033 1031 nand3_x0
xfeed_11176 0 1 decap_w0
xfeed_11175 0 1 decap_w0
xfeed_11174 0 1 decap_w0
xfeed_11173 0 1 decap_w0
xfeed_11172 0 1 decap_w0
xfeed_11171 0 1 decap_w0
xfeed_11170 0 1 decap_w0
xfeed_8749 0 1 decap_w0
xfeed_8748 0 1 decap_w0
xfeed_3909 0 1 decap_w0
xsubckt_902_mux2_x1 0 1 1907 2015 1586 1619 mux2_x1
xsubckt_1510_or21nand_x0 0 1 1086 1088 1111 1120 or21nand_x0
xsubckt_1819_dff_x1 0 1 2021 1913 32 dff_x1
xfeed_11179 0 1 decap_w0
xfeed_11178 0 1 decap_w0
xfeed_11177 0 1 decap_w0
xfeed_10649 0 1 decap_w0
xfeed_10648 0 1 decap_w0
xfeed_10647 0 1 decap_w0
xfeed_10646 0 1 decap_w0
xfeed_10645 0 1 decap_w0
xfeed_10644 0 1 decap_w0
xfeed_10643 0 1 decap_w0
xfeed_10642 0 1 decap_w0
xfeed_10641 0 1 decap_w0
xfeed_10640 0 1 decap_w0
xfeed_9289 0 1 decap_w0
xfeed_9288 0 1 decap_w0
xfeed_9287 0 1 decap_w0
xfeed_9286 0 1 decap_w0
xfeed_9285 0 1 decap_w0
xfeed_9284 0 1 decap_w0
xfeed_9283 0 1 decap_w0
xfeed_9282 0 1 decap_w0
xfeed_9281 0 1 decap_w0
xfeed_9280 0 1 decap_w0
xfeed_8754 0 1 tie
xfeed_8753 0 1 decap_w0
xfeed_8752 0 1 decap_w0
xfeed_8751 0 1 decap_w0
xfeed_8750 0 1 decap_w0
xfeed_4449 0 1 decap_w0
xfeed_4448 0 1 decap_w0
xfeed_4447 0 1 decap_w0
xfeed_4446 0 1 decap_w0
xfeed_4445 0 1 decap_w0
xfeed_4444 0 1 decap_w0
xfeed_4443 0 1 decap_w0
xfeed_4442 0 1 decap_w0
xfeed_4441 0 1 decap_w0
xfeed_4440 0 1 decap_w0
xfeed_3915 0 1 decap_w0
xfeed_3914 0 1 decap_w0
xfeed_3913 0 1 tie
xfeed_3912 0 1 decap_w0
xfeed_3910 0 1 decap_w0
xsubckt_1599_or21nand_x0 0 1 995 1121 116 119 or21nand_x0
xsubckt_1697_and2_x1 0 1 897 899 898 and2_x1
xfeed_11183 0 1 decap_w0
xfeed_11182 0 1 decap_w0
xfeed_11181 0 1 tie
xfeed_11180 0 1 decap_w0
xfeed_8759 0 1 tie
xfeed_8758 0 1 decap_w0
xfeed_8757 0 1 decap_w0
xfeed_8756 0 1 decap_w0
xfeed_8755 0 1 decap_w0
xfeed_3919 0 1 decap_w0
xfeed_3918 0 1 decap_w0
xfeed_3917 0 1 decap_w0
xfeed_3916 0 1 decap_w0
xsubckt_258_nand2_x0 0 1 493 617 495 nand2_x0
xsubckt_213_and3_x1 0 1 541 546 545 542 and3_x1
xsubckt_601_nand2_x0 0 1 155 2036 175 nand2_x0
xsubckt_637_or21nand_x0 0 1 2079 122 129 206 or21nand_x0
xsubckt_1610_or21nand_x0 0 1 984 1105 990 988 or21nand_x0
xsubckt_1635_nand4_x0 0 1 959 2000 1128 1098 1097 nand4_x0
xfeed_11189 0 1 decap_w0
xfeed_11188 0 1 decap_w0
xfeed_11187 0 1 decap_w0
xfeed_11186 0 1 tie
xfeed_11185 0 1 decap_w0
xfeed_11184 0 1 decap_w0
xfeed_10659 0 1 decap_w0
xfeed_10658 0 1 decap_w0
xfeed_10657 0 1 decap_w0
xfeed_10656 0 1 decap_w0
xfeed_10655 0 1 decap_w0
xfeed_10653 0 1 decap_w0
xfeed_10652 0 1 decap_w0
xfeed_10651 0 1 decap_w0
xfeed_10650 0 1 decap_w0
xfeed_9299 0 1 decap_w0
xfeed_9298 0 1 decap_w0
xfeed_9297 0 1 decap_w0
xfeed_9296 0 1 tie
xfeed_9295 0 1 decap_w0
xfeed_9294 0 1 decap_w0
xfeed_9293 0 1 decap_w0
xfeed_9291 0 1 decap_w0
xfeed_9290 0 1 decap_w0
xfeed_8761 0 1 decap_w0
xfeed_8760 0 1 decap_w0
xfeed_4459 0 1 decap_w0
xfeed_4458 0 1 decap_w0
xfeed_4457 0 1 decap_w0
xfeed_4456 0 1 decap_w0
xfeed_4455 0 1 decap_w0
xfeed_4454 0 1 decap_w0
xfeed_4453 0 1 decap_w0
xfeed_4452 0 1 decap_w0
xfeed_4451 0 1 decap_w0
xfeed_4450 0 1 decap_w0
xfeed_3922 0 1 decap_w0
xfeed_3921 0 1 decap_w0
xfeed_3920 0 1 tie
xsubckt_888_nexor2_x0 0 1 1598 1964 2055 nexor2_x0
xsubckt_884_mux2_x1 0 1 1600 1601 2000 445 mux2_x1
xsubckt_1375_or2_x1 0 1 1215 694 1323 or2_x1
xfeed_11190 0 1 tie
xfeed_8769 0 1 decap_w0
xfeed_8768 0 1 decap_w0
xfeed_8767 0 1 decap_w0
xfeed_8766 0 1 decap_w0
xfeed_8764 0 1 tie
xfeed_8763 0 1 decap_w0
xfeed_8762 0 1 decap_w0
xfeed_3929 0 1 decap_w0
xfeed_3928 0 1 decap_w0
xfeed_3927 0 1 decap_w0
xfeed_3926 0 1 decap_w0
xfeed_3925 0 1 decap_w0
xfeed_3924 0 1 decap_w0
xfeed_3923 0 1 decap_w0
xsubckt_52_inv_x0 0 1 730 2074 inv_x0
xsubckt_50_inv_x0 0 1 732 1980 inv_x0
xsubckt_331_nand2_x0 0 1 417 617 418 nand2_x0
xsubckt_459_nor3_x0 0 1 291 298 293 292 nor3_x0
xsubckt_501_and21nor_x0 0 1 250 251 400 557 and21nor_x0
xsubckt_530_and4_x1 0 1 223 365 364 342 341 and4_x1
xsubckt_1710_or21nand_x0 0 1 884 886 887 1075 or21nand_x0
xfeed_11199 0 1 decap_w0
xfeed_11198 0 1 decap_w0
xfeed_11197 0 1 decap_w0
xfeed_11196 0 1 decap_w0
xfeed_11195 0 1 decap_w0
xfeed_11194 0 1 decap_w0
xfeed_11193 0 1 decap_w0
xfeed_11192 0 1 decap_w0
xfeed_11191 0 1 decap_w0
xfeed_10669 0 1 decap_w0
xfeed_10668 0 1 decap_w0
xfeed_10667 0 1 decap_w0
xfeed_10666 0 1 decap_w0
xfeed_10665 0 1 decap_w0
xfeed_10664 0 1 decap_w0
xfeed_10663 0 1 decap_w0
xfeed_10662 0 1 decap_w0
xfeed_10661 0 1 decap_w0
xfeed_10660 0 1 decap_w0
xfeed_4468 0 1 decap_w0
xfeed_4467 0 1 decap_w0
xfeed_4466 0 1 decap_w0
xfeed_4465 0 1 decap_w0
xfeed_4464 0 1 decap_w0
xfeed_4463 0 1 decap_w0
xfeed_4462 0 1 decap_w0
xfeed_4461 0 1 decap_w0
xfeed_4460 0 1 decap_w0
xsubckt_948_nand2_x0 0 1 1571 1959 1575 nand2_x0
xsubckt_58_inv_x0 0 1 724 1946 inv_x0
xsubckt_56_inv_x0 0 1 726 1975 inv_x0
xsubckt_54_inv_x0 0 1 728 1977 inv_x0
xsubckt_151_nand2_x0 0 1 614 712 1926 nand2_x0
xsubckt_526_and4_x1 0 1 226 396 231 230 227 and4_x1
xfeed_8779 0 1 decap_w0
xfeed_8778 0 1 decap_w0
xfeed_8777 0 1 decap_w0
xfeed_8776 0 1 tie
xfeed_8775 0 1 decap_w0
xfeed_8774 0 1 decap_w0
xfeed_8773 0 1 decap_w0
xfeed_8772 0 1 decap_w0
xfeed_8771 0 1 decap_w0
xfeed_8770 0 1 decap_w0
xfeed_4469 0 1 decap_w0
xfeed_3939 0 1 decap_w0
xfeed_3938 0 1 tie
xfeed_3937 0 1 decap_w0
xfeed_3936 0 1 decap_w0
xfeed_3935 0 1 decap_w0
xfeed_3934 0 1 decap_w0
xfeed_3933 0 1 decap_w0
xfeed_3932 0 1 decap_w0
xfeed_3931 0 1 decap_w0
xfeed_3930 0 1 decap_w0
xsubckt_858_nand2_x0 0 1 1623 1946 1625 nand2_x0
xsubckt_768_nand2_x0 0 1 1701 1998 1746 nand2_x0
xsubckt_237_nand3_x0 0 1 514 616 594 556 nand3_x0
xsubckt_1362_nand2_x0 0 1 1227 2052 479 nand2_x0
xsubckt_1452_nand2_x0 0 1 1144 775 2056 nand2_x0
xsubckt_1685_nor2_x0 0 1 909 912 911 nor2_x0
xfeed_10679 0 1 decap_w0
xfeed_10678 0 1 decap_w0
xfeed_10677 0 1 decap_w0
xfeed_10676 0 1 decap_w0
xfeed_10675 0 1 decap_w0
xfeed_10674 0 1 decap_w0
xfeed_10673 0 1 decap_w0
xfeed_10672 0 1 decap_w0
xfeed_10671 0 1 decap_w0
xfeed_10670 0 1 decap_w0
xfeed_4475 0 1 decap_w0
xfeed_4474 0 1 decap_w0
xfeed_4473 0 1 decap_w0
xfeed_4472 0 1 decap_w0
xfeed_4471 0 1 tie
xfeed_4470 0 1 decap_w0
xsubckt_1272_nand2_x0 0 1 1309 774 1981 nand2_x0
xsubckt_1557_mux2_x1 0 1 1037 1109 1039 1142 mux2_x1
xsubckt_1663_and21nor_x0 0 1 931 932 1117 2051 and21nor_x0
xcmpt_abc_11867_new_n522_hfns_0 0 1 558 555 buf_x4
xcmpt_abc_11867_new_n522_hfns_1 0 1 557 555 buf_x4
xcmpt_abc_11867_new_n522_hfns_2 0 1 556 555 buf_x4
xcmpt_abc_11867_new_n522_hfns_3 0 1 555 559 buf_x4
xfeed_8789 0 1 decap_w0
xfeed_8788 0 1 decap_w0
xfeed_8787 0 1 decap_w0
xfeed_8786 0 1 tie
xfeed_8785 0 1 decap_w0
xfeed_8784 0 1 decap_w0
xfeed_8783 0 1 decap_w0
xfeed_8782 0 1 decap_w0
xfeed_8781 0 1 decap_w0
xfeed_8780 0 1 decap_w0
xfeed_4479 0 1 decap_w0
xfeed_4478 0 1 tie
xfeed_4477 0 1 decap_w0
xfeed_4476 0 1 decap_w0
xfeed_3949 0 1 decap_w0
xfeed_3948 0 1 decap_w0
xfeed_3947 0 1 decap_w0
xfeed_3946 0 1 decap_w0
xfeed_3945 0 1 decap_w0
xfeed_3944 0 1 decap_w0
xfeed_3943 0 1 decap_w0
xfeed_3942 0 1 decap_w0
xfeed_3941 0 1 decap_w0
xfeed_3940 0 1 decap_w0
xsubckt_1182_nand2_x0 0 1 1832 1385 1381 nand2_x0
xsubckt_1611_nand3_x0 0 1 983 1103 989 987 nand3_x0
xfeed_10689 0 1 decap_w0
xfeed_10688 0 1 decap_w0
xfeed_10687 0 1 decap_w0
xfeed_10686 0 1 decap_w0
xfeed_10685 0 1 decap_w0
xfeed_10684 0 1 tie
xfeed_10683 0 1 decap_w0
xfeed_10682 0 1 decap_w0
xfeed_10681 0 1 decap_w0
xfeed_10680 0 1 decap_w0
xfeed_9409 0 1 decap_w0
xfeed_9408 0 1 decap_w0
xfeed_9407 0 1 decap_w0
xfeed_9406 0 1 decap_w0
xfeed_9405 0 1 decap_w0
xfeed_9404 0 1 decap_w0
xfeed_9403 0 1 decap_w0
xfeed_9402 0 1 decap_w0
xfeed_9401 0 1 decap_w0
xfeed_4482 0 1 decap_w0
xfeed_4481 0 1 decap_w0
xfeed_4480 0 1 decap_w0
xsubckt_927_nand3_x0 0 1 1578 184 176 1620 nand3_x0
xsubckt_342_and4_x1 0 1 406 419 416 409 407 and4_x1
xsubckt_482_and2_x1 0 1 268 575 558 and2_x1
xsubckt_1431_nand3_x0 0 1 1163 2067 666 657 nand3_x0
xsubckt_1607_nand4_x0 0 1 987 1999 1128 1098 1097 nand4_x0
xsubckt_1634_and4_x1 0 1 960 2000 1128 1098 1097 and4_x1
xsubckt_1748_and3_x1 0 1 846 853 850 847 and3_x1
xfeed_11309 0 1 tie
xfeed_11308 0 1 decap_w0
xfeed_11307 0 1 decap_w0
xfeed_11306 0 1 decap_w0
xfeed_11305 0 1 decap_w0
xfeed_11304 0 1 decap_w0
xfeed_11303 0 1 decap_w0
xfeed_11302 0 1 decap_w0
xfeed_11301 0 1 decap_w0
xfeed_11300 0 1 decap_w0
xfeed_8799 0 1 decap_w0
xfeed_8798 0 1 decap_w0
xfeed_8797 0 1 decap_w0
xfeed_8796 0 1 tie
xfeed_8795 0 1 decap_w0
xfeed_8794 0 1 decap_w0
xfeed_8793 0 1 decap_w0
xfeed_8792 0 1 decap_w0
xfeed_8791 0 1 tie
xfeed_8790 0 1 decap_w0
xfeed_4489 0 1 decap_w0
xfeed_4488 0 1 decap_w0
xfeed_4487 0 1 decap_w0
xfeed_4486 0 1 decap_w0
xfeed_4485 0 1 decap_w0
xfeed_4484 0 1 decap_w0
xfeed_4483 0 1 decap_w0
xfeed_3959 0 1 decap_w0
xfeed_3958 0 1 decap_w0
xfeed_3957 0 1 decap_w0
xfeed_3956 0 1 decap_w0
xfeed_3955 0 1 decap_w0
xfeed_3954 0 1 decap_w0
xfeed_3953 0 1 decap_w0
xfeed_3952 0 1 decap_w0
xfeed_3951 0 1 tie
xfeed_3950 0 1 decap_w0
xsubckt_126_nand4_x0 0 1 642 660 651 648 647 nand4_x0
xsubckt_571_nand2_x0 0 1 184 187 185 nand2_x0
xsubckt_1559_and21nor_x0 0 1 1035 1070 1047 1073 and21nor_x0
xcmpt_abc_11867_new_n488_hfns_0 0 1 595 593 buf_x4
xcmpt_abc_11867_new_n488_hfns_1 0 1 594 593 buf_x4
xcmpt_abc_11867_new_n488_hfns_2 0 1 593 596 buf_x4
xfeed_10699 0 1 decap_w0
xfeed_10698 0 1 decap_w0
xfeed_10697 0 1 decap_w0
xfeed_10696 0 1 decap_w0
xfeed_10695 0 1 decap_w0
xfeed_10694 0 1 decap_w0
xfeed_10693 0 1 decap_w0
xfeed_10692 0 1 decap_w0
xfeed_10691 0 1 tie
xfeed_10690 0 1 decap_w0
xfeed_9419 0 1 decap_w0
xfeed_9418 0 1 decap_w0
xfeed_9417 0 1 decap_w0
xfeed_9416 0 1 decap_w0
xfeed_9415 0 1 decap_w0
xfeed_9414 0 1 decap_w0
xfeed_9413 0 1 decap_w0
xfeed_9412 0 1 decap_w0
xfeed_9411 0 1 decap_w0
xfeed_9410 0 1 decap_w0
xfeed_5109 0 1 decap_w0
xfeed_5108 0 1 decap_w0
xfeed_5107 0 1 decap_w0
xfeed_5106 0 1 decap_w0
xfeed_5105 0 1 decap_w0
xfeed_5104 0 1 decap_w0
xfeed_5103 0 1 tie
xfeed_5102 0 1 decap_w0
xfeed_5101 0 1 decap_w0
xfeed_5100 0 1 decap_w0
xsubckt_793_and21nor_x0 0 1 1679 1680 1740 2053 and21nor_x0
xsubckt_657_nand3_x0 0 1 103 2016 184 177 nand3_x0
xsubckt_312_and2_x1 0 1 436 681 447 and2_x1
xsubckt_303_nand2_x0 0 1 445 616 447 nand2_x0
xsubckt_1818_mux2_x1 0 1 1787 2057 1109 775 mux2_x1
xfeed_11316 0 1 decap_w0
xfeed_11315 0 1 decap_w0
xfeed_11314 0 1 tie
xfeed_11313 0 1 decap_w0
xfeed_11312 0 1 decap_w0
xfeed_11311 0 1 decap_w0
xfeed_11310 0 1 decap_w0
xfeed_4499 0 1 decap_w0
xfeed_4498 0 1 decap_w0
xfeed_4497 0 1 decap_w0
xfeed_4496 0 1 decap_w0
xfeed_4495 0 1 decap_w0
xfeed_4494 0 1 decap_w0
xfeed_4493 0 1 decap_w0
xfeed_4492 0 1 decap_w0
xfeed_4491 0 1 decap_w0
xfeed_3969 0 1 decap_w0
xfeed_3968 0 1 decap_w0
xfeed_3967 0 1 decap_w0
xfeed_3966 0 1 decap_w0
xfeed_3964 0 1 decap_w0
xfeed_3963 0 1 decap_w0
xfeed_3962 0 1 decap_w0
xfeed_3960 0 1 decap_w0
xsubckt_736_or21nand_x0 0 1 1729 2064 1742 1740 or21nand_x0
xsubckt_391_nand2_x0 0 1 358 533 360 nand2_x0
xsubckt_1297_or21nand_x0 0 1 1286 1287 1322 764 or21nand_x0
xfeed_11319 0 1 decap_w0
xfeed_11318 0 1 decap_w0
xfeed_9429 0 1 decap_w0
xfeed_9428 0 1 decap_w0
xfeed_9427 0 1 decap_w0
xfeed_9426 0 1 decap_w0
xfeed_9425 0 1 decap_w0
xfeed_9424 0 1 decap_w0
xfeed_9423 0 1 decap_w0
xfeed_9422 0 1 decap_w0
xfeed_9421 0 1 decap_w0
xfeed_9420 0 1 decap_w0
xfeed_5119 0 1 decap_w0
xfeed_5118 0 1 decap_w0
xfeed_5117 0 1 tie
xfeed_5116 0 1 decap_w0
xfeed_5115 0 1 decap_w0
xfeed_5114 0 1 decap_w0
xfeed_5113 0 1 decap_w0
xfeed_5112 0 1 decap_w0
xfeed_5111 0 1 decap_w0
xfeed_5110 0 1 tie
xsubckt_1155_and2_x1 0 1 1405 1409 1406 and2_x1
xsubckt_743_and2_x1 0 1 1723 2051 1748 and2_x1
xsubckt_308_and2_x1 0 1 440 442 441 and2_x1
xsubckt_293_or2_x1 0 1 455 684 456 or2_x1
xsubckt_209_nand3_x0 0 1 545 617 612 558 nand3_x0
xsubckt_603_and4_x1 0 1 153 157 156 155 154 and4_x1
xsubckt_1334_nand2_x0 0 1 1253 773 1969 nand2_x0
xfeed_11323 0 1 decap_w0
xfeed_11322 0 1 decap_w0
xfeed_11321 0 1 decap_w0
xfeed_11320 0 1 decap_w0
xfeed_3979 0 1 tie
xfeed_3978 0 1 decap_w0
xfeed_3977 0 1 decap_w0
xfeed_3976 0 1 decap_w0
xfeed_3975 0 1 decap_w0
xfeed_3974 0 1 decap_w0
xfeed_3973 0 1 decap_w0
xfeed_3972 0 1 tie
xfeed_3971 0 1 decap_w0
xfeed_3970 0 1 decap_w0
xsubckt_492_and21nor_x0 0 1 259 260 297 535 and21nor_x0
xsubckt_1505_or21nand_x0 0 1 1091 1105 1100 1096 or21nand_x0
xsubckt_1512_and2_x1 0 1 1084 1125 1085 and2_x1
xsubckt_1598_nand3_x0 0 1 996 1005 1001 999 nand3_x0
xsubckt_1759_and21nor_x0 0 1 835 908 839 837 and21nor_x0
xfeed_11329 0 1 decap_w0
xfeed_11328 0 1 decap_w0
xfeed_11327 0 1 decap_w0
xfeed_11326 0 1 decap_w0
xfeed_11325 0 1 decap_w0
xfeed_11324 0 1 decap_w0
xfeed_9439 0 1 decap_w0
xfeed_9438 0 1 decap_w0
xfeed_9437 0 1 decap_w0
xfeed_9436 0 1 decap_w0
xfeed_9435 0 1 decap_w0
xfeed_9434 0 1 decap_w0
xfeed_9433 0 1 decap_w0
xfeed_9432 0 1 decap_w0
xfeed_9431 0 1 decap_w0
xfeed_9430 0 1 decap_w0
xfeed_8901 0 1 decap_w0
xfeed_8900 0 1 decap_w0
xfeed_5129 0 1 tie
xfeed_5128 0 1 decap_w0
xfeed_5127 0 1 decap_w0
xfeed_5126 0 1 decap_w0
xfeed_5125 0 1 decap_w0
xfeed_5124 0 1 tie
xfeed_5123 0 1 decap_w0
xfeed_5122 0 1 decap_w0
xfeed_5121 0 1 decap_w0
xfeed_5120 0 1 decap_w0
xsubckt_993_and21nor_x0 0 1 1535 623 312 1536 and21nor_x0
xsubckt_216_and2_x1 0 1 538 610 595 and2_x1
xsubckt_370_nand3_x0 0 1 379 532 530 382 nand3_x0
xsubckt_460_nand3_x0 0 1 290 309 304 291 nand3_x0
xsubckt_546_nand4_x0 0 1 208 449 410 325 210 nand4_x0
xsubckt_1472_and3_x1 0 1 1124 503 430 192 and3_x1
xfeed_11330 0 1 decap_w0
xfeed_8909 0 1 decap_w0
xfeed_8908 0 1 decap_w0
xfeed_8907 0 1 decap_w0
xfeed_8906 0 1 decap_w0
xfeed_8905 0 1 decap_w0
xfeed_8904 0 1 decap_w0
xfeed_8903 0 1 decap_w0
xfeed_8902 0 1 decap_w0
xfeed_3989 0 1 decap_w0
xfeed_3988 0 1 decap_w0
xfeed_3987 0 1 decap_w0
xfeed_3986 0 1 decap_w0
xfeed_3985 0 1 decap_w0
xfeed_3984 0 1 decap_w0
xfeed_3983 0 1 decap_w0
xfeed_3982 0 1 decap_w0
xfeed_3981 0 1 decap_w0
xfeed_3980 0 1 decap_w0
xsubckt_1050_nand4_x0 0 1 1490 623 525 519 1576 nand4_x0
xsubckt_456_nand4_x0 0 1 294 533 530 524 383 nand4_x0
xsubckt_1420_and2_x1 0 1 1173 1177 1174 and2_x1
xsubckt_1468_and3_x1 0 1 1128 503 482 1340 and3_x1
xsubckt_1494_and2_x1 0 1 1102 1105 1103 and2_x1
xfeed_11339 0 1 decap_w0
xfeed_11338 0 1 decap_w0
xfeed_11337 0 1 decap_w0
xfeed_11336 0 1 decap_w0
xfeed_11335 0 1 decap_w0
xfeed_11334 0 1 decap_w0
xfeed_11333 0 1 decap_w0
xfeed_11332 0 1 decap_w0
xfeed_11331 0 1 tie
xfeed_10809 0 1 decap_w0
xfeed_10808 0 1 decap_w0
xfeed_10807 0 1 decap_w0
xfeed_10806 0 1 decap_w0
xfeed_10805 0 1 decap_w0
xfeed_10804 0 1 tie
xfeed_10803 0 1 decap_w0
xfeed_10802 0 1 decap_w0
xfeed_10801 0 1 decap_w0
xfeed_10800 0 1 decap_w0
xfeed_9447 0 1 decap_w0
xfeed_9446 0 1 decap_w0
xfeed_9445 0 1 decap_w0
xfeed_9444 0 1 decap_w0
xfeed_9443 0 1 decap_w0
xfeed_9442 0 1 tie
xfeed_9441 0 1 decap_w0
xfeed_9440 0 1 decap_w0
xfeed_5139 0 1 decap_w0
xfeed_5138 0 1 decap_w0
xfeed_5137 0 1 decap_w0
xfeed_5136 0 1 decap_w0
xfeed_5135 0 1 decap_w0
xfeed_5134 0 1 decap_w0
xfeed_5133 0 1 decap_w0
xfeed_5132 0 1 decap_w0
xfeed_5131 0 1 decap_w0
xfeed_5130 0 1 decap_w0
xfeed_4608 0 1 decap_w0
xfeed_4607 0 1 decap_w0
xfeed_4606 0 1 decap_w0
xfeed_4605 0 1 decap_w0
xfeed_4604 0 1 decap_w0
xfeed_4603 0 1 decap_w0
xfeed_4602 0 1 decap_w0
xfeed_4601 0 1 decap_w0
xfeed_4600 0 1 decap_w0
xfeed_9449 0 1 decap_w0
xfeed_9448 0 1 decap_w0
xfeed_8919 0 1 decap_w0
xfeed_8918 0 1 decap_w0
xfeed_8917 0 1 decap_w0
xfeed_8916 0 1 tie
xfeed_8915 0 1 decap_w0
xfeed_8914 0 1 decap_w0
xfeed_8913 0 1 decap_w0
xfeed_8912 0 1 decap_w0
xfeed_8911 0 1 decap_w0
xfeed_8910 0 1 decap_w0
xfeed_4609 0 1 decap_w0
xfeed_3999 0 1 decap_w0
xfeed_3998 0 1 tie
xfeed_3997 0 1 decap_w0
xfeed_3996 0 1 decap_w0
xfeed_3995 0 1 decap_w0
xfeed_3994 0 1 decap_w0
xfeed_3993 0 1 decap_w0
xfeed_3992 0 1 decap_w0
xfeed_3991 0 1 tie
xfeed_3990 0 1 decap_w0
xsubckt_1196_or21nand_x0 0 1 1368 680 490 447 or21nand_x0
xsubckt_1128_nexor2_x0 0 1 1429 2055 1430 nexor2_x0
xsubckt_800_and21nor_x0 0 1 1673 695 1755 1754 and21nor_x0
xsubckt_555_and2_x1 0 1 200 505 438 and2_x1
xfeed_11349 0 1 decap_w0
xfeed_11348 0 1 decap_w0
xfeed_11347 0 1 decap_w0
xfeed_11346 0 1 decap_w0
xfeed_11345 0 1 decap_w0
xfeed_11344 0 1 decap_w0
xfeed_11343 0 1 decap_w0
xfeed_11342 0 1 decap_w0
xfeed_11341 0 1 decap_w0
xfeed_11340 0 1 tie
xfeed_10819 0 1 decap_w0
xfeed_10817 0 1 decap_w0
xfeed_10816 0 1 tie
xfeed_10815 0 1 decap_w0
xfeed_10814 0 1 decap_w0
xfeed_10813 0 1 decap_w0
xfeed_10812 0 1 decap_w0
xfeed_10811 0 1 decap_w0
xfeed_10810 0 1 decap_w0
xfeed_9454 0 1 decap_w0
xfeed_9453 0 1 decap_w0
xfeed_9452 0 1 decap_w0
xfeed_9451 0 1 decap_w0
xfeed_5149 0 1 decap_w0
xfeed_5148 0 1 decap_w0
xfeed_5147 0 1 decap_w0
xfeed_5146 0 1 tie
xfeed_5145 0 1 decap_w0
xfeed_5144 0 1 decap_w0
xfeed_5143 0 1 decap_w0
xfeed_5142 0 1 tie
xfeed_5141 0 1 decap_w0
xfeed_4615 0 1 decap_w0
xfeed_4614 0 1 decap_w0
xfeed_4613 0 1 decap_w0
xfeed_4612 0 1 tie
xfeed_4611 0 1 decap_w0
xfeed_4610 0 1 decap_w0
xsubckt_1219_nand4_x0 0 1 1345 1928 1925 711 589 nand4_x0
xsubckt_1043_nand3_x0 0 1 1495 623 526 519 nand3_x0
xsubckt_792_and21nor_x0 0 1 1680 747 600 1745 and21nor_x0
xfeed_9459 0 1 tie
xfeed_9458 0 1 decap_w0
xfeed_9457 0 1 decap_w0
xfeed_9456 0 1 decap_w0
xfeed_9455 0 1 decap_w0
xfeed_8929 0 1 decap_w0
xfeed_8928 0 1 decap_w0
xfeed_8927 0 1 decap_w0
xfeed_8926 0 1 decap_w0
xfeed_8925 0 1 decap_w0
xfeed_8924 0 1 decap_w0
xfeed_8923 0 1 tie
xfeed_8922 0 1 decap_w0
xfeed_8921 0 1 decap_w0
xfeed_8920 0 1 decap_w0
xfeed_4619 0 1 decap_w0
xfeed_4618 0 1 decap_w0
xfeed_4617 0 1 decap_w0
xfeed_4616 0 1 decap_w0
xsubckt_1258_and4_x1 0 1 1322 605 493 476 1756 and4_x1
xsubckt_1170_and4_x1 0 1 1392 778 678 674 670 and4_x1
xsubckt_1039_nand4_x0 0 1 1498 637 633 1563 1515 nand4_x0
xsubckt_872_and3_x1 0 1 1611 1962 1964 2054 and3_x1
xsubckt_790_nand3_x0 0 1 1682 2073 678 489 nand3_x0
xsubckt_612_nand3_x0 0 1 145 2027 184 176 nand3_x0
xfeed_11359 0 1 decap_w0
xfeed_11358 0 1 decap_w0
xfeed_11357 0 1 decap_w0
xfeed_11356 0 1 decap_w0
xfeed_11355 0 1 decap_w0
xfeed_11354 0 1 decap_w0
xfeed_11353 0 1 decap_w0
xfeed_11352 0 1 decap_w0
xfeed_11351 0 1 decap_w0
xfeed_11350 0 1 decap_w0
xfeed_10829 0 1 decap_w0
xfeed_10828 0 1 decap_w0
xfeed_10827 0 1 decap_w0
xfeed_10826 0 1 tie
xfeed_10825 0 1 decap_w0
xfeed_10823 0 1 decap_w0
xfeed_10822 0 1 decap_w0
xfeed_10821 0 1 decap_w0
xfeed_10820 0 1 decap_w0
xfeed_9461 0 1 decap_w0
xfeed_9460 0 1 decap_w0
xfeed_5159 0 1 decap_w0
xfeed_5158 0 1 decap_w0
xfeed_5157 0 1 decap_w0
xfeed_5156 0 1 decap_w0
xfeed_5155 0 1 decap_w0
xfeed_5154 0 1 decap_w0
xfeed_5153 0 1 decap_w0
xfeed_5152 0 1 decap_w0
xfeed_5151 0 1 decap_w0
xfeed_5150 0 1 decap_w0
xfeed_4622 0 1 decap_w0
xfeed_4621 0 1 decap_w0
xfeed_4620 0 1 decap_w0
xsubckt_1820_dff_x1 0 1 2020 1912 35 dff_x1
xsubckt_1822_dff_x1 0 1 2018 1910 32 dff_x1
xsubckt_1824_dff_x1 0 1 2016 1908 32 dff_x1
xfeed_9469 0 1 decap_w0
xfeed_9468 0 1 decap_w0
xfeed_9467 0 1 decap_w0
xfeed_9466 0 1 tie
xfeed_9465 0 1 decap_w0
xfeed_9464 0 1 decap_w0
xfeed_9463 0 1 decap_w0
xfeed_9462 0 1 decap_w0
xfeed_8939 0 1 decap_w0
xfeed_8938 0 1 decap_w0
xfeed_8937 0 1 decap_w0
xfeed_8936 0 1 decap_w0
xfeed_8935 0 1 tie
xfeed_8934 0 1 decap_w0
xfeed_8933 0 1 decap_w0
xfeed_8932 0 1 decap_w0
xfeed_8931 0 1 decap_w0
xfeed_8930 0 1 tie
xfeed_4629 0 1 decap_w0
xfeed_4628 0 1 decap_w0
xfeed_4627 0 1 decap_w0
xfeed_4626 0 1 decap_w0
xfeed_4625 0 1 decap_w0
xfeed_4624 0 1 tie
xfeed_4623 0 1 decap_w0
xsubckt_432_nand3_x0 0 1 28 373 336 318 nand3_x0
xsubckt_635_nor2_x0 0 1 123 125 124 nor2_x0
xsubckt_1826_dff_x1 0 1 2014 1906 32 dff_x1
xsubckt_1828_dff_x1 0 1 1929 28 74 dff_x1
xfeed_11369 0 1 decap_w0
xfeed_11368 0 1 decap_w0
xfeed_11367 0 1 decap_w0
xfeed_11366 0 1 decap_w0
xfeed_11365 0 1 decap_w0
xfeed_11364 0 1 decap_w0
xfeed_11363 0 1 decap_w0
xfeed_11362 0 1 decap_w0
xfeed_11361 0 1 decap_w0
xfeed_11360 0 1 decap_w0
xfeed_10839 0 1 decap_w0
xfeed_10838 0 1 decap_w0
xfeed_10837 0 1 decap_w0
xfeed_10836 0 1 decap_w0
xfeed_10835 0 1 decap_w0
xfeed_10834 0 1 decap_w0
xfeed_10833 0 1 tie
xfeed_10832 0 1 decap_w0
xfeed_10831 0 1 decap_w0
xfeed_10830 0 1 decap_w0
xfeed_5168 0 1 tie
xfeed_5167 0 1 decap_w0
xfeed_5166 0 1 decap_w0
xfeed_5165 0 1 decap_w0
xfeed_5164 0 1 decap_w0
xfeed_5163 0 1 decap_w0
xfeed_5162 0 1 decap_w0
xfeed_5161 0 1 tie
xfeed_5160 0 1 decap_w0
xsubckt_963_nand2_x0 0 1 1560 1957 1575 nand2_x0
xfeed_9479 0 1 decap_w0
xfeed_9478 0 1 decap_w0
xfeed_9477 0 1 decap_w0
xfeed_9476 0 1 decap_w0
xfeed_9475 0 1 decap_w0
xfeed_9474 0 1 decap_w0
xfeed_9473 0 1 decap_w0
xfeed_9472 0 1 decap_w0
xfeed_9471 0 1 decap_w0
xfeed_9470 0 1 decap_w0
xfeed_8949 0 1 decap_w0
xfeed_8948 0 1 decap_w0
xfeed_8947 0 1 tie
xfeed_8946 0 1 decap_w0
xfeed_8945 0 1 decap_w0
xfeed_8944 0 1 decap_w0
xfeed_8943 0 1 decap_w0
xfeed_8941 0 1 decap_w0
xfeed_8940 0 1 decap_w0
xfeed_5169 0 1 decap_w0
xfeed_4639 0 1 decap_w0
xfeed_4638 0 1 decap_w0
xfeed_4637 0 1 decap_w0
xfeed_4636 0 1 decap_w0
xfeed_4635 0 1 tie
xfeed_4634 0 1 decap_w0
xfeed_4633 0 1 decap_w0
xfeed_4632 0 1 decap_w0
xfeed_4631 0 1 tie
xsubckt_1095_or21nand_x0 0 1 1452 1492 312 642 or21nand_x0
xsubckt_938_mux2_x1 0 1 1880 1954 526 774 mux2_x1
xfeed_11379 0 1 decap_w0
xfeed_11378 0 1 decap_w0
xfeed_11377 0 1 decap_w0
xfeed_11376 0 1 decap_w0
xfeed_11375 0 1 decap_w0
xfeed_11374 0 1 decap_w0
xfeed_11373 0 1 decap_w0
xfeed_11372 0 1 decap_w0
xfeed_11371 0 1 decap_w0
xfeed_11370 0 1 decap_w0
xfeed_10849 0 1 decap_w0
xfeed_10848 0 1 decap_w0
xfeed_10847 0 1 decap_w0
xfeed_10846 0 1 decap_w0
xfeed_10845 0 1 decap_w0
xfeed_10844 0 1 decap_w0
xfeed_10843 0 1 decap_w0
xfeed_10842 0 1 decap_w0
xfeed_10841 0 1 decap_w0
xfeed_10840 0 1 decap_w0
xfeed_5175 0 1 decap_w0
xfeed_5174 0 1 decap_w0
xfeed_5173 0 1 decap_w0
xfeed_5172 0 1 decap_w0
xfeed_5171 0 1 decap_w0
xfeed_5170 0 1 decap_w0
xsubckt_610_and3_x1 0 1 146 151 150 147 and3_x1
xsubckt_1707_mux2_x1 0 1 887 929 889 1142 mux2_x1
xfeed_9489 0 1 decap_w0
xfeed_9488 0 1 decap_w0
xfeed_9487 0 1 decap_w0
xfeed_9486 0 1 decap_w0
xfeed_9485 0 1 decap_w0
xfeed_9484 0 1 decap_w0
xfeed_9483 0 1 decap_w0
xfeed_9482 0 1 decap_w0
xfeed_9481 0 1 decap_w0
xfeed_9480 0 1 decap_w0
xfeed_8959 0 1 decap_w0
xfeed_8958 0 1 decap_w0
xfeed_8957 0 1 decap_w0
xfeed_8956 0 1 decap_w0
xfeed_8954 0 1 tie
xfeed_8953 0 1 decap_w0
xfeed_8952 0 1 decap_w0
xfeed_8951 0 1 decap_w0
xfeed_8950 0 1 decap_w0
xfeed_5179 0 1 decap_w0
xfeed_5178 0 1 decap_w0
xfeed_5177 0 1 decap_w0
xfeed_5176 0 1 decap_w0
xfeed_4649 0 1 tie
xfeed_4648 0 1 decap_w0
xfeed_4647 0 1 decap_w0
xfeed_4646 0 1 decap_w0
xfeed_4645 0 1 decap_w0
xfeed_4644 0 1 decap_w0
xfeed_4643 0 1 decap_w0
xfeed_4642 0 1 tie
xfeed_4640 0 1 decap_w0
xsubckt_691_and21nor_x0 0 1 1772 748 449 410 and21nor_x0
xsubckt_404_nexor2_x0 0 1 345 757 346 nexor2_x0
xsubckt_599_nand3_x0 0 1 157 2028 184 176 nand3_x0
xsubckt_1308_nor2_x0 0 1 1276 1280 1277 nor2_x0
xsubckt_1615_mux2_x1 0 1 979 985 980 992 mux2_x1
xfeed_11389 0 1 decap_w0
xfeed_11388 0 1 decap_w0
xfeed_11387 0 1 decap_w0
xfeed_11386 0 1 decap_w0
xfeed_11385 0 1 decap_w0
xfeed_11384 0 1 decap_w0
xfeed_11383 0 1 decap_w0
xfeed_11382 0 1 decap_w0
xfeed_11381 0 1 decap_w0
xfeed_11380 0 1 decap_w0
xfeed_10859 0 1 decap_w0
xfeed_10858 0 1 decap_w0
xfeed_10857 0 1 decap_w0
xfeed_10856 0 1 decap_w0
xfeed_10855 0 1 decap_w0
xfeed_10854 0 1 decap_w0
xfeed_10853 0 1 decap_w0
xfeed_10852 0 1 decap_w0
xfeed_10851 0 1 decap_w0
xfeed_10850 0 1 decap_w0
xfeed_5182 0 1 decap_w0
xfeed_5181 0 1 decap_w0
xfeed_5180 0 1 decap_w0
xsubckt_65_inv_x0 0 1 717 2085 inv_x0
xsubckt_63_inv_x0 0 1 719 2084 inv_x0
xsubckt_61_inv_x0 0 1 721 2083 inv_x0
xfeed_12009 0 1 decap_w0
xfeed_12008 0 1 decap_w0
xfeed_12007 0 1 decap_w0
xfeed_12006 0 1 decap_w0
xfeed_12005 0 1 decap_w0
xfeed_12004 0 1 decap_w0
xfeed_12003 0 1 decap_w0
xfeed_12002 0 1 decap_w0
xfeed_12001 0 1 decap_w0
xfeed_12000 0 1 tie
xfeed_9499 0 1 decap_w0
xfeed_9498 0 1 decap_w0
xfeed_9497 0 1 decap_w0
xfeed_9496 0 1 decap_w0
xfeed_9495 0 1 decap_w0
xfeed_9494 0 1 decap_w0
xfeed_9493 0 1 decap_w0
xfeed_9492 0 1 decap_w0
xfeed_9491 0 1 decap_w0
xfeed_9490 0 1 decap_w0
xfeed_8969 0 1 decap_w0
xfeed_8968 0 1 decap_w0
xfeed_8967 0 1 decap_w0
xfeed_8966 0 1 decap_w0
xfeed_8964 0 1 decap_w0
xfeed_8963 0 1 decap_w0
xfeed_8962 0 1 decap_w0
xfeed_8961 0 1 tie
xfeed_8960 0 1 decap_w0
xfeed_5189 0 1 decap_w0
xfeed_5188 0 1 decap_w0
xfeed_5187 0 1 decap_w0
xfeed_5186 0 1 decap_w0
xfeed_5185 0 1 decap_w0
xfeed_5184 0 1 decap_w0
xfeed_5183 0 1 decap_w0
xfeed_4659 0 1 decap_w0
xfeed_4658 0 1 decap_w0
xfeed_4657 0 1 decap_w0
xfeed_4656 0 1 decap_w0
xfeed_4655 0 1 decap_w0
xfeed_4654 0 1 decap_w0
xfeed_4653 0 1 decap_w0
xfeed_4652 0 1 decap_w0
xfeed_4651 0 1 decap_w0
xfeed_4650 0 1 decap_w0
xsubckt_69_inv_x0 0 1 713 1928 inv_x0
xsubckt_67_inv_x0 0 1 715 1924 inv_x0
xsubckt_155_nand2_x0 0 1 606 1925 711 nand2_x0
xsubckt_514_and3_x1 0 1 237 412 406 328 and3_x1
xsubckt_592_and3_x1 0 1 163 735 608 460 and3_x1
xsubckt_1449_and3_x1 0 1 1146 1169 1159 1148 and3_x1
xfeed_11399 0 1 decap_w0
xfeed_11398 0 1 decap_w0
xfeed_11397 0 1 decap_w0
xfeed_11396 0 1 decap_w0
xfeed_11395 0 1 decap_w0
xfeed_11394 0 1 decap_w0
xfeed_11393 0 1 decap_w0
xfeed_11392 0 1 decap_w0
xfeed_11391 0 1 decap_w0
xfeed_11390 0 1 decap_w0
xfeed_10869 0 1 decap_w0
xfeed_10868 0 1 decap_w0
xfeed_10867 0 1 decap_w0
xfeed_10866 0 1 decap_w0
xfeed_10865 0 1 decap_w0
xfeed_10864 0 1 decap_w0
xfeed_10863 0 1 decap_w0
xfeed_10862 0 1 decap_w0
xfeed_10861 0 1 decap_w0
xfeed_10860 0 1 decap_w0
xsubckt_1276_nand2_x0 0 1 1305 1307 1306 nand2_x0
xsubckt_582_nand3_x0 0 1 173 2029 184 176 nand3_x0
xsubckt_588_and3_x1 0 1 167 1941 608 460 and3_x1
xfeed_12016 0 1 decap_w0
xfeed_12015 0 1 decap_w0
xfeed_12014 0 1 decap_w0
xfeed_12013 0 1 decap_w0
xfeed_12012 0 1 decap_w0
xfeed_12011 0 1 decap_w0
xfeed_12010 0 1 decap_w0
xfeed_8979 0 1 decap_w0
xfeed_8978 0 1 decap_w0
xfeed_8977 0 1 decap_w0
xfeed_8976 0 1 decap_w0
xfeed_8975 0 1 decap_w0
xfeed_8974 0 1 tie
xfeed_8973 0 1 decap_w0
xfeed_8972 0 1 decap_w0
xfeed_8971 0 1 decap_w0
xfeed_8970 0 1 decap_w0
xfeed_5199 0 1 decap_w0
xfeed_5198 0 1 decap_w0
xfeed_5197 0 1 decap_w0
xfeed_5196 0 1 decap_w0
xfeed_5195 0 1 decap_w0
xfeed_5194 0 1 decap_w0
xfeed_5193 0 1 decap_w0
xfeed_5192 0 1 decap_w0
xfeed_5191 0 1 decap_w0
xfeed_5190 0 1 decap_w0
xfeed_4669 0 1 tie
xfeed_4668 0 1 decap_w0
xfeed_4667 0 1 decap_w0
xfeed_4666 0 1 decap_w0
xfeed_4665 0 1 decap_w0
xfeed_4664 0 1 tie
xfeed_4663 0 1 decap_w0
xfeed_4662 0 1 decap_w0
xfeed_4661 0 1 decap_w0
xfeed_4660 0 1 decap_w0
xsubckt_314_nand3_x0 0 1 434 687 681 447 nand3_x0
xsubckt_536_and2_x1 0 1 217 246 218 and2_x1
xsubckt_1714_and3_x1 0 1 880 888 884 882 and3_x1
xfeed_12019 0 1 decap_w0
xfeed_12018 0 1 decap_w0
xfeed_12017 0 1 decap_w0
xfeed_10879 0 1 decap_w0
xfeed_10878 0 1 decap_w0
xfeed_10877 0 1 decap_w0
xfeed_10876 0 1 decap_w0
xfeed_10875 0 1 decap_w0
xfeed_10874 0 1 decap_w0
xfeed_10873 0 1 decap_w0
xfeed_10872 0 1 decap_w0
xfeed_10870 0 1 decap_w0
xsubckt_1096_nand2_x0 0 1 1451 1554 1452 nand2_x0
xsubckt_687_and21nor_x0 0 1 1776 206 1782 1778 and21nor_x0
xsubckt_620_nor2_x0 0 1 137 732 212 nor2_x0
xsubckt_1356_and21nor_x0 0 1 1232 775 1244 1235 and21nor_x0
xsubckt_1379_and2_x1 0 1 1211 1215 1212 and2_x1
xfeed_12023 0 1 decap_w0
xfeed_12022 0 1 decap_w0
xfeed_12021 0 1 decap_w0
xfeed_12020 0 1 tie
xfeed_8989 0 1 tie
xfeed_8988 0 1 decap_w0
xfeed_8987 0 1 decap_w0
xfeed_8986 0 1 decap_w0
xfeed_8985 0 1 decap_w0
xfeed_8984 0 1 decap_w0
xfeed_8983 0 1 decap_w0
xfeed_8982 0 1 decap_w0
xfeed_8981 0 1 decap_w0
xfeed_8980 0 1 decap_w0
xfeed_4679 0 1 decap_w0
xfeed_4678 0 1 decap_w0
xfeed_4677 0 1 decap_w0
xfeed_4676 0 1 decap_w0
xfeed_4675 0 1 decap_w0
xfeed_4674 0 1 decap_w0
xfeed_4673 0 1 decap_w0
xfeed_4672 0 1 decap_w0
xfeed_4671 0 1 decap_w0
xsubckt_330_and3_x1 0 1 418 1927 713 673 and3_x1
xfeed_12029 0 1 decap_w0
xfeed_12028 0 1 decap_w0
xfeed_12027 0 1 decap_w0
xfeed_12026 0 1 tie
xfeed_12025 0 1 decap_w0
xfeed_12024 0 1 decap_w0
xfeed_10889 0 1 decap_w0
xfeed_10888 0 1 decap_w0
xfeed_10887 0 1 decap_w0
xfeed_10886 0 1 decap_w0
xfeed_10885 0 1 tie
xfeed_10884 0 1 decap_w0
xfeed_10883 0 1 decap_w0
xfeed_10882 0 1 decap_w0
xfeed_10881 0 1 decap_w0
xfeed_10880 0 1 decap_w0
xfeed_9601 0 1 decap_w0
xfeed_9600 0 1 decap_w0
xsubckt_801_and2_x1 0 1 1672 2052 1740 and2_x1
xsubckt_378_and4_x1 0 1 371 643 622 532 384 and4_x1
xsubckt_1287_and2_x1 0 1 1295 1298 1296 and2_x1
xsubckt_1456_and21nor_x0 0 1 1140 755 547 1745 and21nor_x0
xfeed_12030 0 1 decap_w0
xfeed_9609 0 1 decap_w0
xfeed_9608 0 1 decap_w0
xfeed_9606 0 1 decap_w0
xfeed_9605 0 1 decap_w0
xfeed_9604 0 1 decap_w0
xfeed_9603 0 1 decap_w0
xfeed_9602 0 1 decap_w0
xfeed_8999 0 1 decap_w0
xfeed_8998 0 1 decap_w0
xfeed_8997 0 1 decap_w0
xfeed_8996 0 1 tie
xfeed_8995 0 1 decap_w0
xfeed_8994 0 1 decap_w0
xfeed_8993 0 1 decap_w0
xfeed_8992 0 1 decap_w0
xfeed_8991 0 1 decap_w0
xfeed_8990 0 1 decap_w0
xfeed_4689 0 1 decap_w0
xfeed_4688 0 1 decap_w0
xfeed_4687 0 1 decap_w0
xfeed_4686 0 1 decap_w0
xfeed_4685 0 1 decap_w0
xfeed_4684 0 1 decap_w0
xfeed_4683 0 1 decap_w0
xfeed_4682 0 1 decap_w0
xfeed_4681 0 1 decap_w0
xfeed_4680 0 1 decap_w0
xsubckt_1194_or21nand_x0 0 1 1370 501 487 614 or21nand_x0
xsubckt_923_mux2_x1 0 1 1893 1599 2033 1579 mux2_x1
xsubckt_217_nand2_x0 0 1 537 610 595 nand2_x0
xsubckt_203_nand4_x0 0 1 551 1925 711 673 669 nand4_x0
xsubckt_381_nand4_x0 0 1 368 652 638 632 530 nand4_x0
xfeed_12039 0 1 decap_w0
xfeed_12038 0 1 decap_w0
xfeed_12037 0 1 decap_w0
xfeed_12036 0 1 decap_w0
xfeed_12035 0 1 decap_w0
xfeed_12034 0 1 decap_w0
xfeed_12033 0 1 decap_w0
xfeed_12032 0 1 decap_w0
xfeed_12031 0 1 decap_w0
xfeed_11509 0 1 decap_w0
xfeed_11508 0 1 decap_w0
xfeed_11507 0 1 decap_w0
xfeed_11506 0 1 decap_w0
xfeed_11505 0 1 decap_w0
xfeed_11504 0 1 decap_w0
xfeed_11503 0 1 decap_w0
xfeed_11502 0 1 decap_w0
xfeed_11501 0 1 decap_w0
xfeed_11500 0 1 decap_w0
xfeed_10899 0 1 decap_w0
xfeed_10898 0 1 decap_w0
xfeed_10897 0 1 decap_w0
xfeed_10896 0 1 decap_w0
xfeed_10895 0 1 decap_w0
xfeed_10894 0 1 decap_w0
xfeed_10893 0 1 decap_w0
xfeed_10892 0 1 decap_w0
xfeed_10891 0 1 decap_w0
xfeed_10890 0 1 decap_w0
xfeed_5308 0 1 decap_w0
xfeed_5307 0 1 decap_w0
xfeed_5306 0 1 decap_w0
xfeed_5305 0 1 decap_w0
xfeed_5304 0 1 decap_w0
xfeed_5303 0 1 decap_w0
xfeed_5302 0 1 decap_w0
xfeed_5301 0 1 decap_w0
xfeed_5300 0 1 decap_w0
xsubckt_1243_mux2_x1 0 1 1818 2102 2069 1334 mux2_x1
xsubckt_919_mux2_x1 0 1 1897 1618 2037 1579 mux2_x1
xsubckt_783_and2_x1 0 1 1688 2046 1748 and2_x1
xsubckt_127_nand2_x0 0 1 641 1986 1994 nand2_x0
xsubckt_1302_or21nand_x0 0 1 1811 1290 1284 1282 or21nand_x0
xsubckt_1428_nand2_x0 0 1 1166 775 1976 nand2_x0
xsubckt_1625_or2_x1 0 1 969 693 1116 or2_x1
xfeed_9619 0 1 decap_w0
xfeed_9618 0 1 decap_w0
xfeed_9617 0 1 decap_w0
xfeed_9615 0 1 decap_w0
xfeed_9614 0 1 decap_w0
xfeed_9613 0 1 decap_w0
xfeed_9612 0 1 decap_w0
xfeed_9611 0 1 decap_w0
xfeed_9610 0 1 decap_w0
xfeed_5309 0 1 tie
xfeed_4699 0 1 decap_w0
xfeed_4698 0 1 decap_w0
xfeed_4696 0 1 decap_w0
xfeed_4695 0 1 decap_w0
xfeed_4694 0 1 decap_w0
xfeed_4693 0 1 decap_w0
xfeed_4692 0 1 tie
xfeed_4691 0 1 decap_w0
xfeed_4690 0 1 decap_w0
xfeed_12049 0 1 decap_w0
xfeed_12048 0 1 decap_w0
xfeed_12047 0 1 decap_w0
xfeed_12046 0 1 decap_w0
xfeed_12045 0 1 decap_w0
xfeed_12044 0 1 decap_w0
xfeed_12043 0 1 decap_w0
xfeed_12042 0 1 decap_w0
xfeed_12041 0 1 decap_w0
xfeed_12040 0 1 decap_w0
xfeed_11519 0 1 decap_w0
xfeed_11518 0 1 decap_w0
xfeed_11517 0 1 decap_w0
xfeed_11516 0 1 decap_w0
xfeed_11515 0 1 decap_w0
xfeed_11514 0 1 decap_w0
xfeed_11513 0 1 decap_w0
xfeed_11512 0 1 decap_w0
xfeed_11511 0 1 decap_w0
xfeed_11510 0 1 decap_w0
xfeed_5315 0 1 decap_w0
xfeed_5314 0 1 tie
xfeed_5313 0 1 decap_w0
xfeed_5312 0 1 decap_w0
xfeed_5311 0 1 decap_w0
xfeed_5310 0 1 decap_w0
xfeed_1009 0 1 decap_w0
xfeed_1008 0 1 decap_w0
xfeed_1007 0 1 decap_w0
xfeed_1006 0 1 decap_w0
xfeed_1005 0 1 decap_w0
xfeed_1004 0 1 decap_w0
xfeed_1003 0 1 decap_w0
xfeed_1002 0 1 decap_w0
xfeed_1001 0 1 decap_w0
xfeed_1000 0 1 decap_w0
xsubckt_1239_mux2_x1 0 1 1822 2092 2073 1334 mux2_x1
xsubckt_665_and3_x1 0 1 95 165 98 96 and3_x1
xsubckt_1656_and21nor_x0 0 1 938 948 945 942 and21nor_x0
xfeed_9629 0 1 decap_w0
xfeed_9628 0 1 decap_w0
xfeed_9627 0 1 decap_w0
xfeed_9626 0 1 decap_w0
xfeed_9625 0 1 decap_w0
xfeed_9624 0 1 decap_w0
xfeed_9623 0 1 decap_w0
xfeed_9622 0 1 decap_w0
xfeed_9621 0 1 decap_w0
xfeed_9620 0 1 decap_w0
xfeed_5319 0 1 decap_w0
xfeed_5318 0 1 decap_w0
xfeed_5317 0 1 decap_w0
xfeed_5316 0 1 decap_w0
xsubckt_995_nand2_x0 0 1 1866 1538 1534 nand2_x0
xsubckt_185_and21nor_x0 0 1 573 575 598 681 and21nor_x0
xsubckt_1321_nand2_x0 0 1 1264 1273 1266 nand2_x0
xcmpt_abc_11867_new_n1848_hfns_0 0 1 1070 1068 buf_x4
xcmpt_abc_11867_new_n1848_hfns_1 0 1 1069 1068 buf_x4
xcmpt_abc_11867_new_n1848_hfns_2 0 1 1068 1071 buf_x4
xfeed_12059 0 1 decap_w0
xfeed_12058 0 1 decap_w0
xfeed_12057 0 1 decap_w0
xfeed_12056 0 1 decap_w0
xfeed_12055 0 1 decap_w0
xfeed_12054 0 1 decap_w0
xfeed_12053 0 1 decap_w0
xfeed_12052 0 1 decap_w0
xfeed_12051 0 1 decap_w0
xfeed_12050 0 1 decap_w0
xfeed_11529 0 1 decap_w0
xfeed_11528 0 1 decap_w0
xfeed_11527 0 1 decap_w0
xfeed_11526 0 1 decap_w0
xfeed_11525 0 1 decap_w0
xfeed_11524 0 1 decap_w0
xfeed_11523 0 1 decap_w0
xfeed_11522 0 1 tie
xfeed_11520 0 1 decap_w0
xfeed_5322 0 1 decap_w0
xfeed_5321 0 1 tie
xfeed_5320 0 1 decap_w0
xfeed_1019 0 1 decap_w0
xfeed_1018 0 1 decap_w0
xfeed_1017 0 1 decap_w0
xfeed_1016 0 1 decap_w0
xfeed_1015 0 1 decap_w0
xfeed_1014 0 1 decap_w0
xfeed_1013 0 1 decap_w0
xfeed_1011 0 1 decap_w0
xfeed_1010 0 1 decap_w0
xsubckt_1147_mux2_x1 0 1 1412 770 2050 780 mux2_x1
xsubckt_1756_and21nor_x0 0 1 838 916 913 910 and21nor_x0
xfeed_9639 0 1 decap_w0
xfeed_9638 0 1 decap_w0
xfeed_9637 0 1 decap_w0
xfeed_9636 0 1 decap_w0
xfeed_9635 0 1 decap_w0
xfeed_9634 0 1 decap_w0
xfeed_9633 0 1 decap_w0
xfeed_9632 0 1 tie
xfeed_9631 0 1 decap_w0
xfeed_9630 0 1 decap_w0
xfeed_5329 0 1 decap_w0
xfeed_5328 0 1 decap_w0
xfeed_5327 0 1 decap_w0
xfeed_5326 0 1 decap_w0
xfeed_5325 0 1 decap_w0
xfeed_5324 0 1 decap_w0
xfeed_5323 0 1 decap_w0
xsubckt_1051_nand2_x0 0 1 1489 1921 1575 nand2_x0
xsubckt_457_nand2_x0 0 1 293 296 294 nand2_x0
xfeed_12069 0 1 decap_w0
xfeed_12068 0 1 decap_w0
xfeed_12067 0 1 decap_w0
xfeed_12066 0 1 decap_w0
xfeed_12065 0 1 decap_w0
xfeed_12064 0 1 decap_w0
xfeed_12063 0 1 decap_w0
xfeed_12062 0 1 decap_w0
xfeed_12061 0 1 tie
xfeed_12060 0 1 decap_w0
xfeed_11539 0 1 tie
xfeed_11538 0 1 decap_w0
xfeed_11537 0 1 decap_w0
xfeed_11536 0 1 decap_w0
xfeed_11535 0 1 decap_w0
xfeed_11534 0 1 decap_w0
xfeed_11533 0 1 decap_w0
xfeed_11532 0 1 decap_w0
xfeed_11531 0 1 decap_w0
xfeed_11530 0 1 decap_w0
xfeed_1029 0 1 decap_w0
xfeed_1028 0 1 decap_w0
xfeed_1027 0 1 decap_w0
xfeed_1026 0 1 decap_w0
xfeed_1025 0 1 decap_w0
xfeed_1024 0 1 decap_w0
xfeed_1023 0 1 decap_w0
xfeed_1022 0 1 decap_w0
xfeed_1021 0 1 decap_w0
xfeed_1020 0 1 decap_w0
xsubckt_517_and2_x1 0 1 234 539 235 and2_x1
xfeed_9649 0 1 decap_w0
xfeed_9648 0 1 decap_w0
xfeed_9647 0 1 decap_w0
xfeed_9646 0 1 tie
xfeed_9645 0 1 decap_w0
xfeed_9644 0 1 decap_w0
xfeed_9643 0 1 decap_w0
xfeed_9642 0 1 tie
xfeed_9641 0 1 decap_w0
xfeed_9640 0 1 decap_w0
xfeed_5339 0 1 decap_w0
xfeed_5338 0 1 decap_w0
xfeed_5337 0 1 decap_w0
xfeed_5336 0 1 decap_w0
xfeed_5334 0 1 decap_w0
xfeed_5333 0 1 tie
xfeed_5332 0 1 decap_w0
xfeed_5331 0 1 decap_w0
xfeed_5330 0 1 decap_w0
xfeed_4809 0 1 decap_w0
xfeed_4808 0 1 tie
xfeed_4807 0 1 decap_w0
xfeed_4805 0 1 decap_w0
xfeed_4804 0 1 decap_w0
xfeed_4803 0 1 decap_w0
xfeed_4802 0 1 decap_w0
xfeed_4801 0 1 decap_w0
xfeed_4800 0 1 decap_w0
xsubckt_729_or21nand_x0 0 1 1735 2065 1742 1740 or21nand_x0
xsubckt_706_nand3_x0 0 1 1758 211 1763 1760 nand3_x0
xsubckt_477_and3_x1 0 1 273 281 278 274 and3_x1
xfeed_12079 0 1 decap_w0
xfeed_12078 0 1 decap_w0
xfeed_12077 0 1 decap_w0
xfeed_12076 0 1 decap_w0
xfeed_12075 0 1 tie
xfeed_12074 0 1 decap_w0
xfeed_12073 0 1 decap_w0
xfeed_12072 0 1 decap_w0
xfeed_12071 0 1 decap_w0
xfeed_12070 0 1 decap_w0
xfeed_11549 0 1 decap_w0
xfeed_11548 0 1 decap_w0
xfeed_11547 0 1 decap_w0
xfeed_11546 0 1 decap_w0
xfeed_11545 0 1 decap_w0
xfeed_11544 0 1 decap_w0
xfeed_11543 0 1 decap_w0
xfeed_11542 0 1 decap_w0
xfeed_11541 0 1 decap_w0
xfeed_11540 0 1 decap_w0
xfeed_1036 0 1 tie
xfeed_1035 0 1 decap_w0
xfeed_1034 0 1 decap_w0
xfeed_1033 0 1 decap_w0
xfeed_1032 0 1 decap_w0
xfeed_1031 0 1 decap_w0
xfeed_1030 0 1 decap_w0
xsubckt_845_or4_x1 0 1 1633 1638 1637 1636 1634 or4_x1
xsubckt_834_and3_x1 0 1 1643 2068 681 490 and3_x1
xsubckt_632_or21nand_x0 0 1 126 2012 436 167 or21nand_x0
xsubckt_1301_or21nand_x0 0 1 1282 1917 1292 1285 or21nand_x0
xsubckt_1831_dff_x1 0 1 1926 25 74 dff_x1
xfeed_9659 0 1 decap_w0
xfeed_9658 0 1 decap_w0
xfeed_9657 0 1 decap_w0
xfeed_9656 0 1 decap_w0
xfeed_9655 0 1 decap_w0
xfeed_9654 0 1 decap_w0
xfeed_9653 0 1 decap_w0
xfeed_9652 0 1 decap_w0
xfeed_9651 0 1 decap_w0
xfeed_9650 0 1 decap_w0
xfeed_5349 0 1 decap_w0
xfeed_5348 0 1 decap_w0
xfeed_5347 0 1 decap_w0
xfeed_5346 0 1 decap_w0
xfeed_5345 0 1 decap_w0
xfeed_5344 0 1 decap_w0
xfeed_5343 0 1 decap_w0
xfeed_5342 0 1 decap_w0
xfeed_5340 0 1 decap_w0
xfeed_4819 0 1 decap_w0
xfeed_4818 0 1 decap_w0
xfeed_4817 0 1 tie
xfeed_4816 0 1 decap_w0
xfeed_4815 0 1 decap_w0
xfeed_4814 0 1 decap_w0
xfeed_4813 0 1 decap_w0
xfeed_4812 0 1 decap_w0
xfeed_4811 0 1 decap_w0
xfeed_4810 0 1 decap_w0
xfeed_1039 0 1 decap_w0
xfeed_1038 0 1 decap_w0
xfeed_1037 0 1 decap_w0
xsubckt_1030_nand3_x0 0 1 1504 1545 1507 1505 nand3_x0
xsubckt_350_nand2_x0 0 1 398 687 400 nand2_x0
xsubckt_359_and4_x1 0 1 389 469 431 425 390 and4_x1
xsubckt_436_nand3_x0 0 1 314 681 489 474 nand3_x0
xsubckt_499_and2_x1 0 1 252 254 253 and2_x1
xsubckt_1384_nand4_x0 0 1 1206 1245 1234 1222 1209 nand4_x0
xsubckt_1398_nand2_x0 0 1 1193 1195 1194 nand2_x0
xsubckt_1694_or21nand_x0 0 1 900 903 1122 153 or21nand_x0
xsubckt_1717_and2_x1 0 1 877 1682 878 and2_x1
xsubckt_1833_dff_x1 0 1 2045 1905 32 dff_x1
xsubckt_1835_dff_x1 0 1 2043 1903 32 dff_x1
xsubckt_1837_dff_x1 0 1 2041 1901 35 dff_x1
xfeed_12089 0 1 decap_w0
xfeed_12088 0 1 decap_w0
xfeed_12087 0 1 decap_w0
xfeed_12086 0 1 decap_w0
xfeed_12085 0 1 decap_w0
xfeed_12084 0 1 decap_w0
xfeed_12083 0 1 decap_w0
xfeed_12082 0 1 decap_w0
xfeed_12081 0 1 decap_w0
xfeed_12080 0 1 decap_w0
xfeed_11559 0 1 decap_w0
xfeed_11558 0 1 decap_w0
xfeed_11557 0 1 decap_w0
xfeed_11556 0 1 decap_w0
xfeed_11555 0 1 decap_w0
xfeed_11554 0 1 decap_w0
xfeed_11553 0 1 decap_w0
xfeed_11552 0 1 decap_w0
xfeed_11551 0 1 decap_w0
xfeed_11550 0 1 decap_w0
xfeed_1043 0 1 decap_w0
xfeed_1042 0 1 decap_w0
xfeed_1041 0 1 decap_w0
xfeed_1040 0 1 decap_w0
xsubckt_742_and3_x1 0 1 1724 1974 1749 1739 and3_x1
xsubckt_1839_dff_x1 0 1 2039 1899 32 dff_x1
xfeed_9669 0 1 decap_w0
xfeed_9668 0 1 decap_w0
xfeed_9667 0 1 tie
xfeed_9665 0 1 decap_w0
xfeed_9664 0 1 decap_w0
xfeed_9663 0 1 decap_w0
xfeed_9662 0 1 decap_w0
xfeed_9661 0 1 decap_w0
xfeed_9660 0 1 decap_w0
xfeed_5359 0 1 decap_w0
xfeed_5358 0 1 decap_w0
xfeed_5357 0 1 tie
xfeed_5356 0 1 decap_w0
xfeed_5355 0 1 decap_w0
xfeed_5354 0 1 decap_w0
xfeed_5353 0 1 decap_w0
xfeed_5352 0 1 decap_w0
xfeed_5351 0 1 decap_w0
xfeed_5350 0 1 tie
xfeed_4829 0 1 decap_w0
xfeed_4828 0 1 decap_w0
xfeed_4827 0 1 decap_w0
xfeed_4826 0 1 decap_w0
xfeed_4824 0 1 tie
xfeed_4823 0 1 decap_w0
xfeed_4821 0 1 decap_w0
xfeed_4820 0 1 decap_w0
xfeed_1049 0 1 decap_w0
xfeed_1048 0 1 decap_w0
xfeed_1047 0 1 decap_w0
xfeed_1046 0 1 decap_w0
xfeed_1045 0 1 decap_w0
xfeed_1044 0 1 decap_w0
xsubckt_1254_and21nor_x0 0 1 1326 395 595 682 and21nor_x0
xsubckt_1089_or21nand_x0 0 1 1848 771 666 784 or21nand_x0
xsubckt_1381_nand2_x0 0 1 1209 1216 1211 nand2_x0
xfeed_12099 0 1 decap_w0
xfeed_12098 0 1 decap_w0
xfeed_12097 0 1 decap_w0
xfeed_12096 0 1 decap_w0
xfeed_12095 0 1 decap_w0
xfeed_12094 0 1 decap_w0
xfeed_12093 0 1 decap_w0
xfeed_12092 0 1 decap_w0
xfeed_12091 0 1 decap_w0
xfeed_12090 0 1 decap_w0
xfeed_11569 0 1 decap_w0
xfeed_11568 0 1 decap_w0
xfeed_11567 0 1 decap_w0
xfeed_11566 0 1 decap_w0
xfeed_11565 0 1 decap_w0
xfeed_11564 0 1 decap_w0
xfeed_11563 0 1 decap_w0
xfeed_11562 0 1 decap_w0
xfeed_11561 0 1 decap_w0
xfeed_11560 0 1 decap_w0
xfeed_1050 0 1 decap_w0
xsubckt_519_nand2_x0 0 1 26 238 233 nand2_x0
xsubckt_1377_nand3_x0 0 1 1213 2071 665 657 nand3_x0
xsubckt_1435_or2_x1 0 1 1159 1165 1161 or2_x1
xfeed_9679 0 1 tie
xfeed_9678 0 1 decap_w0
xfeed_9677 0 1 decap_w0
xfeed_9676 0 1 decap_w0
xfeed_9675 0 1 decap_w0
xfeed_9674 0 1 tie
xfeed_9673 0 1 decap_w0
xfeed_9672 0 1 decap_w0
xfeed_9671 0 1 decap_w0
xfeed_9670 0 1 decap_w0
xfeed_5369 0 1 decap_w0
xfeed_5368 0 1 decap_w0
xfeed_5367 0 1 tie
xfeed_5366 0 1 decap_w0
xfeed_5365 0 1 decap_w0
xfeed_5363 0 1 decap_w0
xfeed_5362 0 1 decap_w0
xfeed_5361 0 1 decap_w0
xfeed_5360 0 1 decap_w0
xfeed_4839 0 1 decap_w0
xfeed_4838 0 1 decap_w0
xfeed_4837 0 1 decap_w0
xfeed_4836 0 1 decap_w0
xfeed_4835 0 1 decap_w0
xfeed_4834 0 1 tie
xfeed_4833 0 1 decap_w0
xfeed_4832 0 1 decap_w0
xfeed_4831 0 1 decap_w0
xfeed_4830 0 1 decap_w0
xfeed_1059 0 1 decap_w0
xfeed_1058 0 1 decap_w0
xfeed_1057 0 1 decap_w0
xfeed_1056 0 1 decap_w0
xfeed_1055 0 1 decap_w0
xfeed_1054 0 1 decap_w0
xfeed_1053 0 1 decap_w0
xfeed_1052 0 1 decap_w0
xfeed_1051 0 1 decap_w0
xsubckt_886_mux2_x1 0 1 1599 1999 2049 446 mux2_x1
xsubckt_325_nand4_x0 0 1 423 653 535 533 530 nand4_x0
xsubckt_415_nand4_x0 0 1 334 653 638 632 530 nand4_x0
xfeed_11579 0 1 decap_w0
xfeed_11578 0 1 decap_w0
xfeed_11577 0 1 decap_w0
xfeed_11576 0 1 decap_w0
xfeed_11575 0 1 decap_w0
xfeed_11574 0 1 decap_w0
xfeed_11573 0 1 decap_w0
xfeed_11572 0 1 decap_w0
xfeed_11571 0 1 decap_w0
xfeed_11570 0 1 decap_w0
xsubckt_1132_mux2_x1 0 1 1425 1426 1997 666 mux2_x1
xsubckt_1092_or21nand_x0 0 1 1455 652 428 1456 or21nand_x0
xsubckt_1006_and2_x1 0 1 1523 623 524 and2_x1
xsubckt_235_nand4_x0 0 1 516 533 530 524 518 nand4_x0
xsubckt_227_or21nand_x0 0 1 524 661 654 527 or21nand_x0
xsubckt_72_inv_x0 0 1 710 1935 inv_x0
xsubckt_70_inv_x0 0 1 712 1925 inv_x0
xsubckt_532_and4_x1 0 1 221 553 550 483 481 and4_x1
xsubckt_1441_and2_x1 0 1 1154 1975 1316 and2_x1
xsubckt_1454_and21nor_x0 0 1 1142 723 547 1745 and21nor_x0
xfeed_9689 0 1 decap_w0
xfeed_9688 0 1 decap_w0
xfeed_9687 0 1 decap_w0
xfeed_9686 0 1 decap_w0
xfeed_9685 0 1 decap_w0
xfeed_9684 0 1 decap_w0
xfeed_9683 0 1 tie
xfeed_9682 0 1 decap_w0
xfeed_9681 0 1 decap_w0
xfeed_9680 0 1 decap_w0
xfeed_5379 0 1 decap_w0
xfeed_5378 0 1 tie
xfeed_5377 0 1 decap_w0
xfeed_5376 0 1 decap_w0
xfeed_5375 0 1 decap_w0
xfeed_5374 0 1 decap_w0
xfeed_5373 0 1 decap_w0
xfeed_5372 0 1 decap_w0
xfeed_5371 0 1 decap_w0
xfeed_5370 0 1 decap_w0
xfeed_4849 0 1 decap_w0
xfeed_4848 0 1 decap_w0
xfeed_4847 0 1 decap_w0
xfeed_4846 0 1 decap_w0
xfeed_4845 0 1 decap_w0
xfeed_4844 0 1 tie
xfeed_4843 0 1 decap_w0
xfeed_4842 0 1 decap_w0
xfeed_4841 0 1 decap_w0
xfeed_4840 0 1 decap_w0
xfeed_1069 0 1 decap_w0
xfeed_1068 0 1 decap_w0
xfeed_1067 0 1 decap_w0
xfeed_1066 0 1 decap_w0
xfeed_1065 0 1 decap_w0
xfeed_1064 0 1 decap_w0
xfeed_1063 0 1 decap_w0
xfeed_1062 0 1 decap_w0
xfeed_1061 0 1 decap_w0
xfeed_1060 0 1 decap_w0
xsubckt_78_inv_x0 0 1 704 2010 inv_x0
xsubckt_76_inv_x0 0 1 706 2011 inv_x0
xsubckt_74_inv_x0 0 1 708 1931 inv_x0
xsubckt_145_and2_x1 0 1 623 661 624 and2_x1
xsubckt_1593_or21nand_x0 0 1 1001 1003 1004 1075 or21nand_x0
xsubckt_1792_nexor2_x0 0 1 802 1084 1062 nexor2_x0
xsubckt_1803_nand2_x0 0 1 792 773 2053 nand2_x0
xfeed_11589 0 1 decap_w0
xfeed_11588 0 1 tie
xfeed_11587 0 1 decap_w0
xfeed_11586 0 1 decap_w0
xfeed_11585 0 1 decap_w0
xfeed_11584 0 1 decap_w0
xfeed_11583 0 1 decap_w0
xfeed_11582 0 1 decap_w0
xfeed_11581 0 1 decap_w0
xfeed_11580 0 1 decap_w0
xsubckt_1192_or21nand_x0 0 1 1372 490 610 616 or21nand_x0
xsubckt_90_mux2_x1 0 1 694 702 701 774 mux2_x1
xsubckt_408_nand3_x0 0 1 341 687 608 595 nand3_x0
xfeed_9699 0 1 decap_w0
xfeed_9698 0 1 decap_w0
xfeed_9697 0 1 decap_w0
xfeed_9696 0 1 decap_w0
xfeed_9695 0 1 decap_w0
xfeed_9694 0 1 decap_w0
xfeed_9693 0 1 decap_w0
xfeed_9692 0 1 decap_w0
xfeed_9691 0 1 decap_w0
xfeed_9690 0 1 decap_w0
xfeed_5389 0 1 decap_w0
xfeed_5388 0 1 decap_w0
xfeed_5387 0 1 decap_w0
xfeed_5386 0 1 decap_w0
xfeed_5385 0 1 decap_w0
xfeed_5384 0 1 decap_w0
xfeed_5383 0 1 decap_w0
xfeed_5382 0 1 decap_w0
xfeed_5381 0 1 decap_w0
xfeed_5380 0 1 decap_w0
xfeed_4859 0 1 decap_w0
xfeed_4858 0 1 decap_w0
xfeed_4857 0 1 decap_w0
xfeed_4856 0 1 decap_w0
xfeed_4855 0 1 decap_w0
xfeed_4854 0 1 decap_w0
xfeed_4853 0 1 decap_w0
xfeed_4852 0 1 decap_w0
xfeed_4851 0 1 tie
xfeed_4850 0 1 decap_w0
xfeed_1079 0 1 decap_w0
xfeed_1078 0 1 decap_w0
xfeed_1077 0 1 decap_w0
xfeed_1076 0 1 decap_w0
xfeed_1075 0 1 decap_w0
xfeed_1074 0 1 decap_w0
xfeed_1073 0 1 decap_w0
xfeed_1072 0 1 decap_w0
xfeed_1071 0 1 decap_w0
xfeed_1070 0 1 decap_w0
xsubckt_1036_mux2_x1 0 1 1859 1500 1934 1576 mux2_x1
xsubckt_232_nand2_x0 0 1 519 661 521 nand2_x0
xsubckt_142_nand2_x0 0 1 626 1986 1987 nand2_x0
xsubckt_484_and21nor_x0 0 1 266 268 267 588 and21nor_x0
xsubckt_631_or21nand_x0 0 1 127 2050 601 163 or21nand_x0
xsubckt_1533_nand2_x0 0 1 1061 774 2055 nand2_x0
xsubckt_1765_nexor2_x0 0 1 829 845 841 nexor2_x0
xfeed_12209 0 1 tie
xfeed_12208 0 1 decap_w0
xfeed_12207 0 1 decap_w0
xfeed_12206 0 1 decap_w0
xfeed_12205 0 1 decap_w0
xfeed_12204 0 1 decap_w0
xfeed_12203 0 1 decap_w0
xfeed_12202 0 1 decap_w0
xfeed_12201 0 1 decap_w0
xfeed_12200 0 1 decap_w0
xfeed_11599 0 1 decap_w0
xfeed_11598 0 1 decap_w0
xfeed_11597 0 1 decap_w0
xfeed_11596 0 1 decap_w0
xfeed_11595 0 1 decap_w0
xfeed_11594 0 1 decap_w0
xfeed_11593 0 1 decap_w0
xfeed_11592 0 1 decap_w0
xfeed_11591 0 1 decap_w0
xfeed_11590 0 1 decap_w0
xfeed_6008 0 1 decap_w0
xfeed_6007 0 1 decap_w0
xfeed_6006 0 1 tie
xfeed_6005 0 1 decap_w0
xfeed_6003 0 1 decap_w0
xfeed_6002 0 1 tie
xfeed_6001 0 1 decap_w0
xfeed_6000 0 1 decap_w0
xsubckt_1205_and4_x1 0 1 1359 574 417 287 197 and4_x1
xsubckt_86_mux2_x1 0 1 696 706 705 774 mux2_x1
xsubckt_1292_or21nand_x0 0 1 1812 1300 1292 1291 or21nand_x0
xsubckt_1702_and2_x1 0 1 892 1101 893 and2_x1
xsubckt_1801_or21nand_x0 0 1 793 1917 795 794 or21nand_x0
xfeed_6009 0 1 decap_w0
xfeed_5399 0 1 decap_w0
xfeed_5398 0 1 decap_w0
xfeed_5397 0 1 decap_w0
xfeed_5396 0 1 decap_w0
xfeed_5395 0 1 decap_w0
xfeed_5394 0 1 decap_w0
xfeed_5393 0 1 decap_w0
xfeed_5392 0 1 decap_w0
xfeed_5391 0 1 decap_w0
xfeed_4869 0 1 decap_w0
xfeed_4868 0 1 decap_w0
xfeed_4867 0 1 decap_w0
xfeed_4866 0 1 decap_w0
xfeed_4865 0 1 decap_w0
xfeed_4864 0 1 decap_w0
xfeed_4863 0 1 decap_w0
xfeed_4862 0 1 decap_w0
xfeed_4861 0 1 decap_w0
xfeed_4860 0 1 decap_w0
xfeed_1089 0 1 decap_w0
xfeed_1088 0 1 decap_w0
xfeed_1087 0 1 decap_w0
xfeed_1086 0 1 decap_w0
xfeed_1085 0 1 decap_w0
xfeed_1084 0 1 decap_w0
xfeed_1083 0 1 decap_w0
xfeed_1082 0 1 decap_w0
xfeed_1081 0 1 decap_w0
xfeed_1080 0 1 decap_w0
xsubckt_1253_and2_x1 0 1 1327 1330 1328 and2_x1
xsubckt_669_nand2_x0 0 1 92 2031 175 nand2_x0
xsubckt_1489_or21nand_x0 0 1 1107 663 597 676 or21nand_x0
xfeed_12219 0 1 decap_w0
xfeed_12218 0 1 decap_w0
xfeed_12217 0 1 decap_w0
xfeed_12216 0 1 tie
xfeed_12215 0 1 decap_w0
xfeed_12214 0 1 decap_w0
xfeed_12213 0 1 decap_w0
xfeed_12212 0 1 decap_w0
xfeed_12211 0 1 decap_w0
xfeed_12210 0 1 decap_w0
xfeed_6015 0 1 decap_w0
xfeed_6014 0 1 decap_w0
xfeed_6013 0 1 decap_w0
xfeed_6012 0 1 decap_w0
xfeed_6011 0 1 decap_w0
xfeed_6010 0 1 decap_w0
xsubckt_841_and2_x1 0 1 1637 2047 1740 and2_x1
xsubckt_815_and3_x1 0 1 1660 1979 1749 1739 and3_x1
xsubckt_565_nand4_x0 0 1 190 501 462 456 403 nand4_x0
xsubckt_1754_and21nor_x0 0 1 840 880 844 842 and21nor_x0
xfeed_6019 0 1 decap_w0
xfeed_6018 0 1 decap_w0
xfeed_6017 0 1 decap_w0
xfeed_6016 0 1 tie
xfeed_4879 0 1 tie
xfeed_4878 0 1 decap_w0
xfeed_4877 0 1 decap_w0
xfeed_4876 0 1 decap_w0
xfeed_4875 0 1 decap_w0
xfeed_4874 0 1 decap_w0
xfeed_4873 0 1 decap_w0
xfeed_4872 0 1 decap_w0
xfeed_4871 0 1 decap_w0
xfeed_4870 0 1 decap_w0
xfeed_1099 0 1 decap_w0
xfeed_1098 0 1 decap_w0
xfeed_1097 0 1 decap_w0
xfeed_1096 0 1 decap_w0
xfeed_1095 0 1 decap_w0
xfeed_1094 0 1 decap_w0
xfeed_1093 0 1 decap_w0
xfeed_1092 0 1 tie
xfeed_1091 0 1 decap_w0
xfeed_1090 0 1 decap_w0
xsubckt_1249_and2_x1 0 1 1331 666 661 and2_x1
xsubckt_1169_nand3_x0 0 1 1393 1934 609 603 nand3_x0
xsubckt_723_and3_x1 0 1 1741 592 574 478 and3_x1
xsubckt_207_nand4_x0 0 1 547 716 1924 682 670 nand4_x0
xsubckt_475_nand4_x0 0 1 275 680 674 670 558 nand4_x0
xsubckt_1805_or3_x1 0 1 790 773 846 791 or3_x1
xfeed_12229 0 1 decap_w0
xfeed_12228 0 1 decap_w0
xfeed_12227 0 1 decap_w0
xfeed_12226 0 1 decap_w0
xfeed_12225 0 1 decap_w0
xfeed_12224 0 1 decap_w0
xfeed_12223 0 1 decap_w0
xfeed_12222 0 1 decap_w0
xfeed_12221 0 1 decap_w0
xfeed_12220 0 1 decap_w0
xfeed_6022 0 1 decap_w0
xfeed_6021 0 1 decap_w0
xfeed_6020 0 1 decap_w0
xsubckt_388_and2_x1 0 1 361 370 362 and2_x1
xsubckt_1492_or21nand_x0 0 1 1104 1106 1143 739 or21nand_x0
xsubckt_1600_or21nand_x0 0 1 994 1649 1116 692 or21nand_x0
xsubckt_1732_mux2_x1 0 1 862 868 864 875 mux2_x1
xfeed_9809 0 1 decap_w0
xfeed_9808 0 1 decap_w0
xfeed_9807 0 1 decap_w0
xfeed_9806 0 1 decap_w0
xfeed_9805 0 1 decap_w0
xfeed_9804 0 1 decap_w0
xfeed_9803 0 1 decap_w0
xfeed_9802 0 1 decap_w0
xfeed_9801 0 1 decap_w0
xfeed_9800 0 1 tie
xfeed_6029 0 1 decap_w0
xfeed_6028 0 1 decap_w0
xfeed_6027 0 1 decap_w0
xfeed_6026 0 1 decap_w0
xfeed_6025 0 1 decap_w0
xfeed_6024 0 1 decap_w0
xfeed_6023 0 1 decap_w0
xfeed_4889 0 1 decap_w0
xfeed_4888 0 1 decap_w0
xfeed_4887 0 1 decap_w0
xfeed_4886 0 1 decap_w0
xfeed_4885 0 1 decap_w0
xfeed_4884 0 1 tie
xfeed_4883 0 1 decap_w0
xfeed_4882 0 1 decap_w0
xfeed_4881 0 1 decap_w0
xfeed_4880 0 1 decap_w0
xsubckt_871_mux2_x1 0 1 1912 2020 1612 1619 mux2_x1
xsubckt_1288_or21nand_x0 0 1 1294 1295 1322 765 or21nand_x0
xsubckt_1592_or21nand_x0 0 1 1002 1067 1014 1072 or21nand_x0
xsubckt_1728_mux2_x1 0 1 866 1103 1105 870 mux2_x1
xfeed_12239 0 1 decap_w0
xfeed_12238 0 1 decap_w0
xfeed_12237 0 1 decap_w0
xfeed_12236 0 1 decap_w0
xfeed_12235 0 1 decap_w0
xfeed_12234 0 1 decap_w0
xfeed_12233 0 1 tie
xfeed_12232 0 1 decap_w0
xfeed_12231 0 1 decap_w0
xfeed_12230 0 1 decap_w0
xfeed_11709 0 1 decap_w0
xfeed_11708 0 1 decap_w0
xfeed_11707 0 1 decap_w0
xfeed_11706 0 1 decap_w0
xfeed_11705 0 1 tie
xfeed_11704 0 1 decap_w0
xfeed_11703 0 1 decap_w0
xfeed_11702 0 1 decap_w0
xfeed_11701 0 1 decap_w0
xfeed_11700 0 1 tie
xsubckt_811_nand3_x0 0 1 1663 2071 680 490 nand3_x0
xsubckt_296_and2_x1 0 1 452 1927 713 and2_x1
xsubckt_204_nand2_x0 0 1 550 687 552 nand2_x0
xsubckt_1553_and21nor_x0 0 1 1041 1102 1044 1043 and21nor_x0
xsubckt_1789_or21nand_x0 0 1 805 1083 1066 1064 or21nand_x0
xfeed_9819 0 1 decap_w0
xfeed_9818 0 1 decap_w0
xfeed_9817 0 1 decap_w0
xfeed_9816 0 1 decap_w0
xfeed_9815 0 1 decap_w0
xfeed_9814 0 1 decap_w0
xfeed_9813 0 1 decap_w0
xfeed_9812 0 1 decap_w0
xfeed_9810 0 1 tie
xfeed_6039 0 1 decap_w0
xfeed_6038 0 1 decap_w0
xfeed_6037 0 1 decap_w0
xfeed_6036 0 1 decap_w0
xfeed_6035 0 1 decap_w0
xfeed_6034 0 1 decap_w0
xfeed_6033 0 1 decap_w0
xfeed_6032 0 1 decap_w0
xfeed_6031 0 1 decap_w0
xfeed_6030 0 1 decap_w0
xfeed_5509 0 1 decap_w0
xfeed_5508 0 1 decap_w0
xfeed_5507 0 1 decap_w0
xfeed_5506 0 1 decap_w0
xfeed_5505 0 1 decap_w0
xfeed_5504 0 1 decap_w0
xfeed_5503 0 1 decap_w0
xfeed_5502 0 1 decap_w0
xfeed_5501 0 1 decap_w0
xfeed_5500 0 1 tie
xfeed_4899 0 1 decap_w0
xfeed_4898 0 1 decap_w0
xfeed_4897 0 1 decap_w0
xfeed_4896 0 1 decap_w0
xfeed_4895 0 1 decap_w0
xfeed_4894 0 1 decap_w0
xfeed_4893 0 1 tie
xfeed_4891 0 1 decap_w0
xfeed_4890 0 1 decap_w0
xsubckt_1152_and21nor_x0 0 1 1408 666 610 603 and21nor_x0
xsubckt_1113_mux2_x1 0 1 1844 2002 1993 1438 mux2_x1
xsubckt_985_nand4_x0 0 1 1542 638 632 622 1544 nand4_x0
xsubckt_130_and2_x1 0 1 638 660 639 and2_x1
xsubckt_1415_nand2_x0 0 1 1178 1977 1316 nand2_x0
xsubckt_1692_or21nand_x0 0 1 902 905 1118 768 or21nand_x0
xfeed_12249 0 1 decap_w0
xfeed_12247 0 1 decap_w0
xfeed_12246 0 1 decap_w0
xfeed_12245 0 1 decap_w0
xfeed_12244 0 1 decap_w0
xfeed_12243 0 1 decap_w0
xfeed_12242 0 1 decap_w0
xfeed_12241 0 1 decap_w0
xfeed_12240 0 1 decap_w0
xfeed_11719 0 1 decap_w0
xfeed_11718 0 1 decap_w0
xfeed_11717 0 1 decap_w0
xfeed_11716 0 1 decap_w0
xfeed_11715 0 1 decap_w0
xfeed_11714 0 1 decap_w0
xfeed_11713 0 1 decap_w0
xfeed_11712 0 1 decap_w0
xfeed_11711 0 1 decap_w0
xfeed_11710 0 1 decap_w0
xsubckt_541_nand3_x0 0 1 24 215 214 213 nand3_x0
xsubckt_1291_or21nand_x0 0 1 1291 1917 1302 1293 or21nand_x0
xdiode_109 0 1 2052 diode_w1
xdiode_108 0 1 2052 diode_w1
xdiode_107 0 1 2052 diode_w1
xdiode_106 0 1 2051 diode_w1
xdiode_105 0 1 2051 diode_w1
xdiode_104 0 1 2051 diode_w1
xdiode_103 0 1 2050 diode_w1
xdiode_102 0 1 2050 diode_w1
xdiode_101 0 1 2050 diode_w1
xdiode_100 0 1 2049 diode_w1
xfeed_9829 0 1 decap_w0
xfeed_9828 0 1 decap_w0
xfeed_9827 0 1 decap_w0
xfeed_9826 0 1 decap_w0
xfeed_9825 0 1 decap_w0
xfeed_9824 0 1 decap_w0
xfeed_9823 0 1 decap_w0
xfeed_9822 0 1 decap_w0
xfeed_9821 0 1 decap_w0
xfeed_9820 0 1 decap_w0
xfeed_6049 0 1 decap_w0
xfeed_6048 0 1 decap_w0
xfeed_6047 0 1 decap_w0
xfeed_6046 0 1 decap_w0
xfeed_6045 0 1 decap_w0
xfeed_6044 0 1 decap_w0
xfeed_6043 0 1 decap_w0
xfeed_6042 0 1 decap_w0
xfeed_6041 0 1 decap_w0
xfeed_6040 0 1 decap_w0
xfeed_5519 0 1 decap_w0
xfeed_5518 0 1 decap_w0
xfeed_5517 0 1 decap_w0
xfeed_5515 0 1 decap_w0
xfeed_5514 0 1 decap_w0
xfeed_5513 0 1 decap_w0
xfeed_5512 0 1 tie
xfeed_5511 0 1 decap_w0
xfeed_5510 0 1 decap_w0
xfeed_1209 0 1 decap_w0
xfeed_1208 0 1 decap_w0
xfeed_1207 0 1 decap_w0
xfeed_1206 0 1 decap_w0
xfeed_1205 0 1 decap_w0
xfeed_1204 0 1 decap_w0
xfeed_1203 0 1 decap_w0
xfeed_1202 0 1 tie
xfeed_1201 0 1 decap_w0
xfeed_1200 0 1 decap_w0
xsubckt_1109_mux2_x1 0 1 1439 1443 1986 1441 mux2_x1
xfeed_12259 0 1 decap_w0
xfeed_12258 0 1 decap_w0
xfeed_12257 0 1 decap_w0
xfeed_12256 0 1 tie
xfeed_12255 0 1 decap_w0
xfeed_12254 0 1 decap_w0
xfeed_12253 0 1 decap_w0
xfeed_12252 0 1 decap_w0
xfeed_12251 0 1 decap_w0
xfeed_12250 0 1 decap_w0
xfeed_11729 0 1 decap_w0
xfeed_11728 0 1 decap_w0
xfeed_11727 0 1 decap_w0
xfeed_11726 0 1 decap_w0
xfeed_11725 0 1 decap_w0
xfeed_11724 0 1 decap_w0
xfeed_11723 0 1 decap_w0
xfeed_11722 0 1 decap_w0
xfeed_11721 0 1 decap_w0
xfeed_11720 0 1 decap_w0
xsubckt_978_nand3_x0 0 1 1549 637 633 383 nand3_x0
xdiode_119 0 1 2047 diode_w1
xdiode_118 0 1 2046 diode_w1
xdiode_117 0 1 2046 diode_w1
xdiode_116 0 1 2046 diode_w1
xdiode_115 0 1 2046 diode_w1
xdiode_114 0 1 2046 diode_w1
xdiode_113 0 1 2053 diode_w1
xdiode_112 0 1 2053 diode_w1
xdiode_111 0 1 2053 diode_w1
xdiode_110 0 1 2053 diode_w1
xfeed_9838 0 1 decap_w0
xfeed_9837 0 1 decap_w0
xfeed_9835 0 1 tie
xfeed_9834 0 1 decap_w0
xfeed_9833 0 1 decap_w0
xfeed_9831 0 1 decap_w0
xfeed_9830 0 1 decap_w0
xfeed_6059 0 1 decap_w0
xfeed_6058 0 1 decap_w0
xfeed_6057 0 1 decap_w0
xfeed_6056 0 1 decap_w0
xfeed_6055 0 1 decap_w0
xfeed_6054 0 1 decap_w0
xfeed_6053 0 1 decap_w0
xfeed_6052 0 1 decap_w0
xfeed_6051 0 1 decap_w0
xfeed_6050 0 1 decap_w0
xfeed_5529 0 1 decap_w0
xfeed_5528 0 1 decap_w0
xfeed_5527 0 1 decap_w0
xfeed_5526 0 1 decap_w0
xfeed_5525 0 1 decap_w0
xfeed_5524 0 1 decap_w0
xfeed_5523 0 1 decap_w0
xfeed_5522 0 1 decap_w0
xfeed_5521 0 1 tie
xfeed_5520 0 1 decap_w0
xfeed_1219 0 1 decap_w0
xfeed_1218 0 1 decap_w0
xfeed_1217 0 1 decap_w0
xfeed_1216 0 1 decap_w0
xfeed_1215 0 1 decap_w0
xfeed_1214 0 1 decap_w0
xfeed_1213 0 1 decap_w0
xfeed_1212 0 1 decap_w0
xfeed_1211 0 1 tie
xfeed_1210 0 1 decap_w0
xsubckt_379_and21nor_x0 0 1 370 372 371 535 and21nor_x0
xsubckt_443_and3_x1 0 1 307 379 375 308 and3_x1
xsubckt_1290_and3_x1 0 1 1292 1311 1303 1293 and3_x1
xfeed_12269 0 1 decap_w0
xfeed_12268 0 1 tie
xfeed_12267 0 1 decap_w0
xfeed_12266 0 1 decap_w0
xfeed_12265 0 1 decap_w0
xfeed_12264 0 1 decap_w0
xfeed_12263 0 1 decap_w0
xfeed_12262 0 1 decap_w0
xfeed_12261 0 1 decap_w0
xfeed_12260 0 1 decap_w0
xfeed_11739 0 1 decap_w0
xfeed_11738 0 1 decap_w0
xfeed_11737 0 1 decap_w0
xfeed_11736 0 1 decap_w0
xfeed_11735 0 1 decap_w0
xfeed_11734 0 1 decap_w0
xfeed_11733 0 1 decap_w0
xfeed_11732 0 1 decap_w0
xfeed_11731 0 1 decap_w0
xfeed_11730 0 1 decap_w0
xsubckt_465_and2_x1 0 1 285 287 286 and2_x1
xsubckt_1549_and21nor_x0 0 1 1045 1104 1050 1048 and21nor_x0
xsubckt_1745_nand2_x0 0 1 849 852 851 nand2_x0
xdiode_129 0 1 581 diode_w1
xdiode_128 0 1 581 diode_w1
xdiode_127 0 1 524 diode_w1
xdiode_126 0 1 524 diode_w1
xdiode_125 0 1 524 diode_w1
xdiode_124 0 1 623 diode_w1
xdiode_123 0 1 623 diode_w1
xdiode_122 0 1 623 diode_w1
xdiode_121 0 1 2047 diode_w1
xdiode_120 0 1 2047 diode_w1
xfeed_9849 0 1 decap_w0
xfeed_9848 0 1 decap_w0
xfeed_9847 0 1 decap_w0
xfeed_9846 0 1 decap_w0
xfeed_9845 0 1 tie
xfeed_9844 0 1 decap_w0
xfeed_9843 0 1 decap_w0
xfeed_9842 0 1 decap_w0
xfeed_9841 0 1 decap_w0
xfeed_9840 0 1 tie
xfeed_6069 0 1 decap_w0
xfeed_6068 0 1 decap_w0
xfeed_6067 0 1 decap_w0
xfeed_6066 0 1 decap_w0
xfeed_6064 0 1 decap_w0
xfeed_6063 0 1 decap_w0
xfeed_6062 0 1 decap_w0
xfeed_6061 0 1 tie
xfeed_6060 0 1 decap_w0
xfeed_5539 0 1 decap_w0
xfeed_5538 0 1 decap_w0
xfeed_5537 0 1 decap_w0
xfeed_5536 0 1 decap_w0
xfeed_5535 0 1 decap_w0
xfeed_5534 0 1 decap_w0
xfeed_5533 0 1 tie
xfeed_5532 0 1 decap_w0
xfeed_5531 0 1 decap_w0
xfeed_5530 0 1 decap_w0
xfeed_1229 0 1 decap_w0
xfeed_1227 0 1 decap_w0
xfeed_1226 0 1 decap_w0
xfeed_1225 0 1 decap_w0
xfeed_1224 0 1 decap_w0
xfeed_1223 0 1 decap_w0
xfeed_1222 0 1 decap_w0
xfeed_1221 0 1 decap_w0
xfeed_1220 0 1 decap_w0
xsubckt_1208_and3_x1 0 1 1356 1379 1359 1357 and3_x1
xsubckt_479_and21nor_x0 0 1 271 272 289 687 and21nor_x0
xsubckt_1840_dff_x1 0 1 2038 1898 32 dff_x1
xsubckt_1842_dff_x1 0 1 2036 1896 35 dff_x1
xsubckt_1844_dff_x1 0 1 2034 1894 32 dff_x1
xfeed_12279 0 1 decap_w0
xfeed_12278 0 1 decap_w0
xfeed_12277 0 1 decap_w0
xfeed_12276 0 1 decap_w0
xfeed_12275 0 1 decap_w0
xfeed_12274 0 1 decap_w0
xfeed_12273 0 1 decap_w0
xfeed_12272 0 1 decap_w0
xfeed_12271 0 1 decap_w0
xfeed_12270 0 1 decap_w0
xfeed_11749 0 1 tie
xfeed_11748 0 1 decap_w0
xfeed_11747 0 1 decap_w0
xfeed_11746 0 1 decap_w0
xfeed_11745 0 1 decap_w0
xfeed_11744 0 1 decap_w0
xfeed_11743 0 1 decap_w0
xfeed_11742 0 1 decap_w0
xfeed_11741 0 1 decap_w0
xfeed_11740 0 1 decap_w0
xsubckt_782_and3_x1 0 1 1689 1969 1749 1739 and3_x1
xsubckt_264_nand2_x0 0 1 484 609 495 nand2_x0
xsubckt_250_nand4_x0 0 1 501 1929 715 679 670 nand4_x0
xsubckt_233_and4_x1 0 1 518 661 626 625 521 and4_x1
xsubckt_1788_or21nand_x0 0 1 806 1028 812 810 or21nand_x0
xsubckt_1846_dff_x1 0 1 2032 1892 32 dff_x1
xsubckt_1848_dff_x1 0 1 2030 1890 32 dff_x1
xdiode_139 0 1 2055 diode_w1
xdiode_138 0 1 2055 diode_w1
xdiode_137 0 1 1961 diode_w1
xdiode_136 0 1 1961 diode_w1
xdiode_135 0 1 1961 diode_w1
xdiode_134 0 1 1961 diode_w1
xdiode_133 0 1 67 diode_w1
xdiode_132 0 1 67 diode_w1
xdiode_131 0 1 581 diode_w1
xdiode_130 0 1 581 diode_w1
xfeed_9859 0 1 decap_w0
xfeed_9857 0 1 decap_w0
xfeed_9856 0 1 decap_w0
xfeed_9855 0 1 decap_w0
xfeed_9854 0 1 decap_w0
xfeed_9853 0 1 decap_w0
xfeed_9852 0 1 decap_w0
xfeed_9851 0 1 decap_w0
xfeed_9850 0 1 decap_w0
xfeed_6079 0 1 decap_w0
xfeed_6078 0 1 decap_w0
xfeed_6077 0 1 decap_w0
xfeed_6076 0 1 decap_w0
xfeed_6075 0 1 tie
xfeed_6074 0 1 decap_w0
xfeed_6073 0 1 decap_w0
xfeed_6072 0 1 decap_w0
xfeed_6071 0 1 decap_w0
xfeed_6070 0 1 decap_w0
xfeed_5549 0 1 decap_w0
xfeed_5548 0 1 decap_w0
xfeed_5547 0 1 decap_w0
xfeed_5546 0 1 decap_w0
xfeed_5545 0 1 decap_w0
xfeed_5544 0 1 decap_w0
xfeed_5543 0 1 decap_w0
xfeed_5542 0 1 decap_w0
xfeed_5541 0 1 decap_w0
xfeed_5540 0 1 tie
xfeed_1239 0 1 decap_w0
xfeed_1238 0 1 decap_w0
xfeed_1237 0 1 decap_w0
xfeed_1236 0 1 decap_w0
xfeed_1235 0 1 decap_w0
xfeed_1234 0 1 decap_w0
xfeed_1233 0 1 decap_w0
xfeed_1232 0 1 decap_w0
xfeed_1231 0 1 decap_w0
xfeed_1230 0 1 decap_w0
xsubckt_513_nand3_x0 0 1 238 315 271 239 nand3_x0
xsubckt_1385_nand2_x0 0 1 1205 1916 1206 nand2_x0
xfeed_12289 0 1 decap_w0
xfeed_12288 0 1 decap_w0
xfeed_12287 0 1 decap_w0
xfeed_12286 0 1 decap_w0
xfeed_12285 0 1 decap_w0
xfeed_12284 0 1 decap_w0
xfeed_12283 0 1 decap_w0
xfeed_12282 0 1 decap_w0
xfeed_12281 0 1 decap_w0
xfeed_12280 0 1 decap_w0
xfeed_11759 0 1 decap_w0
xfeed_11758 0 1 decap_w0
xfeed_11757 0 1 decap_w0
xfeed_11756 0 1 decap_w0
xfeed_11755 0 1 decap_w0
xfeed_11754 0 1 decap_w0
xfeed_11753 0 1 decap_w0
xfeed_11752 0 1 decap_w0
xfeed_11751 0 1 decap_w0
xfeed_11750 0 1 decap_w0
xsubckt_1138_and2_x1 0 1 1420 1423 1421 and2_x1
xsubckt_423_nand3_x0 0 1 326 687 610 598 nand3_x0
xsubckt_1749_and21nor_x0 0 1 845 854 850 847 and21nor_x0
xdiode_149 0 1 558 diode_w1
xdiode_148 0 1 558 diode_w1
xdiode_147 0 1 558 diode_w1
xdiode_146 0 1 557 diode_w1
xdiode_145 0 1 557 diode_w1
xdiode_144 0 1 557 diode_w1
xdiode_143 0 1 557 diode_w1
xdiode_142 0 1 557 diode_w1
xdiode_141 0 1 2055 diode_w1
xdiode_140 0 1 2055 diode_w1
xfeed_9869 0 1 decap_w0
xfeed_9868 0 1 decap_w0
xfeed_9867 0 1 decap_w0
xfeed_9866 0 1 decap_w0
xfeed_9865 0 1 decap_w0
xfeed_9864 0 1 decap_w0
xfeed_9863 0 1 decap_w0
xfeed_9862 0 1 decap_w0
xfeed_9861 0 1 decap_w0
xfeed_9860 0 1 decap_w0
xfeed_6089 0 1 decap_w0
xfeed_6088 0 1 decap_w0
xfeed_6087 0 1 decap_w0
xfeed_6086 0 1 decap_w0
xfeed_6085 0 1 decap_w0
xfeed_6084 0 1 decap_w0
xfeed_6083 0 1 decap_w0
xfeed_6082 0 1 tie
xfeed_6081 0 1 decap_w0
xfeed_6080 0 1 decap_w0
xfeed_5559 0 1 decap_w0
xfeed_5558 0 1 decap_w0
xfeed_5557 0 1 decap_w0
xfeed_5556 0 1 tie
xfeed_5555 0 1 decap_w0
xfeed_5553 0 1 decap_w0
xfeed_5552 0 1 decap_w0
xfeed_5551 0 1 decap_w0
xfeed_5550 0 1 decap_w0
xfeed_1249 0 1 decap_w0
xfeed_1248 0 1 decap_w0
xfeed_1247 0 1 decap_w0
xfeed_1246 0 1 decap_w0
xfeed_1245 0 1 decap_w0
xfeed_1244 0 1 decap_w0
xfeed_1243 0 1 decap_w0
xfeed_1242 0 1 decap_w0
xfeed_1241 0 1 decap_w0
xfeed_1240 0 1 decap_w0
xsubckt_1191_nand4_x0 0 1 1373 1929 715 711 670 nand4_x0
xsubckt_333_nand3_x0 0 1 415 609 557 421 nand3_x0
xsubckt_1544_nand3_x0 0 1 1050 1970 679 595 nand3_x0
xfeed_12299 0 1 decap_w0
xfeed_12298 0 1 decap_w0
xfeed_12297 0 1 decap_w0
xfeed_12296 0 1 tie
xfeed_12295 0 1 decap_w0
xfeed_12294 0 1 decap_w0
xfeed_12293 0 1 decap_w0
xfeed_12292 0 1 decap_w0
xfeed_12291 0 1 tie
xfeed_12290 0 1 decap_w0
xfeed_11769 0 1 decap_w0
xfeed_11768 0 1 decap_w0
xfeed_11767 0 1 decap_w0
xfeed_11766 0 1 decap_w0
xfeed_11765 0 1 decap_w0
xfeed_11764 0 1 decap_w0
xfeed_11763 0 1 decap_w0
xfeed_11762 0 1 decap_w0
xfeed_11761 0 1 decap_w0
xfeed_11760 0 1 decap_w0
xsubckt_905_nexor2_x0 0 1 1583 759 1584 nexor2_x0
xsubckt_163_and3_x1 0 1 598 716 1924 599 and3_x1
xsubckt_137_and4_x1 0 1 631 660 639 636 635 and4_x1
xsubckt_572_and4_x1 0 1 183 1951 681 674 670 and4_x1
xsubckt_1569_and2_x1 0 1 1025 1642 1026 and2_x1
xsubckt_1617_mux2_x1 0 1 977 1020 979 1142 mux2_x1
xdiode_159 0 1 548 diode_w1
xdiode_158 0 1 1917 diode_w1
xdiode_157 0 1 1917 diode_w1
xdiode_156 0 1 1917 diode_w1
xdiode_155 0 1 1917 diode_w1
xdiode_154 0 1 1917 diode_w1
xdiode_153 0 1 1917 diode_w1
xdiode_152 0 1 1917 diode_w1
xdiode_151 0 1 1917 diode_w1
xdiode_150 0 1 1917 diode_w1
xfeed_9879 0 1 decap_w0
xfeed_9878 0 1 decap_w0
xfeed_9877 0 1 decap_w0
xfeed_9876 0 1 decap_w0
xfeed_9875 0 1 tie
xfeed_9874 0 1 decap_w0
xfeed_9873 0 1 decap_w0
xfeed_9872 0 1 decap_w0
xfeed_9871 0 1 decap_w0
xfeed_9870 0 1 decap_w0
xfeed_6099 0 1 decap_w0
xfeed_6098 0 1 decap_w0
xfeed_6097 0 1 decap_w0
xfeed_6096 0 1 tie
xfeed_6095 0 1 decap_w0
xfeed_6094 0 1 decap_w0
xfeed_6093 0 1 decap_w0
xfeed_6092 0 1 tie
xfeed_6091 0 1 decap_w0
xfeed_6090 0 1 decap_w0
xfeed_5569 0 1 decap_w0
xfeed_5568 0 1 decap_w0
xfeed_5567 0 1 tie
xfeed_5566 0 1 decap_w0
xfeed_5565 0 1 decap_w0
xfeed_5564 0 1 decap_w0
xfeed_5563 0 1 tie
xfeed_5562 0 1 decap_w0
xfeed_5561 0 1 decap_w0
xfeed_5560 0 1 decap_w0
xfeed_1259 0 1 decap_w0
xfeed_1257 0 1 decap_w0
xfeed_1256 0 1 decap_w0
xfeed_1255 0 1 decap_w0
xfeed_1254 0 1 decap_w0
xfeed_1253 0 1 decap_w0
xfeed_1252 0 1 decap_w0
xfeed_1251 0 1 decap_w0
xfeed_1250 0 1 decap_w0
xsubckt_1100_nand2_x0 0 1 1447 1476 1448 nand2_x0
xsubckt_684_nand2_x0 0 1 1779 2038 172 nand2_x0
xsubckt_81_inv_x0 0 1 701 2088 inv_x0
xsubckt_83_inv_x0 0 1 699 2087 inv_x0
xsubckt_85_inv_x0 0 1 697 2086 inv_x0
xfeed_11779 0 1 decap_w0
xfeed_11778 0 1 tie
xfeed_11777 0 1 decap_w0
xfeed_11776 0 1 decap_w0
xfeed_11775 0 1 decap_w0
xfeed_11774 0 1 decap_w0
xfeed_11773 0 1 decap_w0
xfeed_11772 0 1 decap_w0
xfeed_11771 0 1 decap_w0
xfeed_11770 0 1 decap_w0
xsubckt_1274_nand3_x0 0 1 1307 2064 665 657 nand3_x0
xsubckt_87_inv_x0 0 1 2003 696 inv_x0
xsubckt_89_inv_x0 0 1 2002 695 inv_x0
xsubckt_107_and2_x1 0 1 671 1927 1928 and2_x1
xdiode_169 0 1 603 diode_w1
xdiode_168 0 1 603 diode_w1
xdiode_167 0 1 714 diode_w1
xdiode_166 0 1 714 diode_w1
xdiode_165 0 1 460 diode_w1
xdiode_164 0 1 460 diode_w1
xdiode_163 0 1 460 diode_w1
xdiode_162 0 1 548 diode_w1
xdiode_161 0 1 548 diode_w1
xdiode_160 0 1 548 diode_w1
xfeed_9889 0 1 decap_w0
xfeed_9888 0 1 decap_w0
xfeed_9887 0 1 decap_w0
xfeed_9886 0 1 decap_w0
xfeed_9885 0 1 decap_w0
xfeed_9884 0 1 decap_w0
xfeed_9883 0 1 decap_w0
xfeed_9882 0 1 tie
xfeed_9881 0 1 decap_w0
xfeed_9880 0 1 decap_w0
xfeed_5579 0 1 decap_w0
xfeed_5578 0 1 decap_w0
xfeed_5577 0 1 decap_w0
xfeed_5576 0 1 decap_w0
xfeed_5575 0 1 tie
xfeed_5574 0 1 decap_w0
xfeed_5573 0 1 decap_w0
xfeed_5572 0 1 decap_w0
xfeed_5571 0 1 tie
xfeed_5570 0 1 decap_w0
xfeed_1269 0 1 decap_w0
xfeed_1268 0 1 decap_w0
xfeed_1267 0 1 decap_w0
xfeed_1266 0 1 decap_w0
xfeed_1265 0 1 decap_w0
xfeed_1264 0 1 decap_w0
xfeed_1263 0 1 decap_w0
xfeed_1262 0 1 decap_w0
xfeed_1261 0 1 decap_w0
xfeed_1260 0 1 decap_w0
xsubckt_843_nand3_x0 0 1 1635 2067 682 490 nand3_x0
xsubckt_1720_and3_x1 0 1 874 1982 678 595 and3_x1
xfeed_11789 0 1 decap_w0
xfeed_11788 0 1 decap_w0
xfeed_11787 0 1 decap_w0
xfeed_11786 0 1 decap_w0
xfeed_11785 0 1 decap_w0
xfeed_11784 0 1 decap_w0
xfeed_11783 0 1 decap_w0
xfeed_11782 0 1 decap_w0
xfeed_11781 0 1 decap_w0
xfeed_11780 0 1 decap_w0
xsubckt_146_nand2_x0 0 1 622 661 624 nand2_x0
xsubckt_450_and2_x1 0 1 300 652 360 and2_x1
xsubckt_538_and2_x1 0 1 215 252 216 and2_x1
xsubckt_1343_nand4_x0 0 1 1244 1273 1266 1257 1247 nand4_x0
xsubckt_1357_nand2_x0 0 1 1231 1233 1232 nand2_x0
xsubckt_1648_and21nor_x0 0 1 946 1070 958 1073 and21nor_x0
xsubckt_1700_nand2_x0 0 1 894 1105 896 nand2_x0
xdiode_179 0 1 490 diode_w1
xdiode_178 0 1 490 diode_w1
xdiode_177 0 1 490 diode_w1
xdiode_176 0 1 490 diode_w1
xdiode_175 0 1 490 diode_w1
xdiode_174 0 1 489 diode_w1
xdiode_173 0 1 489 diode_w1
xdiode_172 0 1 489 diode_w1
xdiode_171 0 1 489 diode_w1
xdiode_170 0 1 603 diode_w1
xfeed_9899 0 1 decap_w0
xfeed_9898 0 1 decap_w0
xfeed_9897 0 1 decap_w0
xfeed_9896 0 1 decap_w0
xfeed_9895 0 1 decap_w0
xfeed_9894 0 1 decap_w0
xfeed_9893 0 1 decap_w0
xfeed_9892 0 1 tie
xfeed_9891 0 1 decap_w0
xfeed_9890 0 1 decap_w0
xfeed_5589 0 1 decap_w0
xfeed_5588 0 1 decap_w0
xfeed_5587 0 1 decap_w0
xfeed_5586 0 1 decap_w0
xfeed_5585 0 1 decap_w0
xfeed_5584 0 1 tie
xfeed_5583 0 1 decap_w0
xfeed_5582 0 1 decap_w0
xfeed_5581 0 1 decap_w0
xfeed_5580 0 1 tie
xfeed_1279 0 1 decap_w0
xfeed_1278 0 1 decap_w0
xfeed_1277 0 1 decap_w0
xfeed_1276 0 1 decap_w0
xfeed_1275 0 1 decap_w0
xfeed_1274 0 1 decap_w0
xfeed_1273 0 1 decap_w0
xfeed_1272 0 1 decap_w0
xfeed_1271 0 1 decap_w0
xfeed_1270 0 1 decap_w0
xsubckt_622_nor2_x0 0 1 135 137 136 nor2_x0
xsubckt_1386_or21nand_x0 0 1 1804 1217 1208 1205 or21nand_x0
xfeed_12409 0 1 decap_w0
xfeed_12408 0 1 decap_w0
xfeed_12407 0 1 decap_w0
xfeed_12406 0 1 decap_w0
xfeed_12405 0 1 decap_w0
xfeed_12404 0 1 decap_w0
xfeed_12403 0 1 decap_w0
xfeed_12402 0 1 decap_w0
xfeed_12401 0 1 decap_w0
xfeed_12400 0 1 decap_w0
xfeed_11799 0 1 decap_w0
xfeed_11798 0 1 decap_w0
xfeed_11797 0 1 decap_w0
xfeed_11796 0 1 decap_w0
xfeed_11795 0 1 decap_w0
xfeed_11794 0 1 decap_w0
xfeed_11793 0 1 decap_w0
xfeed_11792 0 1 decap_w0
xfeed_11791 0 1 decap_w0
xfeed_11790 0 1 decap_w0
xsubckt_1215_and2_x1 0 1 1349 547 467 and2_x1
xsubckt_446_and2_x1 0 1 304 307 305 and2_x1
xsubckt_569_nand4_x0 0 1 186 1950 681 674 670 nand4_x0
xsubckt_1430_nand2_x0 0 1 1164 2047 479 nand2_x0
xsubckt_1690_or21nand_x0 0 1 904 1670 1116 695 or21nand_x0
xdiode_189 0 1 773 diode_w1
xdiode_188 0 1 617 diode_w1
xdiode_187 0 1 617 diode_w1
xdiode_186 0 1 616 diode_w1
xdiode_185 0 1 616 diode_w1
xdiode_184 0 1 616 diode_w1
xdiode_183 0 1 616 diode_w1
xdiode_182 0 1 616 diode_w1
xdiode_181 0 1 616 diode_w1
xdiode_180 0 1 616 diode_w1
xfeed_6209 0 1 decap_w0
xfeed_6208 0 1 decap_w0
xfeed_6207 0 1 decap_w0
xfeed_6206 0 1 decap_w0
xfeed_6205 0 1 decap_w0
xfeed_6204 0 1 tie
xfeed_6203 0 1 decap_w0
xfeed_6202 0 1 decap_w0
xfeed_6201 0 1 decap_w0
xfeed_6200 0 1 decap_w0
xfeed_5599 0 1 decap_w0
xfeed_5597 0 1 decap_w0
xfeed_5596 0 1 decap_w0
xfeed_5594 0 1 decap_w0
xfeed_5593 0 1 decap_w0
xfeed_5592 0 1 decap_w0
xfeed_5591 0 1 decap_w0
xfeed_5590 0 1 decap_w0
xfeed_1289 0 1 decap_w0
xfeed_1288 0 1 decap_w0
xfeed_1287 0 1 decap_w0
xfeed_1286 0 1 decap_w0
xfeed_1285 0 1 decap_w0
xfeed_1284 0 1 decap_w0
xfeed_1283 0 1 decap_w0
xfeed_1282 0 1 decap_w0
xfeed_1281 0 1 decap_w0
xfeed_1280 0 1 decap_w0
xsubckt_746_nand2_x0 0 1 1720 1722 1721 nand2_x0
xfeed_12419 0 1 decap_w0
xfeed_12418 0 1 decap_w0
xfeed_12417 0 1 decap_w0
xfeed_12416 0 1 decap_w0
xfeed_12415 0 1 decap_w0
xfeed_12414 0 1 decap_w0
xfeed_12413 0 1 decap_w0
xfeed_12412 0 1 decap_w0
xfeed_12411 0 1 decap_w0
xfeed_12410 0 1 decap_w0
xsubckt_1250_nand2_x0 0 1 1330 665 661 nand2_x0
xsubckt_925_mux2_x1 0 1 1891 1586 2031 1579 mux2_x1
xsubckt_402_mux2_x1 0 1 347 2013 1985 1952 mux2_x1
xsubckt_1336_nand3_x0 0 1 1251 2058 666 657 nand3_x0
xdiode_197 0 1 775 diode_w1
xdiode_196 0 1 775 diode_w1
xdiode_195 0 1 774 diode_w1
xdiode_194 0 1 774 diode_w1
xdiode_193 0 1 773 diode_w1
xdiode_192 0 1 773 diode_w1
xdiode_191 0 1 773 diode_w1
xdiode_190 0 1 773 diode_w1
xfeed_6219 0 1 decap_w0
xfeed_6218 0 1 decap_w0
xfeed_6217 0 1 decap_w0
xfeed_6216 0 1 decap_w0
xfeed_6215 0 1 decap_w0
xfeed_6214 0 1 decap_w0
xfeed_6213 0 1 decap_w0
xfeed_6211 0 1 tie
xfeed_6210 0 1 decap_w0
xfeed_1299 0 1 decap_w0
xfeed_1298 0 1 decap_w0
xfeed_1297 0 1 decap_w0
xfeed_1296 0 1 decap_w0
xfeed_1295 0 1 decap_w0
xfeed_1294 0 1 decap_w0
xfeed_1293 0 1 decap_w0
xfeed_1292 0 1 decap_w0
xfeed_1291 0 1 decap_w0
xfeed_1290 0 1 decap_w0
xsubckt_1057_and4_x1 0 1 1485 645 623 525 519 and4_x1
xsubckt_1751_and21nor_x0 0 1 843 888 885 882 and21nor_x0
xdiode_199 0 1 775 diode_w1
xdiode_198 0 1 775 diode_w1
xfeed_12429 0 1 decap_w0
xfeed_12428 0 1 decap_w0
xfeed_12427 0 1 decap_w0
xfeed_12426 0 1 decap_w0
xfeed_12425 0 1 decap_w0
xfeed_12424 0 1 decap_w0
xfeed_12423 0 1 decap_w0
xfeed_12422 0 1 decap_w0
xfeed_12421 0 1 decap_w0
xfeed_12420 0 1 decap_w0
xsubckt_1245_mux2_x1 0 1 1816 2100 2067 1334 mux2_x1
xsubckt_892_nexor2_x0 0 1 1594 762 1597 nexor2_x0
xsubckt_208_nand2_x0 0 1 546 558 548 nand2_x0
xfeed_6229 0 1 decap_w0
xfeed_6228 0 1 decap_w0
xfeed_6227 0 1 tie
xfeed_6226 0 1 decap_w0
xfeed_6225 0 1 decap_w0
xfeed_6224 0 1 decap_w0
xfeed_6223 0 1 tie
xfeed_6222 0 1 decap_w0
xfeed_6221 0 1 decap_w0
xfeed_6220 0 1 decap_w0
xsubckt_883_nexor2_x0 0 1 1601 1604 1602 nexor2_x0
xsubckt_781_and21nor_x0 0 1 1690 1767 1778 1782 and21nor_x0
xsubckt_192_nand4_x0 0 1 566 716 1924 599 568 nand4_x0
xsubckt_624_or21nand_x0 0 1 2080 134 141 206 or21nand_x0
xsubckt_1676_mux2_x1 0 1 918 923 919 929 mux2_x1
xfeed_12439 0 1 decap_w0
xfeed_12438 0 1 decap_w0
xfeed_12437 0 1 decap_w0
xfeed_12436 0 1 decap_w0
xfeed_12435 0 1 decap_w0
xfeed_12434 0 1 decap_w0
xfeed_12433 0 1 decap_w0
xfeed_12432 0 1 decap_w0
xfeed_12431 0 1 decap_w0
xfeed_12430 0 1 decap_w0
xfeed_11909 0 1 decap_w0
xfeed_11908 0 1 decap_w0
xfeed_11907 0 1 decap_w0
xfeed_11906 0 1 decap_w0
xfeed_11905 0 1 decap_w0
xfeed_11904 0 1 decap_w0
xfeed_11903 0 1 decap_w0
xfeed_11902 0 1 decap_w0
xfeed_11901 0 1 decap_w0
xfeed_11900 0 1 decap_w0
xsubckt_865_nexor2_x0 0 1 1617 1964 2054 nexor2_x0
xsubckt_1686_nor3_x0 0 1 908 915 912 911 nor3_x0
xfeed_6239 0 1 decap_w0
xfeed_6238 0 1 decap_w0
xfeed_6237 0 1 decap_w0
xfeed_6236 0 1 decap_w0
xfeed_6235 0 1 tie
xfeed_6234 0 1 decap_w0
xfeed_6233 0 1 decap_w0
xfeed_6231 0 1 tie
xfeed_6230 0 1 decap_w0
xfeed_5709 0 1 decap_w0
xfeed_5707 0 1 decap_w0
xfeed_5706 0 1 decap_w0
xfeed_5705 0 1 decap_w0
xfeed_5704 0 1 tie
xfeed_5703 0 1 decap_w0
xfeed_5702 0 1 decap_w0
xfeed_5701 0 1 decap_w0
xfeed_5700 0 1 decap_w0
xsubckt_1149_mux2_x1 0 1 1835 1411 2012 1413 mux2_x1
xsubckt_1135_nand4_x0 0 1 1423 758 710 610 581 nand4_x0
xsubckt_984_and4_x1 0 1 1543 638 632 622 1544 and4_x1
xsubckt_1580_nand2_x0 0 1 1014 1018 1016 nand2_x0
xsubckt_1670_nand2_x0 0 1 924 927 926 nand2_x0
xfeed_12449 0 1 decap_w0
xfeed_12448 0 1 decap_w0
xfeed_12447 0 1 decap_w0
xfeed_12446 0 1 decap_w0
xfeed_12445 0 1 decap_w0
xfeed_12444 0 1 decap_w0
xfeed_12443 0 1 decap_w0
xfeed_12442 0 1 decap_w0
xfeed_12441 0 1 decap_w0
xfeed_12440 0 1 decap_w0
xfeed_11919 0 1 decap_w0
xfeed_11918 0 1 decap_w0
xfeed_11917 0 1 decap_w0
xfeed_11916 0 1 decap_w0
xfeed_11915 0 1 decap_w0
xfeed_11914 0 1 decap_w0
xfeed_11913 0 1 decap_w0
xfeed_11912 0 1 decap_w0
xfeed_11911 0 1 decap_w0
xfeed_11910 0 1 decap_w0
xsubckt_747_nor3_x0 0 1 1719 1724 1723 1720 nor3_x0
xsubckt_1576_nand3_x0 0 1 1018 1971 678 595 nand3_x0
xfeed_6249 0 1 decap_w0
xfeed_6248 0 1 decap_w0
xfeed_6247 0 1 decap_w0
xfeed_6246 0 1 decap_w0
xfeed_6245 0 1 tie
xfeed_6244 0 1 decap_w0
xfeed_6243 0 1 decap_w0
xfeed_6242 0 1 decap_w0
xfeed_6241 0 1 decap_w0
xfeed_6240 0 1 decap_w0
xfeed_5719 0 1 decap_w0
xfeed_5718 0 1 decap_w0
xfeed_5717 0 1 decap_w0
xfeed_5716 0 1 decap_w0
xfeed_5715 0 1 decap_w0
xfeed_5713 0 1 decap_w0
xfeed_5712 0 1 decap_w0
xfeed_5711 0 1 decap_w0
xfeed_5710 0 1 decap_w0
xfeed_1409 0 1 decap_w0
xfeed_1408 0 1 decap_w0
xfeed_1407 0 1 decap_w0
xfeed_1406 0 1 tie
xfeed_1405 0 1 decap_w0
xfeed_1404 0 1 decap_w0
xfeed_1403 0 1 decap_w0
xfeed_1402 0 1 decap_w0
xfeed_1401 0 1 decap_w0
xfeed_1400 0 1 decap_w0
xsubckt_122_mux2_x1 0 1 646 1992 2001 1986 mux2_x1
xsubckt_483_and3_x1 0 1 267 1917 771 583 and3_x1
xsubckt_628_nand2_x0 0 1 130 2042 172 nand2_x0
xsubckt_1366_and2_x1 0 1 1223 1229 1224 and2_x1
xfeed_12459 0 1 decap_w0
xfeed_12458 0 1 decap_w0
xfeed_12457 0 1 decap_w0
xfeed_12456 0 1 decap_w0
xfeed_12455 0 1 decap_w0
xfeed_12454 0 1 decap_w0
xfeed_12453 0 1 decap_w0
xfeed_12452 0 1 decap_w0
xfeed_12451 0 1 decap_w0
xfeed_12450 0 1 decap_w0
xfeed_11929 0 1 decap_w0
xfeed_11928 0 1 decap_w0
xfeed_11927 0 1 decap_w0
xfeed_11926 0 1 decap_w0
xfeed_11925 0 1 decap_w0
xfeed_11924 0 1 decap_w0
xfeed_11923 0 1 decap_w0
xfeed_11922 0 1 decap_w0
xfeed_11921 0 1 decap_w0
xfeed_11920 0 1 decap_w0
xsubckt_1485_or21nand_x0 0 1 1111 1114 1118 759 or21nand_x0
xfeed_6259 0 1 decap_w0
xfeed_6258 0 1 decap_w0
xfeed_6257 0 1 decap_w0
xfeed_6256 0 1 decap_w0
xfeed_6255 0 1 decap_w0
xfeed_6254 0 1 decap_w0
xfeed_6253 0 1 decap_w0
xfeed_6252 0 1 decap_w0
xfeed_6251 0 1 decap_w0
xfeed_6250 0 1 decap_w0
xfeed_5729 0 1 decap_w0
xfeed_5728 0 1 decap_w0
xfeed_5727 0 1 decap_w0
xfeed_5726 0 1 decap_w0
xfeed_5725 0 1 decap_w0
xfeed_5724 0 1 decap_w0
xfeed_5723 0 1 decap_w0
xfeed_5722 0 1 tie
xfeed_5721 0 1 decap_w0
xfeed_5720 0 1 decap_w0
xfeed_1419 0 1 decap_w0
xfeed_1418 0 1 decap_w0
xfeed_1417 0 1 decap_w0
xfeed_1416 0 1 decap_w0
xfeed_1415 0 1 decap_w0
xfeed_1414 0 1 decap_w0
xfeed_1413 0 1 decap_w0
xfeed_1412 0 1 decap_w0
xfeed_1411 0 1 decap_w0
xfeed_1410 0 1 tie
xsubckt_1134_and4_x1 0 1 1424 758 710 610 581 and4_x1
xsubckt_1038_nand3_x0 0 1 1499 643 533 1527 nand3_x0
xsubckt_365_and4_x1 0 1 384 660 656 655 527 and4_x1
xsubckt_1683_and3_x1 0 1 911 1070 927 926 and3_x1
xsubckt_1851_dff_x1 0 1 2027 1887 32 dff_x1
xfeed_12469 0 1 decap_w0
xfeed_12468 0 1 decap_w0
xfeed_12467 0 1 decap_w0
xfeed_12466 0 1 decap_w0
xfeed_12465 0 1 decap_w0
xfeed_12464 0 1 decap_w0
xfeed_12463 0 1 decap_w0
xfeed_12462 0 1 tie
xfeed_12461 0 1 decap_w0
xfeed_12460 0 1 decap_w0
xfeed_11939 0 1 decap_w0
xfeed_11938 0 1 decap_w0
xfeed_11937 0 1 decap_w0
xfeed_11936 0 1 decap_w0
xfeed_11935 0 1 decap_w0
xfeed_11934 0 1 decap_w0
xfeed_11933 0 1 decap_w0
xfeed_11932 0 1 decap_w0
xfeed_11931 0 1 tie
xfeed_11930 0 1 decap_w0
xsubckt_910_mux2_x1 0 1 1905 1618 2045 1580 mux2_x1
xsubckt_1446_nor2_x0 0 1 1149 1154 1150 nor2_x0
xsubckt_1853_dff_x1 0 1 2025 1885 35 dff_x1
xsubckt_1855_dff_x1 0 1 2023 1883 32 dff_x1
xsubckt_1857_dff_x1 0 1 1983 1881 54 dff_x1
xfeed_6269 0 1 tie
xfeed_6268 0 1 decap_w0
xfeed_6267 0 1 decap_w0
xfeed_6266 0 1 decap_w0
xfeed_6265 0 1 tie
xfeed_6264 0 1 decap_w0
xfeed_6263 0 1 decap_w0
xfeed_6262 0 1 decap_w0
xfeed_6261 0 1 decap_w0
xfeed_6260 0 1 decap_w0
xfeed_5739 0 1 decap_w0
xfeed_5738 0 1 decap_w0
xfeed_5737 0 1 decap_w0
xfeed_5736 0 1 decap_w0
xfeed_5735 0 1 decap_w0
xfeed_5734 0 1 decap_w0
xfeed_5733 0 1 decap_w0
xfeed_5732 0 1 decap_w0
xfeed_5731 0 1 decap_w0
xfeed_5730 0 1 decap_w0
xfeed_1429 0 1 decap_w0
xfeed_1428 0 1 decap_w0
xfeed_1427 0 1 decap_w0
xfeed_1426 0 1 decap_w0
xfeed_1425 0 1 tie
xfeed_1424 0 1 decap_w0
xfeed_1423 0 1 decap_w0
xfeed_1422 0 1 decap_w0
xfeed_1421 0 1 decap_w0
xfeed_1420 0 1 decap_w0
xsubckt_1104_or2_x1 0 1 1847 1457 1444 or2_x1
xsubckt_1859_dff_x1 0 1 1954 1880 67 dff_x1
xfeed_12479 0 1 decap_w0
xfeed_12478 0 1 decap_w0
xfeed_12477 0 1 decap_w0
xfeed_12476 0 1 decap_w0
xfeed_12475 0 1 decap_w0
xfeed_12474 0 1 decap_w0
xfeed_12473 0 1 decap_w0
xfeed_12472 0 1 decap_w0
xfeed_12471 0 1 decap_w0
xfeed_12470 0 1 decap_w0
xfeed_11947 0 1 decap_w0
xfeed_11946 0 1 decap_w0
xfeed_11945 0 1 decap_w0
xfeed_11944 0 1 tie
xfeed_11943 0 1 decap_w0
xfeed_11942 0 1 decap_w0
xfeed_11941 0 1 decap_w0
xfeed_11940 0 1 decap_w0
xsubckt_269_and4_x1 0 1 479 714 1928 678 589 and4_x1
xsubckt_341_nand2_x0 0 1 407 687 408 nand2_x0
xfeed_11949 0 1 decap_w0
xfeed_11948 0 1 decap_w0
xfeed_6279 0 1 decap_w0
xfeed_6278 0 1 tie
xfeed_6277 0 1 decap_w0
xfeed_6276 0 1 decap_w0
xfeed_6275 0 1 decap_w0
xfeed_6274 0 1 decap_w0
xfeed_6273 0 1 tie
xfeed_6272 0 1 decap_w0
xfeed_6271 0 1 decap_w0
xfeed_6270 0 1 decap_w0
xfeed_5749 0 1 decap_w0
xfeed_5748 0 1 decap_w0
xfeed_5747 0 1 decap_w0
xfeed_5745 0 1 decap_w0
xfeed_5744 0 1 decap_w0
xfeed_5743 0 1 decap_w0
xfeed_5742 0 1 decap_w0
xfeed_5741 0 1 decap_w0
xfeed_5740 0 1 tie
xfeed_1439 0 1 tie
xfeed_1438 0 1 decap_w0
xfeed_1437 0 1 decap_w0
xfeed_1436 0 1 decap_w0
xfeed_1435 0 1 decap_w0
xfeed_1434 0 1 decap_w0
xfeed_1433 0 1 decap_w0
xfeed_1432 0 1 tie
xfeed_1431 0 1 decap_w0
xsubckt_1199_or3_x1 0 1 1365 1371 1370 1366 or3_x1
xsubckt_1090_and2_x1 0 1 1457 1946 1575 and2_x1
xsubckt_1017_nand4_x0 0 1 1514 637 633 622 1515 nand4_x0
xsubckt_944_nand4_x0 0 1 1573 650 644 533 1576 nand4_x0
xsubckt_766_and2_x1 0 1 1703 2048 1748 and2_x1
xsubckt_161_nand2_x0 0 1 600 610 603 nand2_x0
xsubckt_1552_nand2_x0 0 1 1042 1044 1043 nand2_x0
xsubckt_1785_or21nand_x0 0 1 809 1036 1035 1032 or21nand_x0
xfeed_12489 0 1 decap_w0
xfeed_12488 0 1 decap_w0
xfeed_12487 0 1 decap_w0
xfeed_12486 0 1 decap_w0
xfeed_12485 0 1 decap_w0
xfeed_12484 0 1 decap_w0
xfeed_12483 0 1 decap_w0
xfeed_12482 0 1 decap_w0
xfeed_12481 0 1 decap_w0
xfeed_12480 0 1 decap_w0
xfeed_11954 0 1 decap_w0
xfeed_11953 0 1 decap_w0
xfeed_11952 0 1 decap_w0
xfeed_11951 0 1 tie
xfeed_11950 0 1 decap_w0
xsubckt_1086_and2_x1 0 1 1459 1461 1460 and2_x1
xsubckt_880_and21nor_x0 0 1 1604 1609 1608 1615 and21nor_x0
xsubckt_239_and2_x1 0 1 512 514 513 and2_x1
xsubckt_1746_and21nor_x0 0 1 848 860 858 855 and21nor_x0
xfeed_11959 0 1 decap_w0
xfeed_11958 0 1 decap_w0
xfeed_11957 0 1 decap_w0
xfeed_11956 0 1 decap_w0
xfeed_11955 0 1 decap_w0
xfeed_6289 0 1 decap_w0
xfeed_6288 0 1 decap_w0
xfeed_6287 0 1 decap_w0
xfeed_6286 0 1 decap_w0
xfeed_6285 0 1 decap_w0
xfeed_6284 0 1 decap_w0
xfeed_6283 0 1 decap_w0
xfeed_6282 0 1 decap_w0
xfeed_6281 0 1 decap_w0
xfeed_6280 0 1 decap_w0
xfeed_5759 0 1 decap_w0
xfeed_5758 0 1 decap_w0
xfeed_5757 0 1 tie
xfeed_5756 0 1 decap_w0
xfeed_5755 0 1 decap_w0
xfeed_5754 0 1 decap_w0
xfeed_5753 0 1 decap_w0
xfeed_5752 0 1 decap_w0
xfeed_5751 0 1 decap_w0
xfeed_5750 0 1 decap_w0
xfeed_1449 0 1 decap_w0
xfeed_1448 0 1 decap_w0
xfeed_1447 0 1 decap_w0
xfeed_1446 0 1 decap_w0
xfeed_1445 0 1 decap_w0
xfeed_1444 0 1 decap_w0
xfeed_1443 0 1 decap_w0
xfeed_1442 0 1 decap_w0
xfeed_1441 0 1 decap_w0
xfeed_1440 0 1 decap_w0
xsubckt_534_and4_x1 0 1 219 223 222 221 220 and4_x1
xsubckt_560_and3_x1 0 1 195 198 197 196 and3_x1
xsubckt_1282_nand2_x0 0 1 1300 775 1974 nand2_x0
xsubckt_1621_nand3_x0 0 1 973 1070 989 987 nand3_x0
xfeed_13109 0 1 decap_w0
xfeed_13108 0 1 decap_w0
xfeed_13107 0 1 decap_w0
xfeed_13106 0 1 decap_w0
xfeed_13105 0 1 decap_w0
xfeed_13104 0 1 decap_w0
xfeed_13103 0 1 tie
xfeed_13102 0 1 decap_w0
xfeed_13101 0 1 decap_w0
xfeed_13100 0 1 decap_w0
xfeed_12499 0 1 decap_w0
xfeed_12498 0 1 decap_w0
xfeed_12497 0 1 decap_w0
xfeed_12496 0 1 decap_w0
xfeed_12495 0 1 tie
xfeed_12494 0 1 decap_w0
xfeed_12493 0 1 decap_w0
xfeed_12492 0 1 decap_w0
xfeed_12491 0 1 decap_w0
xfeed_12490 0 1 decap_w0
xfeed_11961 0 1 decap_w0
xfeed_11960 0 1 decap_w0
xsubckt_1144_nor3_x0 0 1 1415 1940 1958 1936 nor3_x0
xsubckt_619_or21nand_x0 0 1 138 1995 436 167 or21nand_x0
xfeed_11969 0 1 decap_w0
xfeed_11968 0 1 decap_w0
xfeed_11967 0 1 decap_w0
xfeed_11966 0 1 decap_w0
xfeed_11965 0 1 tie
xfeed_11964 0 1 decap_w0
xfeed_11963 0 1 decap_w0
xfeed_11962 0 1 decap_w0
xfeed_6299 0 1 decap_w0
xfeed_6298 0 1 decap_w0
xfeed_6297 0 1 tie
xfeed_6296 0 1 decap_w0
xfeed_6295 0 1 decap_w0
xfeed_6294 0 1 decap_w0
xfeed_6293 0 1 tie
xfeed_6292 0 1 decap_w0
xfeed_6291 0 1 decap_w0
xfeed_6290 0 1 decap_w0
xfeed_5769 0 1 decap_w0
xfeed_5768 0 1 decap_w0
xfeed_5767 0 1 tie
xfeed_5766 0 1 decap_w0
xfeed_5764 0 1 decap_w0
xfeed_5763 0 1 decap_w0
xfeed_5762 0 1 tie
xfeed_5761 0 1 decap_w0
xfeed_5760 0 1 decap_w0
xfeed_1459 0 1 decap_w0
xfeed_1458 0 1 decap_w0
xfeed_1457 0 1 decap_w0
xfeed_1456 0 1 decap_w0
xfeed_1455 0 1 decap_w0
xfeed_1454 0 1 decap_w0
xfeed_1453 0 1 decap_w0
xfeed_1452 0 1 decap_w0
xfeed_1451 0 1 decap_w0
xfeed_1450 0 1 decap_w0
xsubckt_761_nand2_x0 0 1 1707 1999 1746 nand2_x0
xsubckt_92_mux2_x1 0 1 693 700 699 774 mux2_x1
xfeed_13119 0 1 decap_w0
xfeed_13118 0 1 decap_w0
xfeed_13117 0 1 decap_w0
xfeed_13116 0 1 decap_w0
xfeed_13115 0 1 decap_w0
xfeed_13114 0 1 decap_w0
xfeed_13113 0 1 decap_w0
xfeed_13112 0 1 decap_w0
xfeed_13111 0 1 decap_w0
xfeed_13110 0 1 tie
xsubckt_667_nand3_x0 0 1 94 2023 184 176 nand3_x0
xsubckt_375_and21nor_x0 0 1 374 377 376 535 and21nor_x0
xsubckt_581_nand2_x0 0 1 174 2037 175 nand2_x0
xfeed_11979 0 1 decap_w0
xfeed_11978 0 1 decap_w0
xfeed_11977 0 1 decap_w0
xfeed_11976 0 1 tie
xfeed_11975 0 1 decap_w0
xfeed_11974 0 1 decap_w0
xfeed_11973 0 1 decap_w0
xfeed_11972 0 1 tie
xfeed_11971 0 1 decap_w0
xfeed_11970 0 1 decap_w0
xfeed_5779 0 1 decap_w0
xfeed_5778 0 1 decap_w0
xfeed_5777 0 1 decap_w0
xfeed_5776 0 1 decap_w0
xfeed_5775 0 1 decap_w0
xfeed_5774 0 1 tie
xfeed_5773 0 1 decap_w0
xfeed_5772 0 1 decap_w0
xfeed_5771 0 1 decap_w0
xfeed_5770 0 1 decap_w0
xfeed_1469 0 1 decap_w0
xfeed_1468 0 1 decap_w0
xfeed_1467 0 1 decap_w0
xfeed_1466 0 1 decap_w0
xfeed_1465 0 1 decap_w0
xfeed_1464 0 1 decap_w0
xfeed_1463 0 1 decap_w0
xfeed_1462 0 1 decap_w0
xfeed_1461 0 1 decap_w0
xfeed_1460 0 1 decap_w0
xsubckt_1207_and4_x1 0 1 1357 414 193 1769 1358 and4_x1
xsubckt_313_nand2_x0 0 1 435 681 447 nand2_x0
xsubckt_88_mux2_x1 0 1 695 704 703 774 mux2_x1
xsubckt_412_and2_x1 0 1 337 340 338 and2_x1
xsubckt_1614_nand2_x0 0 1 980 1101 982 nand2_x0
xfeed_13129 0 1 decap_w0
xfeed_13128 0 1 decap_w0
xfeed_13127 0 1 decap_w0
xfeed_13126 0 1 decap_w0
xfeed_13125 0 1 decap_w0
xfeed_13124 0 1 decap_w0
xfeed_13123 0 1 decap_w0
xfeed_13122 0 1 decap_w0
xfeed_13121 0 1 decap_w0
xfeed_13120 0 1 decap_w0
xsubckt_1081_nand3_x0 0 1 1463 426 1465 1464 nand3_x0
xsubckt_895_and3_x1 0 1 1592 1962 1964 2055 and3_x1
xsubckt_223_nand2_x0 0 1 528 785 1998 nand2_x0
xsubckt_221_or21nand_x0 0 1 530 661 651 646 or21nand_x0
xsubckt_133_nand2_x0 0 1 635 785 2002 nand2_x0
xsubckt_346_and4_x1 0 1 402 1917 771 568 405 and4_x1
xsubckt_372_and3_x1 0 1 377 609 557 447 and3_x1
xsubckt_486_and2_x1 0 1 264 469 422 and2_x1
xsubckt_1524_nand2_x0 0 1 1072 1081 1077 nand2_x0
xfeed_11989 0 1 decap_w0
xfeed_11988 0 1 decap_w0
xfeed_11987 0 1 decap_w0
xfeed_11986 0 1 decap_w0
xfeed_11985 0 1 decap_w0
xfeed_11984 0 1 decap_w0
xfeed_11983 0 1 decap_w0
xfeed_11982 0 1 decap_w0
xfeed_11981 0 1 decap_w0
xfeed_11980 0 1 decap_w0
xfeed_5789 0 1 decap_w0
xfeed_5788 0 1 decap_w0
xfeed_5787 0 1 decap_w0
xfeed_5786 0 1 decap_w0
xfeed_5785 0 1 decap_w0
xfeed_5784 0 1 decap_w0
xfeed_5783 0 1 decap_w0
xfeed_5782 0 1 tie
xfeed_5780 0 1 decap_w0
xfeed_1479 0 1 decap_w0
xfeed_1478 0 1 decap_w0
xfeed_1477 0 1 decap_w0
xfeed_1476 0 1 decap_w0
xfeed_1475 0 1 decap_w0
xfeed_1474 0 1 decap_w0
xfeed_1473 0 1 decap_w0
xfeed_1472 0 1 tie
xfeed_1471 0 1 decap_w0
xfeed_1470 0 1 decap_w0
xsubckt_703_and4_x1 0 1 1761 1927 1925 711 674 and4_x1
xsubckt_1344_nand2_x0 0 1 1243 1917 1244 nand2_x0
xfeed_13139 0 1 decap_w0
xfeed_13138 0 1 decap_w0
xfeed_13137 0 1 decap_w0
xfeed_13136 0 1 decap_w0
xfeed_13135 0 1 decap_w0
xfeed_13134 0 1 decap_w0
xfeed_13133 0 1 decap_w0
xfeed_13132 0 1 decap_w0
xfeed_13131 0 1 decap_w0
xfeed_13130 0 1 decap_w0
xfeed_12609 0 1 decap_w0
xfeed_12608 0 1 decap_w0
xfeed_12607 0 1 decap_w0
xfeed_12606 0 1 decap_w0
xfeed_12605 0 1 decap_w0
xfeed_12604 0 1 decap_w0
xfeed_12603 0 1 decap_w0
xfeed_12602 0 1 decap_w0
xfeed_12601 0 1 decap_w0
xfeed_12600 0 1 decap_w0
xsubckt_806_or2_x1 0 1 2091 1674 1668 or2_x1
xsubckt_470_nand3_x0 0 1 280 686 617 451 nand3_x0
xfeed_11999 0 1 decap_w0
xfeed_11998 0 1 decap_w0
xfeed_11997 0 1 decap_w0
xfeed_11996 0 1 decap_w0
xfeed_11995 0 1 decap_w0
xfeed_11994 0 1 decap_w0
xfeed_11993 0 1 decap_w0
xfeed_11992 0 1 decap_w0
xfeed_11991 0 1 decap_w0
xfeed_11990 0 1 decap_w0
xfeed_6409 0 1 decap_w0
xfeed_6408 0 1 decap_w0
xfeed_6407 0 1 decap_w0
xfeed_6406 0 1 tie
xfeed_6405 0 1 decap_w0
xfeed_6404 0 1 decap_w0
xfeed_6403 0 1 decap_w0
xfeed_6402 0 1 decap_w0
xfeed_6401 0 1 tie
xfeed_6400 0 1 decap_w0
xfeed_5799 0 1 decap_w0
xfeed_5798 0 1 decap_w0
xfeed_5797 0 1 decap_w0
xfeed_5796 0 1 decap_w0
xfeed_5795 0 1 decap_w0
xfeed_5794 0 1 decap_w0
xfeed_5793 0 1 decap_w0
xfeed_5792 0 1 decap_w0
xfeed_5790 0 1 decap_w0
xfeed_1489 0 1 tie
xfeed_1488 0 1 decap_w0
xfeed_1487 0 1 decap_w0
xfeed_1486 0 1 decap_w0
xfeed_1485 0 1 decap_w0
xfeed_1484 0 1 decap_w0
xfeed_1483 0 1 decap_w0
xfeed_1482 0 1 decap_w0
xfeed_1481 0 1 decap_w0
xfeed_1480 0 1 decap_w0
xsubckt_799_and3_x1 0 1 1674 1967 1749 1739 and3_x1
xsubckt_751_and2_x1 0 1 1716 2050 1748 and2_x1
xsubckt_675_and21nor_x0 0 1 86 749 449 410 and21nor_x0
xsubckt_466_nand4_x0 0 1 284 714 1928 712 589 nand4_x0
xsubckt_1309_or2_x1 0 1 1275 1280 1277 or2_x1
xsubckt_1520_and2_x1 0 1 1076 1082 1078 and2_x1
xsubckt_1608_and2_x1 0 1 986 989 987 and2_x1
xsubckt_1734_mux2_x1 0 1 860 900 862 1142 mux2_x1
xfeed_13149 0 1 decap_w0
xfeed_13148 0 1 decap_w0
xfeed_13147 0 1 decap_w0
xfeed_13146 0 1 decap_w0
xfeed_13145 0 1 decap_w0
xfeed_13144 0 1 decap_w0
xfeed_13143 0 1 decap_w0
xfeed_13142 0 1 decap_w0
xfeed_13141 0 1 decap_w0
xfeed_13140 0 1 decap_w0
xfeed_12619 0 1 decap_w0
xfeed_12618 0 1 decap_w0
xfeed_12617 0 1 tie
xfeed_12616 0 1 decap_w0
xfeed_12615 0 1 decap_w0
xfeed_12614 0 1 tie
xfeed_12613 0 1 decap_w0
xfeed_12612 0 1 decap_w0
xfeed_12611 0 1 decap_w0
xfeed_12610 0 1 decap_w0
xsubckt_1159_and2_x1 0 1 1402 1940 768 and2_x1
xsubckt_819_nand3_x0 0 1 1656 2070 680 489 nand3_x0
xsubckt_733_nand2_x0 0 1 1732 152 1766 nand2_x0
xsubckt_643_nand2_x0 0 1 116 118 117 nand2_x0
xsubckt_618_or21nand_x0 0 1 139 2051 601 163 or21nand_x0
xsubckt_1483_or21nand_x0 0 1 1113 1628 1116 689 or21nand_x0
xfeed_6419 0 1 decap_w0
xfeed_6418 0 1 decap_w0
xfeed_6417 0 1 decap_w0
xfeed_6416 0 1 decap_w0
xfeed_6415 0 1 decap_w0
xfeed_6414 0 1 decap_w0
xfeed_6412 0 1 decap_w0
xfeed_6411 0 1 decap_w0
xfeed_6410 0 1 decap_w0
xfeed_2109 0 1 decap_w0
xfeed_2108 0 1 decap_w0
xfeed_2107 0 1 decap_w0
xfeed_2106 0 1 decap_w0
xfeed_2105 0 1 decap_w0
xfeed_2104 0 1 decap_w0
xfeed_2103 0 1 decap_w0
xfeed_2102 0 1 decap_w0
xfeed_2101 0 1 decap_w0
xfeed_2100 0 1 decap_w0
xfeed_1499 0 1 decap_w0
xfeed_1498 0 1 decap_w0
xfeed_1497 0 1 decap_w0
xfeed_1496 0 1 decap_w0
xfeed_1495 0 1 decap_w0
xfeed_1494 0 1 decap_w0
xfeed_1493 0 1 decap_w0
xfeed_1492 0 1 decap_w0
xfeed_1491 0 1 decap_w0
xfeed_1490 0 1 decap_w0
xsubckt_1129_nexor2_x0 0 1 1428 759 1429 nexor2_x0
xsubckt_298_and2_x1 0 1 450 616 451 and2_x1
xsubckt_286_nand4_x0 0 1 462 712 1926 599 589 nand4_x0
xsubckt_553_nand2_x0 0 1 201 1921 202 nand2_x0
xfeed_13159 0 1 decap_w0
xfeed_13158 0 1 decap_w0
xfeed_13157 0 1 decap_w0
xfeed_13156 0 1 tie
xfeed_13155 0 1 decap_w0
xfeed_13154 0 1 decap_w0
xfeed_13153 0 1 decap_w0
xfeed_13152 0 1 decap_w0
xfeed_13151 0 1 decap_w0
xfeed_13150 0 1 decap_w0
xfeed_12629 0 1 decap_w0
xfeed_12628 0 1 decap_w0
xfeed_12627 0 1 decap_w0
xfeed_12626 0 1 decap_w0
xfeed_12625 0 1 decap_w0
xfeed_12624 0 1 decap_w0
xfeed_12623 0 1 tie
xfeed_12622 0 1 decap_w0
xfeed_12621 0 1 decap_w0
xfeed_12620 0 1 decap_w0
xsubckt_1115_mux2_x1 0 1 1842 2000 1991 1438 mux2_x1
xsubckt_718_or21nand_x0 0 1 1746 569 459 614 or21nand_x0
xsubckt_463_nand2_x0 0 1 287 609 581 nand2_x0
xsubckt_515_and4_x1 0 1 236 507 496 432 237 and4_x1
xsubckt_639_nand3_x0 0 1 120 2017 184 177 nand3_x0
xsubckt_1764_nand2_x0 0 1 830 1964 548 nand2_x0
xfeed_6429 0 1 decap_w0
xfeed_6428 0 1 decap_w0
xfeed_6427 0 1 decap_w0
xfeed_6426 0 1 decap_w0
xfeed_6425 0 1 decap_w0
xfeed_6424 0 1 decap_w0
xfeed_6423 0 1 decap_w0
xfeed_6422 0 1 decap_w0
xfeed_6421 0 1 decap_w0
xfeed_6420 0 1 tie
xfeed_2119 0 1 decap_w0
xfeed_2118 0 1 decap_w0
xfeed_2117 0 1 decap_w0
xfeed_2116 0 1 decap_w0
xfeed_2115 0 1 decap_w0
xfeed_2114 0 1 decap_w0
xfeed_2113 0 1 decap_w0
xfeed_2112 0 1 decap_w0
xfeed_2111 0 1 decap_w0
xfeed_2110 0 1 decap_w0
xfeed_13169 0 1 decap_w0
xfeed_13168 0 1 tie
xfeed_13167 0 1 decap_w0
xfeed_13166 0 1 decap_w0
xfeed_13165 0 1 decap_w0
xfeed_13164 0 1 decap_w0
xfeed_13163 0 1 decap_w0
xfeed_13162 0 1 decap_w0
xfeed_13161 0 1 decap_w0
xfeed_13160 0 1 decap_w0
xfeed_12639 0 1 decap_w0
xfeed_12638 0 1 decap_w0
xfeed_12637 0 1 decap_w0
xfeed_12636 0 1 decap_w0
xfeed_12635 0 1 decap_w0
xfeed_12634 0 1 decap_w0
xfeed_12633 0 1 decap_w0
xfeed_12632 0 1 decap_w0
xfeed_12631 0 1 decap_w0
xfeed_12630 0 1 tie
xsubckt_1023_mux2_x1 0 1 1861 1511 1955 1576 mux2_x1
xsubckt_220_or21nand_x0 0 1 534 661 639 634 or21nand_x0
xsubckt_563_and2_x1 0 1 192 501 462 and2_x1
xsubckt_1584_nand2_x0 0 1 1010 1012 1011 nand2_x0
xfeed_6439 0 1 decap_w0
xfeed_6438 0 1 decap_w0
xfeed_6437 0 1 decap_w0
xfeed_6436 0 1 tie
xfeed_6435 0 1 decap_w0
xfeed_6434 0 1 decap_w0
xfeed_6433 0 1 decap_w0
xfeed_6432 0 1 decap_w0
xfeed_6431 0 1 decap_w0
xfeed_6430 0 1 decap_w0
xfeed_5909 0 1 decap_w0
xfeed_5908 0 1 decap_w0
xfeed_5907 0 1 decap_w0
xfeed_5906 0 1 decap_w0
xfeed_5905 0 1 decap_w0
xfeed_5904 0 1 decap_w0
xfeed_5903 0 1 decap_w0
xfeed_5902 0 1 decap_w0
xfeed_5901 0 1 decap_w0
xfeed_5900 0 1 decap_w0
xfeed_2129 0 1 decap_w0
xfeed_2128 0 1 decap_w0
xfeed_2127 0 1 decap_w0
xfeed_2126 0 1 decap_w0
xfeed_2125 0 1 decap_w0
xfeed_2124 0 1 decap_w0
xfeed_2123 0 1 decap_w0
xfeed_2122 0 1 decap_w0
xfeed_2121 0 1 decap_w0
xfeed_2120 0 1 decap_w0
xsubckt_189_nand3_x0 0 1 569 1925 711 571 nand3_x0
xfeed_13179 0 1 decap_w0
xfeed_13178 0 1 decap_w0
xfeed_13177 0 1 decap_w0
xfeed_13176 0 1 decap_w0
xfeed_13175 0 1 decap_w0
xfeed_13174 0 1 decap_w0
xfeed_13173 0 1 decap_w0
xfeed_13172 0 1 decap_w0
xfeed_13171 0 1 decap_w0
xfeed_13170 0 1 decap_w0
xfeed_12647 0 1 decap_w0
xfeed_12646 0 1 decap_w0
xfeed_12645 0 1 decap_w0
xfeed_12644 0 1 decap_w0
xfeed_12643 0 1 decap_w0
xfeed_12642 0 1 decap_w0
xfeed_12641 0 1 decap_w0
xfeed_12640 0 1 tie
xsubckt_1078_or21nand_x0 0 1 1466 1468 1467 1495 or21nand_x0
xsubckt_1019_mux2_x1 0 1 1863 1513 1938 1576 mux2_x1
xsubckt_442_nand3_x0 0 1 308 653 632 530 nand3_x0
xsubckt_1763_and2_x1 0 1 831 1964 548 and2_x1
xsubckt_1783_or21nand_x0 0 1 811 996 817 815 or21nand_x0
xsubckt_1900_dff_x1 0 1 1946 1847 67 dff_x1
xsubckt_1902_dff_x1 0 1 1994 1845 67 dff_x1
xfeed_101 0 1 decap_w0
xfeed_102 0 1 decap_w0
xfeed_103 0 1 decap_w0
xfeed_104 0 1 decap_w0
xfeed_105 0 1 decap_w0
xfeed_106 0 1 decap_w0
xfeed_107 0 1 decap_w0
xfeed_108 0 1 decap_w0
xfeed_12649 0 1 decap_w0
xfeed_12648 0 1 decap_w0
xfeed_6449 0 1 decap_w0
xfeed_6448 0 1 tie
xfeed_6447 0 1 decap_w0
xfeed_6446 0 1 decap_w0
xfeed_6444 0 1 decap_w0
xfeed_6443 0 1 decap_w0
xfeed_6442 0 1 decap_w0
xfeed_6441 0 1 decap_w0
xfeed_6440 0 1 decap_w0
xfeed_5919 0 1 decap_w0
xfeed_5918 0 1 decap_w0
xfeed_5917 0 1 decap_w0
xfeed_5916 0 1 decap_w0
xfeed_5915 0 1 decap_w0
xfeed_5914 0 1 decap_w0
xfeed_5913 0 1 decap_w0
xfeed_5912 0 1 decap_w0
xfeed_5911 0 1 decap_w0
xfeed_5910 0 1 decap_w0
xfeed_2139 0 1 decap_w0
xfeed_2138 0 1 decap_w0
xfeed_2137 0 1 decap_w0
xfeed_2136 0 1 decap_w0
xfeed_2135 0 1 decap_w0
xfeed_2134 0 1 decap_w0
xfeed_2133 0 1 decap_w0
xfeed_2132 0 1 decap_w0
xfeed_2131 0 1 decap_w0
xfeed_2130 0 1 decap_w0
xfeed_1609 0 1 decap_w0
xfeed_1608 0 1 decap_w0
xfeed_1607 0 1 decap_w0
xfeed_1606 0 1 decap_w0
xfeed_1605 0 1 decap_w0
xfeed_1604 0 1 decap_w0
xfeed_1603 0 1 decap_w0
xfeed_1602 0 1 decap_w0
xfeed_1601 0 1 decap_w0
xfeed_1600 0 1 decap_w0
xsubckt_802_and3_x1 0 1 1671 2072 679 490 and3_x1
xsubckt_262_nand3_x0 0 1 486 687 617 490 nand3_x0
xsubckt_327_and4_x1 0 1 421 716 1924 1927 713 and4_x1
xsubckt_438_nand4_x0 0 1 312 659 641 640 634 nand4_x0
xsubckt_1563_nand3_x0 0 1 1031 1070 1050 1048 nand3_x0
xsubckt_1904_dff_x1 0 1 1992 1843 67 dff_x1
xsubckt_1906_dff_x1 0 1 1990 1841 64 dff_x1
xfeed_13189 0 1 decap_w0
xfeed_13188 0 1 decap_w0
xfeed_13187 0 1 decap_w0
xfeed_13186 0 1 decap_w0
xfeed_13185 0 1 decap_w0
xfeed_13184 0 1 decap_w0
xfeed_13183 0 1 decap_w0
xfeed_13182 0 1 decap_w0
xfeed_13181 0 1 decap_w0
xfeed_13180 0 1 decap_w0
xfeed_12654 0 1 decap_w0
xfeed_12653 0 1 decap_w0
xfeed_12652 0 1 decap_w0
xfeed_12651 0 1 decap_w0
xfeed_12650 0 1 decap_w0
xsubckt_710_and3_x1 0 1 1754 587 579 493 and3_x1
xsubckt_615_nand2_x0 0 1 142 2043 172 nand2_x0
xsubckt_1807_mux2_x1 0 1 1795 2052 829 774 mux2_x1
xsubckt_1860_dff_x1 0 1 1953 1879 67 dff_x1
xsubckt_1862_dff_x1 0 1 1940 1877 64 dff_x1
xsubckt_1864_dff_x1 0 1 1959 1875 67 dff_x1
xsubckt_1908_dff_x1 0 1 1988 1839 67 dff_x1
xfeed_110 0 1 decap_w0
xfeed_111 0 1 decap_w0
xfeed_112 0 1 decap_w0
xfeed_113 0 1 decap_w0
xfeed_114 0 1 decap_w0
xfeed_115 0 1 decap_w0
xfeed_116 0 1 decap_w0
xfeed_117 0 1 decap_w0
xfeed_118 0 1 decap_w0
xfeed_119 0 1 decap_w0
xfeed_12659 0 1 decap_w0
xfeed_12658 0 1 decap_w0
xfeed_12657 0 1 decap_w0
xfeed_12656 0 1 decap_w0
xfeed_12655 0 1 decap_w0
xfeed_6459 0 1 decap_w0
xfeed_6458 0 1 tie
xfeed_6457 0 1 decap_w0
xfeed_6456 0 1 decap_w0
xfeed_6455 0 1 decap_w0
xfeed_6454 0 1 decap_w0
xfeed_6453 0 1 decap_w0
xfeed_6451 0 1 decap_w0
xfeed_6450 0 1 decap_w0
xfeed_5929 0 1 decap_w0
xfeed_5928 0 1 decap_w0
xfeed_5927 0 1 decap_w0
xfeed_5926 0 1 decap_w0
xfeed_5925 0 1 decap_w0
xfeed_5924 0 1 decap_w0
xfeed_5923 0 1 decap_w0
xfeed_5922 0 1 decap_w0
xfeed_5921 0 1 decap_w0
xfeed_5920 0 1 decap_w0
xfeed_2149 0 1 tie
xfeed_2148 0 1 decap_w0
xfeed_2147 0 1 decap_w0
xfeed_2146 0 1 decap_w0
xfeed_2145 0 1 decap_w0
xfeed_2144 0 1 decap_w0
xfeed_2143 0 1 decap_w0
xfeed_2142 0 1 tie
xfeed_2141 0 1 decap_w0
xfeed_2140 0 1 decap_w0
xfeed_1619 0 1 decap_w0
xfeed_1618 0 1 decap_w0
xfeed_1617 0 1 decap_w0
xfeed_1616 0 1 decap_w0
xfeed_1615 0 1 decap_w0
xfeed_1614 0 1 decap_w0
xfeed_1613 0 1 decap_w0
xfeed_1612 0 1 decap_w0
xfeed_1611 0 1 tie
xfeed_1610 0 1 decap_w0
xsubckt_551_nor2_x0 0 1 203 570 204 nor2_x0
xsubckt_1866_dff_x1 0 1 1958 1873 67 dff_x1
xsubckt_1868_dff_x1 0 1 1957 1871 67 dff_x1
xfeed_13199 0 1 decap_w0
xfeed_13198 0 1 decap_w0
xfeed_13197 0 1 decap_w0
xfeed_13196 0 1 decap_w0
xfeed_13195 0 1 decap_w0
xfeed_13194 0 1 decap_w0
xfeed_13193 0 1 decap_w0
xfeed_13192 0 1 decap_w0
xfeed_13191 0 1 decap_w0
xfeed_13190 0 1 decap_w0
xfeed_12661 0 1 decap_w0
xfeed_12660 0 1 decap_w0
xsubckt_862_nand3_x0 0 1 1619 184 177 1620 nand3_x0
xsubckt_345_nand2_x0 0 1 403 568 405 nand2_x0
xsubckt_405_nexor2_x0 0 1 344 1954 346 nexor2_x0
xsubckt_1582_or21nand_x0 0 1 1012 1105 1019 1017 or21nand_x0
xfeed_120 0 1 decap_w0
xfeed_121 0 1 decap_w0
xfeed_122 0 1 decap_w0
xfeed_123 0 1 decap_w0
xfeed_124 0 1 decap_w0
xfeed_125 0 1 decap_w0
xfeed_126 0 1 decap_w0
xfeed_127 0 1 decap_w0
xfeed_128 0 1 decap_w0
xfeed_129 0 1 decap_w0
xfeed_12669 0 1 tie
xfeed_12668 0 1 decap_w0
xfeed_12667 0 1 decap_w0
xfeed_12666 0 1 decap_w0
xfeed_12665 0 1 decap_w0
xfeed_12664 0 1 decap_w0
xfeed_12663 0 1 decap_w0
xfeed_12662 0 1 decap_w0
xfeed_6469 0 1 tie
xfeed_6467 0 1 decap_w0
xfeed_6466 0 1 decap_w0
xfeed_6464 0 1 decap_w0
xfeed_6463 0 1 decap_w0
xfeed_6462 0 1 decap_w0
xfeed_6461 0 1 decap_w0
xfeed_6460 0 1 decap_w0
xfeed_5939 0 1 decap_w0
xfeed_5938 0 1 decap_w0
xfeed_5937 0 1 decap_w0
xfeed_5936 0 1 decap_w0
xfeed_5935 0 1 decap_w0
xfeed_5934 0 1 decap_w0
xfeed_5933 0 1 decap_w0
xfeed_5932 0 1 tie
xfeed_5931 0 1 decap_w0
xfeed_5930 0 1 decap_w0
xfeed_2159 0 1 decap_w0
xfeed_2158 0 1 decap_w0
xfeed_2157 0 1 decap_w0
xfeed_2156 0 1 tie
xfeed_2155 0 1 decap_w0
xfeed_2154 0 1 decap_w0
xfeed_2153 0 1 decap_w0
xfeed_2152 0 1 decap_w0
xfeed_2151 0 1 decap_w0
xfeed_2150 0 1 decap_w0
xfeed_1629 0 1 decap_w0
xfeed_1628 0 1 decap_w0
xfeed_1627 0 1 decap_w0
xfeed_1626 0 1 decap_w0
xfeed_1625 0 1 decap_w0
xfeed_1624 0 1 decap_w0
xfeed_1623 0 1 decap_w0
xfeed_1622 0 1 decap_w0
xfeed_1621 0 1 decap_w0
xfeed_1620 0 1 decap_w0
xsubckt_1181_or21nand_x0 0 1 1381 1382 1387 1394 or21nand_x0
xsubckt_1162_nor4_x0 0 1 1399 2049 2048 2047 2046 nor4_x0
xsubckt_1142_and21nor_x0 0 1 1416 439 1420 1417 and21nor_x0
xsubckt_205_and2_x1 0 1 549 553 550 and2_x1
xsubckt_500_and4_x1 0 1 251 1916 771 679 571 and4_x1
xsubckt_1376_nand2_x0 0 1 1214 2051 479 nand2_x0
xfeed_130 0 1 decap_w0
xfeed_131 0 1 decap_w0
xfeed_132 0 1 decap_w0
xfeed_133 0 1 decap_w0
xfeed_134 0 1 decap_w0
xfeed_135 0 1 decap_w0
xfeed_136 0 1 decap_w0
xfeed_137 0 1 decap_w0
xfeed_138 0 1 decap_w0
xfeed_139 0 1 decap_w0
xfeed_12679 0 1 decap_w0
xfeed_12678 0 1 decap_w0
xfeed_12677 0 1 decap_w0
xfeed_12676 0 1 decap_w0
xfeed_12675 0 1 tie
xfeed_12674 0 1 decap_w0
xfeed_12673 0 1 decap_w0
xfeed_12672 0 1 decap_w0
xfeed_12671 0 1 decap_w0
xfeed_12670 0 1 decap_w0
xfeed_6479 0 1 tie
xfeed_6478 0 1 decap_w0
xfeed_6477 0 1 decap_w0
xfeed_6476 0 1 decap_w0
xfeed_6475 0 1 decap_w0
xfeed_6474 0 1 decap_w0
xfeed_6473 0 1 decap_w0
xfeed_6472 0 1 decap_w0
xfeed_6471 0 1 decap_w0
xfeed_6470 0 1 decap_w0
xfeed_5946 0 1 decap_w0
xfeed_5945 0 1 decap_w0
xfeed_5944 0 1 decap_w0
xfeed_5943 0 1 decap_w0
xfeed_5942 0 1 decap_w0
xfeed_5941 0 1 decap_w0
xfeed_5940 0 1 decap_w0
xfeed_2169 0 1 decap_w0
xfeed_2168 0 1 decap_w0
xfeed_2167 0 1 decap_w0
xfeed_2166 0 1 decap_w0
xfeed_2165 0 1 decap_w0
xfeed_2164 0 1 decap_w0
xfeed_2163 0 1 tie
xfeed_2162 0 1 decap_w0
xfeed_2161 0 1 decap_w0
xfeed_2160 0 1 decap_w0
xfeed_1639 0 1 decap_w0
xfeed_1638 0 1 decap_w0
xfeed_1637 0 1 decap_w0
xfeed_1636 0 1 decap_w0
xfeed_1635 0 1 decap_w0
xfeed_1634 0 1 decap_w0
xfeed_1633 0 1 decap_w0
xfeed_1632 0 1 decap_w0
xfeed_1631 0 1 decap_w0
xfeed_1630 0 1 decap_w0
xsubckt_720_or21nand_x0 0 1 1744 467 580 606 or21nand_x0
xsubckt_324_nand3_x0 0 1 424 682 595 557 nand3_x0
xsubckt_414_nand3_x0 0 1 335 616 558 460 nand3_x0
xsubckt_1281_or21nand_x0 0 1 1813 1309 1302 1301 or21nand_x0
xsubckt_1715_nand3_x0 0 1 879 888 884 882 nand3_x0
xfeed_5949 0 1 decap_w0
xfeed_5948 0 1 decap_w0
xfeed_5947 0 1 decap_w0
xsubckt_1018_nand2_x0 0 1 1513 1516 1514 nand2_x0
xsubckt_498_nand4_x0 0 1 253 653 649 645 535 nand4_x0
xsubckt_573_and21nor_x0 0 1 182 183 190 1948 and21nor_x0
xfeed_140 0 1 decap_w0
xfeed_141 0 1 decap_w0
xfeed_142 0 1 decap_w0
xfeed_143 0 1 decap_w0
xfeed_144 0 1 decap_w0
xfeed_145 0 1 decap_w0
xfeed_146 0 1 decap_w0
xfeed_147 0 1 decap_w0
xfeed_148 0 1 decap_w0
xfeed_149 0 1 decap_w0
xfeed_12689 0 1 decap_w0
xfeed_12688 0 1 decap_w0
xfeed_12687 0 1 decap_w0
xfeed_12686 0 1 tie
xfeed_12685 0 1 decap_w0
xfeed_12684 0 1 decap_w0
xfeed_12683 0 1 decap_w0
xfeed_12682 0 1 decap_w0
xfeed_12681 0 1 decap_w0
xfeed_12680 0 1 decap_w0
xfeed_6489 0 1 decap_w0
xfeed_6488 0 1 decap_w0
xfeed_6487 0 1 tie
xfeed_6486 0 1 decap_w0
xfeed_6485 0 1 decap_w0
xfeed_6484 0 1 decap_w0
xfeed_6483 0 1 tie
xfeed_6482 0 1 decap_w0
xfeed_6481 0 1 decap_w0
xfeed_6480 0 1 decap_w0
xfeed_5953 0 1 decap_w0
xfeed_5952 0 1 decap_w0
xfeed_5951 0 1 decap_w0
xfeed_5950 0 1 decap_w0
xfeed_2179 0 1 decap_w0
xfeed_2178 0 1 decap_w0
xfeed_2177 0 1 tie
xfeed_2176 0 1 decap_w0
xfeed_2175 0 1 decap_w0
xfeed_2174 0 1 decap_w0
xfeed_2173 0 1 decap_w0
xfeed_2172 0 1 decap_w0
xfeed_2171 0 1 decap_w0
xfeed_2170 0 1 tie
xfeed_1649 0 1 decap_w0
xfeed_1648 0 1 decap_w0
xfeed_1647 0 1 tie
xfeed_1646 0 1 decap_w0
xfeed_1645 0 1 decap_w0
xfeed_1644 0 1 decap_w0
xfeed_1643 0 1 decap_w0
xfeed_1642 0 1 decap_w0
xfeed_1641 0 1 decap_w0
xfeed_1640 0 1 decap_w0
xsubckt_1082_mux2_x1 0 1 1850 1463 1951 1576 mux2_x1
xsubckt_953_and3_x1 0 1 1567 660 654 527 and3_x1
xsubckt_1743_and21nor_x0 0 1 851 1142 1137 1126 and21nor_x0
xfeed_13309 0 1 tie
xfeed_13308 0 1 decap_w0
xfeed_13307 0 1 decap_w0
xfeed_13306 0 1 decap_w0
xfeed_13305 0 1 decap_w0
xfeed_13304 0 1 decap_w0
xfeed_13303 0 1 decap_w0
xfeed_13302 0 1 decap_w0
xfeed_13301 0 1 decap_w0
xfeed_13300 0 1 decap_w0
xfeed_5959 0 1 decap_w0
xfeed_5958 0 1 decap_w0
xfeed_5957 0 1 decap_w0
xfeed_5956 0 1 decap_w0
xfeed_5955 0 1 decap_w0
xfeed_5954 0 1 decap_w0
xsubckt_1001_nand2_x0 0 1 1528 1563 1529 nand2_x0
xsubckt_1539_and21nor_x0 0 1 1055 1056 1117 2047 and21nor_x0
xsubckt_1800_nexor2_x0 0 1 794 804 803 nexor2_x0
xfeed_150 0 1 decap_w0
xfeed_151 0 1 decap_w0
xfeed_152 0 1 decap_w0
xfeed_153 0 1 decap_w0
xfeed_154 0 1 decap_w0
xfeed_155 0 1 decap_w0
xfeed_156 0 1 decap_w0
xfeed_157 0 1 decap_w0
xfeed_158 0 1 decap_w0
xfeed_159 0 1 decap_w0
xfeed_12699 0 1 decap_w0
xfeed_12698 0 1 decap_w0
xfeed_12697 0 1 decap_w0
xfeed_12696 0 1 decap_w0
xfeed_12695 0 1 decap_w0
xfeed_12694 0 1 decap_w0
xfeed_12693 0 1 decap_w0
xfeed_12692 0 1 decap_w0
xfeed_12691 0 1 decap_w0
xfeed_12690 0 1 decap_w0
xfeed_7109 0 1 decap_w0
xfeed_7108 0 1 decap_w0
xfeed_7107 0 1 tie
xfeed_7106 0 1 decap_w0
xfeed_7105 0 1 decap_w0
xfeed_7104 0 1 decap_w0
xfeed_7103 0 1 decap_w0
xfeed_7102 0 1 decap_w0
xfeed_7101 0 1 decap_w0
xfeed_7100 0 1 decap_w0
xfeed_6499 0 1 decap_w0
xfeed_6498 0 1 decap_w0
xfeed_6497 0 1 decap_w0
xfeed_6496 0 1 decap_w0
xfeed_6495 0 1 decap_w0
xfeed_6494 0 1 tie
xfeed_6493 0 1 decap_w0
xfeed_6492 0 1 decap_w0
xfeed_6491 0 1 decap_w0
xfeed_6490 0 1 decap_w0
xfeed_5960 0 1 decap_w0
xfeed_2189 0 1 decap_w0
xfeed_2188 0 1 decap_w0
xfeed_2187 0 1 decap_w0
xfeed_2186 0 1 decap_w0
xfeed_2185 0 1 decap_w0
xfeed_2184 0 1 tie
xfeed_2183 0 1 decap_w0
xfeed_2182 0 1 decap_w0
xfeed_2181 0 1 decap_w0
xfeed_2180 0 1 decap_w0
xfeed_1659 0 1 decap_w0
xfeed_1658 0 1 decap_w0
xfeed_1657 0 1 decap_w0
xfeed_1656 0 1 decap_w0
xfeed_1655 0 1 decap_w0
xfeed_1654 0 1 decap_w0
xfeed_1653 0 1 decap_w0
xfeed_1652 0 1 decap_w0
xfeed_1651 0 1 decap_w0
xfeed_1650 0 1 decap_w0
xsubckt_975_and2_x1 0 1 1551 382 1552 and2_x1
xfeed_13319 0 1 decap_w0
xfeed_13318 0 1 decap_w0
xfeed_13317 0 1 decap_w0
xfeed_13316 0 1 decap_w0
xfeed_13315 0 1 decap_w0
xfeed_13314 0 1 tie
xfeed_13313 0 1 decap_w0
xfeed_13312 0 1 decap_w0
xfeed_13311 0 1 decap_w0
xfeed_13310 0 1 decap_w0
xfeed_5969 0 1 decap_w0
xfeed_5968 0 1 decap_w0
xfeed_5967 0 1 decap_w0
xfeed_5966 0 1 decap_w0
xfeed_5965 0 1 decap_w0
xfeed_5964 0 1 decap_w0
xfeed_5963 0 1 decap_w0
xfeed_5962 0 1 decap_w0
xfeed_5961 0 1 decap_w0
xsubckt_1744_and2_x1 0 1 850 852 851 and2_x1
xfeed_160 0 1 decap_w0
xfeed_161 0 1 decap_w0
xfeed_162 0 1 decap_w0
xfeed_163 0 1 decap_w0
xfeed_164 0 1 decap_w0
xfeed_165 0 1 decap_w0
xfeed_166 0 1 decap_w0
xfeed_167 0 1 decap_w0
xfeed_168 0 1 decap_w0
xfeed_169 0 1 decap_w0
xfeed_7119 0 1 tie
xfeed_7118 0 1 decap_w0
xfeed_7117 0 1 decap_w0
xfeed_7116 0 1 decap_w0
xfeed_7115 0 1 decap_w0
xfeed_7114 0 1 decap_w0
xfeed_7113 0 1 decap_w0
xfeed_7112 0 1 decap_w0
xfeed_7111 0 1 decap_w0
xfeed_7110 0 1 decap_w0
xfeed_2199 0 1 decap_w0
xfeed_2198 0 1 decap_w0
xfeed_2197 0 1 decap_w0
xfeed_2196 0 1 decap_w0
xfeed_2195 0 1 tie
xfeed_2194 0 1 decap_w0
xfeed_2193 0 1 decap_w0
xfeed_2192 0 1 decap_w0
xfeed_2191 0 1 tie
xfeed_2190 0 1 decap_w0
xfeed_1667 0 1 decap_w0
xfeed_1666 0 1 decap_w0
xfeed_1665 0 1 decap_w0
xfeed_1664 0 1 decap_w0
xfeed_1663 0 1 decap_w0
xfeed_1662 0 1 decap_w0
xfeed_1660 0 1 decap_w0
xsubckt_1217_and2_x1 0 1 1347 605 1348 and2_x1
xsubckt_931_mux2_x1 0 1 1886 2026 1600 1578 mux2_x1
xsubckt_360_and2_x1 0 1 388 510 389 and2_x1
xsubckt_1438_nand2_x0 0 1 1156 1158 1157 nand2_x0
xsubckt_1778_or21nand_x0 0 1 816 970 821 818 or21nand_x0
xfeed_13329 0 1 decap_w0
xfeed_13328 0 1 decap_w0
xfeed_13327 0 1 decap_w0
xfeed_13326 0 1 tie
xfeed_13325 0 1 decap_w0
xfeed_13324 0 1 decap_w0
xfeed_13323 0 1 decap_w0
xfeed_13322 0 1 decap_w0
xfeed_13321 0 1 decap_w0
xfeed_13320 0 1 decap_w0
xfeed_5979 0 1 decap_w0
xfeed_5978 0 1 tie
xfeed_5977 0 1 decap_w0
xfeed_5976 0 1 decap_w0
xfeed_5975 0 1 decap_w0
xfeed_5974 0 1 decap_w0
xfeed_5973 0 1 decap_w0
xfeed_5972 0 1 decap_w0
xfeed_5971 0 1 tie
xfeed_5970 0 1 decap_w0
xfeed_1669 0 1 decap_w0
xfeed_1668 0 1 decap_w0
xsubckt_422_or2_x1 0 1 327 554 456 or2_x1
xsubckt_1681_or21nand_x0 0 1 913 1067 924 1072 or21nand_x0
xfeed_170 0 1 decap_w0
xfeed_171 0 1 decap_w0
xfeed_172 0 1 decap_w0
xfeed_173 0 1 decap_w0
xfeed_174 0 1 decap_w0
xfeed_175 0 1 decap_w0
xfeed_176 0 1 decap_w0
xfeed_177 0 1 decap_w0
xfeed_178 0 1 decap_w0
xfeed_179 0 1 decap_w0
xfeed_7129 0 1 decap_w0
xfeed_7128 0 1 decap_w0
xfeed_7127 0 1 decap_w0
xfeed_7126 0 1 decap_w0
xfeed_7125 0 1 decap_w0
xfeed_7124 0 1 decap_w0
xfeed_7123 0 1 decap_w0
xfeed_7122 0 1 decap_w0
xfeed_7121 0 1 decap_w0
xfeed_7120 0 1 decap_w0
xfeed_1674 0 1 decap_w0
xfeed_1673 0 1 decap_w0
xfeed_1672 0 1 tie
xfeed_1671 0 1 decap_w0
xfeed_1670 0 1 decap_w0
xsubckt_1280_or21nand_x0 0 1 1301 1916 1311 1303 or21nand_x0
xsubckt_765_and3_x1 0 1 1704 1971 1749 1739 and3_x1
xsubckt_120_nand2_x0 0 1 648 1986 1992 nand2_x0
xsubckt_356_and2_x1 0 1 392 394 393 and2_x1
xsubckt_384_nand3_x0 0 1 365 608 603 557 nand3_x0
xsubckt_1312_or2_x1 0 1 1272 775 1273 or2_x1
xsubckt_1642_and21nor_x0 0 1 952 1102 955 954 and21nor_x0
xfeed_13339 0 1 decap_w0
xfeed_13338 0 1 decap_w0
xfeed_13337 0 1 decap_w0
xfeed_13336 0 1 decap_w0
xfeed_13335 0 1 decap_w0
xfeed_13334 0 1 decap_w0
xfeed_13333 0 1 decap_w0
xfeed_13332 0 1 decap_w0
xfeed_13331 0 1 decap_w0
xfeed_13330 0 1 decap_w0
xfeed_12801 0 1 decap_w0
xfeed_12800 0 1 tie
xfeed_5989 0 1 decap_w0
xfeed_5988 0 1 decap_w0
xfeed_5987 0 1 decap_w0
xfeed_5986 0 1 decap_w0
xfeed_5985 0 1 tie
xfeed_5984 0 1 decap_w0
xfeed_5983 0 1 decap_w0
xfeed_5982 0 1 decap_w0
xfeed_5981 0 1 decap_w0
xfeed_5980 0 1 decap_w0
xfeed_1679 0 1 decap_w0
xfeed_1678 0 1 decap_w0
xfeed_1677 0 1 decap_w0
xfeed_1676 0 1 decap_w0
xfeed_1675 0 1 decap_w0
xsubckt_1059_and4_x1 0 1 1483 653 623 525 519 and4_x1
xsubckt_737_nand2_x0 0 1 1728 2002 1746 nand2_x0
xsubckt_713_and2_x1 0 1 1751 566 1752 and2_x1
xsubckt_1477_or21nand_x0 0 1 1119 1121 1777 1781 or21nand_x0
xsubckt_1595_nand3_x0 0 1 999 1070 1018 1016 nand3_x0
xfeed_180 0 1 decap_w0
xfeed_181 0 1 decap_w0
xfeed_182 0 1 decap_w0
xfeed_183 0 1 decap_w0
xfeed_184 0 1 decap_w0
xfeed_185 0 1 decap_w0
xfeed_186 0 1 decap_w0
xfeed_187 0 1 decap_w0
xfeed_188 0 1 decap_w0
xfeed_189 0 1 decap_w0
xfeed_12809 0 1 tie
xfeed_12808 0 1 decap_w0
xfeed_12807 0 1 decap_w0
xfeed_12806 0 1 decap_w0
xfeed_12805 0 1 decap_w0
xfeed_12804 0 1 decap_w0
xfeed_12803 0 1 decap_w0
xfeed_12802 0 1 decap_w0
xfeed_7139 0 1 decap_w0
xfeed_7138 0 1 decap_w0
xfeed_7137 0 1 tie
xfeed_7136 0 1 decap_w0
xfeed_7135 0 1 decap_w0
xfeed_7134 0 1 decap_w0
xfeed_7133 0 1 decap_w0
xfeed_7132 0 1 decap_w0
xfeed_7131 0 1 decap_w0
xfeed_7130 0 1 decap_w0
xfeed_6609 0 1 decap_w0
xfeed_6608 0 1 decap_w0
xfeed_6607 0 1 tie
xfeed_6606 0 1 decap_w0
xfeed_6605 0 1 decap_w0
xfeed_6604 0 1 decap_w0
xfeed_6603 0 1 decap_w0
xfeed_6602 0 1 decap_w0
xfeed_6601 0 1 decap_w0
xfeed_6600 0 1 decap_w0
xfeed_1681 0 1 decap_w0
xfeed_1680 0 1 decap_w0
xsubckt_1007_and3_x1 0 1 1522 643 533 1523 and3_x1
xsubckt_709_and2_x1 0 1 1755 1757 1756 and2_x1
xfeed_13347 0 1 decap_w0
xfeed_13346 0 1 decap_w0
xfeed_13345 0 1 decap_w0
xfeed_13344 0 1 decap_w0
xfeed_13343 0 1 decap_w0
xfeed_13342 0 1 decap_w0
xfeed_13341 0 1 decap_w0
xfeed_13340 0 1 tie
xfeed_5999 0 1 decap_w0
xfeed_5998 0 1 decap_w0
xfeed_5997 0 1 decap_w0
xfeed_5996 0 1 decap_w0
xfeed_5995 0 1 decap_w0
xfeed_5994 0 1 decap_w0
xfeed_5993 0 1 decap_w0
xfeed_5992 0 1 decap_w0
xfeed_5991 0 1 decap_w0
xfeed_5990 0 1 tie
xfeed_1689 0 1 decap_w0
xfeed_1688 0 1 decap_w0
xfeed_1687 0 1 decap_w0
xfeed_1686 0 1 decap_w0
xfeed_1685 0 1 decap_w0
xfeed_1684 0 1 decap_w0
xfeed_1683 0 1 decap_w0
xfeed_1682 0 1 tie
xsubckt_1678_mux2_x1 0 1 916 963 918 1142 mux2_x1
xfeed_190 0 1 decap_w0
xfeed_191 0 1 decap_w0
xfeed_192 0 1 decap_w0
xfeed_193 0 1 decap_w0
xfeed_194 0 1 decap_w0
xfeed_195 0 1 decap_w0
xfeed_196 0 1 decap_w0
xfeed_197 0 1 decap_w0
xfeed_198 0 1 decap_w0
xfeed_199 0 1 decap_w0
xfeed_13349 0 1 decap_w0
xfeed_13348 0 1 decap_w0
xfeed_12819 0 1 decap_w0
xfeed_12818 0 1 decap_w0
xfeed_12817 0 1 decap_w0
xfeed_12816 0 1 decap_w0
xfeed_12815 0 1 decap_w0
xfeed_12814 0 1 decap_w0
xfeed_12813 0 1 decap_w0
xfeed_12812 0 1 decap_w0
xfeed_12811 0 1 decap_w0
xfeed_12810 0 1 decap_w0
xfeed_7149 0 1 tie
xfeed_7148 0 1 decap_w0
xfeed_7147 0 1 decap_w0
xfeed_7146 0 1 decap_w0
xfeed_7145 0 1 decap_w0
xfeed_7144 0 1 decap_w0
xfeed_7143 0 1 decap_w0
xfeed_7142 0 1 decap_w0
xfeed_7141 0 1 decap_w0
xfeed_7140 0 1 decap_w0
xfeed_6619 0 1 decap_w0
xfeed_6618 0 1 decap_w0
xfeed_6617 0 1 decap_w0
xfeed_6616 0 1 decap_w0
xfeed_6615 0 1 decap_w0
xfeed_6614 0 1 tie
xfeed_6613 0 1 decap_w0
xfeed_6612 0 1 decap_w0
xfeed_6611 0 1 decap_w0
xfeed_6610 0 1 decap_w0
xfeed_2309 0 1 decap_w0
xfeed_2308 0 1 decap_w0
xfeed_2307 0 1 decap_w0
xfeed_2306 0 1 decap_w0
xfeed_2305 0 1 decap_w0
xfeed_2304 0 1 decap_w0
xfeed_2303 0 1 decap_w0
xfeed_2302 0 1 decap_w0
xfeed_2301 0 1 decap_w0
xfeed_2300 0 1 decap_w0
xsubckt_1590_mux2_x1 0 1 1004 1053 1006 1142 mux2_x1
xfeed_13354 0 1 decap_w0
xfeed_13353 0 1 decap_w0
xfeed_13352 0 1 decap_w0
xfeed_13351 0 1 decap_w0
xfeed_13350 0 1 decap_w0
xfeed_1699 0 1 decap_w0
xfeed_1698 0 1 decap_w0
xfeed_1697 0 1 decap_w0
xfeed_1696 0 1 tie
xfeed_1695 0 1 decap_w0
xfeed_1694 0 1 decap_w0
xfeed_1693 0 1 decap_w0
xfeed_1692 0 1 decap_w0
xfeed_1691 0 1 decap_w0
xfeed_1690 0 1 decap_w0
xsubckt_986_and4_x1 0 1 1541 1550 1549 1547 1542 and4_x1
xsubckt_716_nand3_x0 0 1 1748 476 1759 1750 nand3_x0
xsubckt_626_nand3_x0 0 1 132 2018 184 177 nand3_x0
xfeed_13359 0 1 decap_w0
xfeed_13358 0 1 decap_w0
xfeed_13357 0 1 decap_w0
xfeed_13356 0 1 decap_w0
xfeed_13355 0 1 decap_w0
xfeed_12829 0 1 decap_w0
xfeed_12828 0 1 decap_w0
xfeed_12827 0 1 decap_w0
xfeed_12826 0 1 tie
xfeed_12825 0 1 decap_w0
xfeed_12824 0 1 decap_w0
xfeed_12823 0 1 decap_w0
xfeed_12822 0 1 decap_w0
xfeed_12821 0 1 decap_w0
xfeed_12820 0 1 decap_w0
xfeed_7159 0 1 decap_w0
xfeed_7158 0 1 tie
xfeed_7157 0 1 decap_w0
xfeed_7156 0 1 decap_w0
xfeed_7155 0 1 decap_w0
xfeed_7154 0 1 decap_w0
xfeed_7153 0 1 decap_w0
xfeed_7152 0 1 decap_w0
xfeed_7151 0 1 decap_w0
xfeed_7150 0 1 decap_w0
xfeed_6629 0 1 decap_w0
xfeed_6628 0 1 tie
xfeed_6627 0 1 decap_w0
xfeed_6626 0 1 decap_w0
xfeed_6625 0 1 decap_w0
xfeed_6624 0 1 decap_w0
xfeed_6623 0 1 decap_w0
xfeed_6622 0 1 decap_w0
xfeed_6621 0 1 tie
xfeed_6620 0 1 decap_w0
xfeed_2319 0 1 decap_w0
xfeed_2318 0 1 decap_w0
xfeed_2317 0 1 decap_w0
xfeed_2316 0 1 decap_w0
xfeed_2315 0 1 decap_w0
xfeed_2314 0 1 decap_w0
xfeed_2313 0 1 decap_w0
xfeed_2312 0 1 decap_w0
xfeed_2311 0 1 decap_w0
xfeed_2310 0 1 decap_w0
xsubckt_371_and21nor_x0 0 1 378 387 380 535 and21nor_x0
xsubckt_1638_and21nor_x0 0 1 956 1104 961 959 and21nor_x0
xcmpt_abc_11867_new_n425_hfns_0 0 1 687 685 buf_x4
xcmpt_abc_11867_new_n425_hfns_1 0 1 686 685 buf_x4
xcmpt_abc_11867_new_n425_hfns_2 0 1 685 688 buf_x4
xfeed_13361 0 1 decap_w0
xfeed_13360 0 1 decap_w0
xsubckt_485_and3_x1 0 1 265 270 269 266 and3_x1
xsubckt_1518_nor3_x0 0 1 1078 208 1080 1079 nor3_x0
xcmpt_abc_11867_new_n427_hfns_0 0 1 682 677 buf_x4
xcmpt_abc_11867_new_n427_hfns_1 0 1 681 677 buf_x4
xcmpt_abc_11867_new_n427_hfns_2 0 1 680 677 buf_x4
xcmpt_abc_11867_new_n427_hfns_3 0 1 679 677 buf_x4
xcmpt_abc_11867_new_n427_hfns_4 0 1 678 677 buf_x4
xcmpt_abc_11867_new_n427_hfns_5 0 1 677 683 buf_x4
xcmpt_abc_11867_new_n429_hfns_0 0 1 674 672 buf_x4
xcmpt_abc_11867_new_n429_hfns_1 0 1 673 672 buf_x4
xcmpt_abc_11867_new_n429_hfns_2 0 1 672 675 buf_x4
xfeed_13369 0 1 decap_w0
xfeed_13368 0 1 decap_w0
xfeed_13367 0 1 decap_w0
xfeed_13366 0 1 decap_w0
xfeed_13365 0 1 decap_w0
xfeed_13364 0 1 decap_w0
xfeed_13363 0 1 decap_w0
xfeed_13362 0 1 decap_w0
xfeed_12839 0 1 decap_w0
xfeed_12838 0 1 decap_w0
xfeed_12837 0 1 decap_w0
xfeed_12836 0 1 decap_w0
xfeed_12835 0 1 decap_w0
xfeed_12834 0 1 decap_w0
xfeed_12833 0 1 decap_w0
xfeed_12832 0 1 decap_w0
xfeed_12831 0 1 decap_w0
xfeed_12830 0 1 decap_w0
xfeed_7169 0 1 decap_w0
xfeed_7168 0 1 decap_w0
xfeed_7167 0 1 decap_w0
xfeed_7166 0 1 decap_w0
xfeed_7165 0 1 decap_w0
xfeed_7164 0 1 decap_w0
xfeed_7163 0 1 decap_w0
xfeed_7162 0 1 decap_w0
xfeed_7161 0 1 decap_w0
xfeed_7160 0 1 decap_w0
xfeed_6639 0 1 tie
xfeed_6638 0 1 decap_w0
xfeed_6637 0 1 decap_w0
xfeed_6636 0 1 decap_w0
xfeed_6635 0 1 tie
xfeed_6634 0 1 decap_w0
xfeed_6633 0 1 decap_w0
xfeed_6632 0 1 decap_w0
xfeed_6631 0 1 decap_w0
xfeed_6630 0 1 decap_w0
xfeed_2329 0 1 decap_w0
xfeed_2328 0 1 decap_w0
xfeed_2327 0 1 decap_w0
xfeed_2326 0 1 decap_w0
xfeed_2325 0 1 decap_w0
xfeed_2324 0 1 decap_w0
xfeed_2323 0 1 decap_w0
xfeed_2322 0 1 decap_w0
xfeed_2321 0 1 decap_w0
xfeed_2320 0 1 decap_w0
xsubckt_842_and3_x1 0 1 1636 2067 682 490 and3_x1
xsubckt_274_nexor2_x0 0 1 474 2055 1961 nexor2_x0
xsubckt_1303_nand2_x0 0 1 1281 775 1972 nand2_x0
xsubckt_1911_dff_x1 0 1 1995 1836 71 dff_x1
xsubckt_1913_dff_x1 0 1 1985 1834 61 dff_x1
xsubckt_797_nand2_x0 0 1 1675 1678 1676 nand2_x0
xsubckt_1780_or21nand_x0 0 1 814 1004 1003 1000 or21nand_x0
xsubckt_1799_and2_x1 0 1 795 801 796 and2_x1
xsubckt_1871_dff_x1 0 1 1960 1868 67 dff_x1
xsubckt_1915_dff_x1 0 1 2013 1832 67 dff_x1
xsubckt_1917_dff_x1 0 1 1961 1831 64 dff_x1
xsubckt_1919_dff_x1 0 1 2064 1829 45 dff_x1
xfeed_300 0 1 decap_w0
xfeed_301 0 1 decap_w0
xfeed_302 0 1 decap_w0
xfeed_303 0 1 decap_w0
xfeed_304 0 1 decap_w0
xfeed_305 0 1 decap_w0
xfeed_306 0 1 decap_w0
xfeed_307 0 1 decap_w0
xfeed_308 0 1 tie
xfeed_309 0 1 decap_w0
xfeed_13379 0 1 decap_w0
xfeed_13378 0 1 decap_w0
xfeed_13377 0 1 decap_w0
xfeed_13376 0 1 decap_w0
xfeed_13375 0 1 decap_w0
xfeed_13374 0 1 decap_w0
xfeed_13373 0 1 decap_w0
xfeed_13372 0 1 decap_w0
xfeed_13371 0 1 decap_w0
xfeed_13370 0 1 decap_w0
xfeed_12849 0 1 decap_w0
xfeed_12848 0 1 decap_w0
xfeed_12847 0 1 decap_w0
xfeed_12846 0 1 decap_w0
xfeed_12845 0 1 decap_w0
xfeed_12844 0 1 decap_w0
xfeed_12843 0 1 tie
xfeed_12842 0 1 decap_w0
xfeed_12841 0 1 decap_w0
xfeed_12840 0 1 decap_w0
xfeed_7179 0 1 decap_w0
xfeed_7178 0 1 tie
xfeed_7177 0 1 decap_w0
xfeed_7176 0 1 decap_w0
xfeed_7175 0 1 decap_w0
xfeed_7174 0 1 decap_w0
xfeed_7173 0 1 decap_w0
xfeed_7172 0 1 decap_w0
xfeed_7171 0 1 decap_w0
xfeed_7170 0 1 decap_w0
xfeed_6646 0 1 decap_w0
xfeed_6645 0 1 decap_w0
xfeed_6644 0 1 decap_w0
xfeed_6643 0 1 decap_w0
xfeed_6642 0 1 decap_w0
xfeed_6641 0 1 decap_w0
xfeed_6640 0 1 decap_w0
xfeed_2339 0 1 decap_w0
xfeed_2338 0 1 decap_w0
xfeed_2337 0 1 decap_w0
xfeed_2336 0 1 decap_w0
xfeed_2335 0 1 decap_w0
xfeed_2334 0 1 decap_w0
xfeed_2333 0 1 decap_w0
xfeed_2332 0 1 decap_w0
xfeed_2331 0 1 decap_w0
xfeed_2330 0 1 decap_w0
xfeed_1807 0 1 decap_w0
xfeed_1806 0 1 decap_w0
xfeed_1805 0 1 decap_w0
xfeed_1804 0 1 decap_w0
xfeed_1803 0 1 decap_w0
xfeed_1802 0 1 decap_w0
xfeed_1801 0 1 decap_w0
xfeed_1800 0 1 decap_w0
xsubckt_1110_and2_x1 0 1 1846 771 1439 and2_x1
xsubckt_912_mux2_x1 0 1 1903 1605 2043 1580 mux2_x1
xsubckt_750_and3_x1 0 1 1717 1973 1749 1739 and3_x1
xsubckt_389_and3_x1 0 1 360 660 651 646 and3_x1
xsubckt_529_nand2_x0 0 1 25 232 224 nand2_x0
xsubckt_1437_and21nor_x0 0 1 1157 775 1168 1160 and21nor_x0
xsubckt_1640_nand3_x0 0 1 954 1103 961 959 nand3_x0
xsubckt_1873_dff_x1 0 1 1944 1866 77 dff_x1
xsubckt_1875_dff_x1 0 1 1942 1864 77 dff_x1
xsubckt_1877_dff_x1 0 1 1933 1862 77 dff_x1
xfeed_6649 0 1 decap_w0
xfeed_6648 0 1 decap_w0
xfeed_6647 0 1 decap_w0
xfeed_1809 0 1 decap_w0
xfeed_1808 0 1 decap_w0
xsubckt_1232_mux2_x1 0 1 1829 2105 2064 1334 mux2_x1
xsubckt_1070_and3_x1 0 1 1473 652 526 1563 and3_x1
xsubckt_908_mux2_x1 0 1 1906 2014 1581 1619 mux2_x1
xsubckt_337_and2_x1 0 1 411 682 421 and2_x1
xsubckt_602_nand2_x0 0 1 154 2044 172 nand2_x0
xsubckt_1879_dff_x1 0 1 1964 1860 77 dff_x1
xfeed_310 0 1 decap_w0
xfeed_311 0 1 decap_w0
xfeed_312 0 1 decap_w0
xfeed_313 0 1 decap_w0
xfeed_314 0 1 decap_w0
xfeed_315 0 1 tie
xfeed_316 0 1 decap_w0
xfeed_317 0 1 decap_w0
xfeed_318 0 1 decap_w0
xfeed_319 0 1 decap_w0
xfeed_13389 0 1 tie
xfeed_13388 0 1 decap_w0
xfeed_13387 0 1 decap_w0
xfeed_13386 0 1 decap_w0
xfeed_13385 0 1 decap_w0
xfeed_13384 0 1 decap_w0
xfeed_13383 0 1 decap_w0
xfeed_13382 0 1 decap_w0
xfeed_13381 0 1 decap_w0
xfeed_13380 0 1 decap_w0
xfeed_12859 0 1 tie
xfeed_12858 0 1 decap_w0
xfeed_12857 0 1 decap_w0
xfeed_12856 0 1 decap_w0
xfeed_12855 0 1 decap_w0
xfeed_12854 0 1 decap_w0
xfeed_12853 0 1 decap_w0
xfeed_12852 0 1 decap_w0
xfeed_12851 0 1 decap_w0
xfeed_12850 0 1 decap_w0
xfeed_7189 0 1 decap_w0
xfeed_7188 0 1 decap_w0
xfeed_7187 0 1 decap_w0
xfeed_7186 0 1 decap_w0
xfeed_7185 0 1 decap_w0
xfeed_7184 0 1 decap_w0
xfeed_7183 0 1 decap_w0
xfeed_7182 0 1 decap_w0
xfeed_7181 0 1 decap_w0
xfeed_7180 0 1 decap_w0
xfeed_6653 0 1 decap_w0
xfeed_6652 0 1 decap_w0
xfeed_6651 0 1 decap_w0
xfeed_6650 0 1 decap_w0
xfeed_2349 0 1 decap_w0
xfeed_2348 0 1 decap_w0
xfeed_2347 0 1 decap_w0
xfeed_2346 0 1 decap_w0
xfeed_2345 0 1 decap_w0
xfeed_2344 0 1 decap_w0
xfeed_2343 0 1 decap_w0
xfeed_2342 0 1 decap_w0
xfeed_2341 0 1 decap_w0
xfeed_2340 0 1 decap_w0
xfeed_1814 0 1 decap_w0
xfeed_1813 0 1 decap_w0
xfeed_1812 0 1 decap_w0
xfeed_1811 0 1 decap_w0
xfeed_1810 0 1 decap_w0
xsubckt_297_and3_x1 0 1 451 1927 713 589 and3_x1
xsubckt_194_or2_x1 0 1 564 570 567 or2_x1
xsubckt_183_and4_x1 0 1 575 714 1928 681 674 and4_x1
xsubckt_1370_nand3_x0 0 1 1219 1245 1234 1222 nand3_x0
xsubckt_1546_nand4_x0 0 1 1048 1997 1128 1098 1097 nand4_x0
xsubckt_1791_nor2_x0 0 1 803 1141 875 nor2_x0
xsubckt_1793_nexor2_x0 0 1 801 807 802 nexor2_x0
xfeed_14009 0 1 tie
xfeed_14008 0 1 tie
xfeed_14007 0 1 tie
xfeed_14006 0 1 tie
xfeed_14005 0 1 tie
xfeed_14004 0 1 tie
xfeed_14003 0 1 tie
xfeed_14002 0 1 tie
xfeed_14001 0 1 tie
xfeed_14000 0 1 tie
xfeed_6659 0 1 decap_w0
xfeed_6658 0 1 tie
xfeed_6657 0 1 decap_w0
xfeed_6656 0 1 decap_w0
xfeed_6655 0 1 decap_w0
xfeed_6654 0 1 decap_w0
xfeed_1819 0 1 decap_w0
xfeed_1818 0 1 decap_w0
xfeed_1817 0 1 decap_w0
xfeed_1816 0 1 decap_w0
xfeed_1815 0 1 decap_w0
xsubckt_1140_mux2_x1 0 1 1418 758 2051 288 mux2_x1
xsubckt_1136_and21nor_x0 0 1 1422 288 1624 1435 and21nor_x0
xsubckt_894_mux2_x1 0 1 1908 2016 1593 1619 mux2_x1
xsubckt_467_and21nor_x0 0 1 283 548 421 608 and21nor_x0
xsubckt_1537_and2_x1 0 1 1057 1635 1058 and2_x1
xfeed_320 0 1 decap_w0
xfeed_321 0 1 decap_w0
xfeed_322 0 1 tie
xfeed_323 0 1 decap_w0
xfeed_324 0 1 decap_w0
xfeed_325 0 1 decap_w0
xfeed_326 0 1 decap_w0
xfeed_327 0 1 decap_w0
xfeed_328 0 1 decap_w0
xfeed_329 0 1 decap_w0
xfeed_13399 0 1 decap_w0
xfeed_13398 0 1 decap_w0
xfeed_13397 0 1 decap_w0
xfeed_13396 0 1 decap_w0
xfeed_13395 0 1 decap_w0
xfeed_13394 0 1 decap_w0
xfeed_13393 0 1 decap_w0
xfeed_13392 0 1 decap_w0
xfeed_13391 0 1 decap_w0
xfeed_13390 0 1 decap_w0
xfeed_12869 0 1 decap_w0
xfeed_12868 0 1 decap_w0
xfeed_12867 0 1 decap_w0
xfeed_12866 0 1 decap_w0
xfeed_12865 0 1 decap_w0
xfeed_12864 0 1 decap_w0
xfeed_12863 0 1 decap_w0
xfeed_12862 0 1 decap_w0
xfeed_12861 0 1 decap_w0
xfeed_12860 0 1 decap_w0
xfeed_7199 0 1 decap_w0
xfeed_7198 0 1 decap_w0
xfeed_7197 0 1 decap_w0
xfeed_7196 0 1 decap_w0
xfeed_7195 0 1 tie
xfeed_7194 0 1 decap_w0
xfeed_7193 0 1 decap_w0
xfeed_7192 0 1 tie
xfeed_7191 0 1 decap_w0
xfeed_7190 0 1 decap_w0
xfeed_6660 0 1 decap_w0
xfeed_2359 0 1 decap_w0
xfeed_2358 0 1 decap_w0
xfeed_2357 0 1 decap_w0
xfeed_2355 0 1 tie
xfeed_2354 0 1 decap_w0
xfeed_2353 0 1 decap_w0
xfeed_2352 0 1 decap_w0
xfeed_2351 0 1 decap_w0
xfeed_2350 0 1 decap_w0
xfeed_1821 0 1 decap_w0
xfeed_1820 0 1 decap_w0
xsubckt_1190_nand3_x0 0 1 1374 1378 1377 1376 nand3_x0
xsubckt_1775_nexor2_x0 0 1 819 976 972 nexor2_x0
xfeed_14019 0 1 tie
xfeed_14018 0 1 tie
xfeed_14017 0 1 tie
xfeed_14016 0 1 tie
xfeed_14015 0 1 tie
xfeed_14014 0 1 tie
xfeed_14013 0 1 tie
xfeed_14010 0 1 tie
xfeed_6669 0 1 decap_w0
xfeed_6668 0 1 decap_w0
xfeed_6667 0 1 decap_w0
xfeed_6666 0 1 decap_w0
xfeed_6665 0 1 tie
xfeed_6664 0 1 decap_w0
xfeed_6663 0 1 decap_w0
xfeed_6662 0 1 decap_w0
xfeed_6661 0 1 decap_w0
xfeed_1829 0 1 decap_w0
xfeed_1828 0 1 decap_w0
xfeed_1827 0 1 decap_w0
xfeed_1826 0 1 decap_w0
xfeed_1825 0 1 decap_w0
xfeed_1824 0 1 decap_w0
xfeed_1823 0 1 decap_w0
xfeed_1822 0 1 decap_w0
xsubckt_1383_and4_x1 0 1 1207 1245 1234 1222 1209 and4_x1
xsubckt_1766_nexor2_x0 0 1 828 844 841 nexor2_x0
xfeed_330 0 1 decap_w0
xfeed_331 0 1 tie
xfeed_332 0 1 decap_w0
xfeed_333 0 1 decap_w0
xfeed_334 0 1 decap_w0
xfeed_335 0 1 decap_w0
xfeed_336 0 1 decap_w0
xfeed_337 0 1 decap_w0
xfeed_338 0 1 decap_w0
xfeed_12879 0 1 decap_w0
xfeed_12878 0 1 decap_w0
xfeed_12877 0 1 decap_w0
xfeed_12876 0 1 tie
xfeed_12875 0 1 decap_w0
xfeed_12874 0 1 decap_w0
xfeed_12873 0 1 decap_w0
xfeed_12872 0 1 decap_w0
xfeed_12871 0 1 decap_w0
xfeed_12870 0 1 decap_w0
xfeed_2367 0 1 decap_w0
xfeed_2366 0 1 decap_w0
xfeed_2365 0 1 decap_w0
xfeed_2364 0 1 decap_w0
xfeed_2363 0 1 decap_w0
xfeed_2362 0 1 decap_w0
xfeed_2361 0 1 decap_w0
xfeed_2360 0 1 decap_w0
xsubckt_148_nand3_x0 0 1 620 627 623 621 nand3_x0
xfeed_14029 0 1 tie
xfeed_14028 0 1 tie
xfeed_14027 0 1 tie
xfeed_14026 0 1 tie
xfeed_14025 0 1 tie
xfeed_14024 0 1 tie
xfeed_14023 0 1 tie
xfeed_14022 0 1 tie
xfeed_14021 0 1 tie
xfeed_14020 0 1 tie
xfeed_6679 0 1 decap_w0
xfeed_6678 0 1 decap_w0
xfeed_6677 0 1 decap_w0
xfeed_6676 0 1 decap_w0
xfeed_6675 0 1 decap_w0
xfeed_6674 0 1 decap_w0
xfeed_6673 0 1 decap_w0
xfeed_6672 0 1 decap_w0
xfeed_6671 0 1 decap_w0
xfeed_6670 0 1 tie
xfeed_2369 0 1 decap_w0
xfeed_2368 0 1 tie
xfeed_1839 0 1 decap_w0
xfeed_1838 0 1 decap_w0
xfeed_1837 0 1 decap_w0
xfeed_1836 0 1 decap_w0
xfeed_1835 0 1 decap_w0
xfeed_1834 0 1 decap_w0
xfeed_1833 0 1 decap_w0
xfeed_1832 0 1 decap_w0
xfeed_1831 0 1 decap_w0
xfeed_1830 0 1 decap_w0
xsubckt_1044_mux2_x1 0 1 1856 1496 1947 1576 mux2_x1
xsubckt_94_mux2_x1 0 1 692 698 697 774 mux2_x1
xsubckt_575_nand4_x0 0 1 180 195 194 188 182 nand4_x0
xsubckt_1353_and2_x1 0 1 1235 1241 1236 and2_x1
xfeed_340 0 1 decap_w0
xfeed_341 0 1 decap_w0
xfeed_342 0 1 decap_w0
xfeed_343 0 1 decap_w0
xfeed_344 0 1 decap_w0
xfeed_345 0 1 decap_w0
xfeed_346 0 1 decap_w0
xfeed_347 0 1 decap_w0
xfeed_348 0 1 decap_w0
xfeed_349 0 1 decap_w0
xfeed_12889 0 1 decap_w0
xfeed_12888 0 1 decap_w0
xfeed_12887 0 1 decap_w0
xfeed_12886 0 1 decap_w0
xfeed_12885 0 1 decap_w0
xfeed_12884 0 1 decap_w0
xfeed_12883 0 1 decap_w0
xfeed_12882 0 1 tie
xfeed_12881 0 1 decap_w0
xfeed_12880 0 1 decap_w0
xfeed_2374 0 1 decap_w0
xfeed_2373 0 1 decap_w0
xfeed_2372 0 1 decap_w0
xfeed_2371 0 1 decap_w0
xfeed_2370 0 1 decap_w0
xfeed_14039 0 1 tie
xfeed_14038 0 1 tie
xfeed_14037 0 1 tie
xfeed_14036 0 1 tie
xfeed_14035 0 1 tie
xfeed_14034 0 1 tie
xfeed_14032 0 1 tie
xfeed_14031 0 1 tie
xfeed_13501 0 1 decap_w0
xfeed_13500 0 1 decap_w0
xfeed_6689 0 1 decap_w0
xfeed_6688 0 1 decap_w0
xfeed_6687 0 1 decap_w0
xfeed_6686 0 1 decap_w0
xfeed_6685 0 1 decap_w0
xfeed_6684 0 1 decap_w0
xfeed_6683 0 1 decap_w0
xfeed_6682 0 1 decap_w0
xfeed_6681 0 1 decap_w0
xfeed_6680 0 1 decap_w0
xfeed_2379 0 1 decap_w0
xfeed_2378 0 1 decap_w0
xfeed_2377 0 1 decap_w0
xfeed_2376 0 1 decap_w0
xfeed_2375 0 1 decap_w0
xfeed_1849 0 1 decap_w0
xfeed_1848 0 1 decap_w0
xfeed_1847 0 1 decap_w0
xfeed_1846 0 1 decap_w0
xfeed_1845 0 1 decap_w0
xfeed_1844 0 1 decap_w0
xfeed_1843 0 1 decap_w0
xfeed_1842 0 1 decap_w0
xfeed_1841 0 1 decap_w0
xfeed_1840 0 1 decap_w0
xfeed_359 0 1 decap_w0
xfeed_358 0 1 decap_w0
xfeed_357 0 1 decap_w0
xfeed_356 0 1 decap_w0
xsubckt_1261_and2_x1 0 1 1319 435 1320 and2_x1
xsubckt_823_and3_x1 0 1 1653 1978 1749 1739 and3_x1
xsubckt_344_or4_x1 0 1 404 1929 1923 1927 1928 or4_x1
xsubckt_1696_nand4_x0 0 1 898 2002 1128 1098 1097 nand4_x0
xfeed_350 0 1 decap_w0
xfeed_351 0 1 decap_w0
xfeed_352 0 1 decap_w0
xfeed_353 0 1 decap_w0
xfeed_354 0 1 decap_w0
xfeed_355 0 1 decap_w0
xfeed_13509 0 1 decap_w0
xfeed_13508 0 1 decap_w0
xfeed_13507 0 1 decap_w0
xfeed_13506 0 1 decap_w0
xfeed_13505 0 1 decap_w0
xfeed_13504 0 1 decap_w0
xfeed_13503 0 1 decap_w0
xfeed_13502 0 1 decap_w0
xfeed_12899 0 1 tie
xfeed_12898 0 1 decap_w0
xfeed_12897 0 1 decap_w0
xfeed_12896 0 1 decap_w0
xfeed_12895 0 1 decap_w0
xfeed_12894 0 1 decap_w0
xfeed_12893 0 1 decap_w0
xfeed_12892 0 1 decap_w0
xfeed_12891 0 1 decap_w0
xfeed_12890 0 1 tie
xfeed_7309 0 1 decap_w0
xfeed_7308 0 1 decap_w0
xfeed_7307 0 1 decap_w0
xfeed_7306 0 1 decap_w0
xfeed_7305 0 1 decap_w0
xfeed_7304 0 1 tie
xfeed_7303 0 1 decap_w0
xfeed_7302 0 1 decap_w0
xfeed_7301 0 1 decap_w0
xfeed_7300 0 1 decap_w0
xfeed_2381 0 1 tie
xfeed_2380 0 1 decap_w0
xsubckt_260_and4_x1 0 1 491 1929 715 714 1928 and4_x1
xfeed_14047 0 1 tie
xfeed_14046 0 1 tie
xfeed_14045 0 1 tie
xfeed_14043 0 1 tie
xfeed_14041 0 1 tie
xfeed_14040 0 1 tie
xfeed_6699 0 1 decap_w0
xfeed_6698 0 1 decap_w0
xfeed_6697 0 1 decap_w0
xfeed_6696 0 1 decap_w0
xfeed_6695 0 1 decap_w0
xfeed_6694 0 1 decap_w0
xfeed_6693 0 1 decap_w0
xfeed_6692 0 1 decap_w0
xfeed_6691 0 1 decap_w0
xfeed_6690 0 1 decap_w0
xfeed_2389 0 1 decap_w0
xfeed_2388 0 1 tie
xfeed_2386 0 1 decap_w0
xfeed_2385 0 1 decap_w0
xfeed_2384 0 1 decap_w0
xfeed_2383 0 1 decap_w0
xfeed_2382 0 1 decap_w0
xfeed_1859 0 1 decap_w0
xfeed_1858 0 1 decap_w0
xfeed_1857 0 1 decap_w0
xfeed_1856 0 1 decap_w0
xfeed_1855 0 1 decap_w0
xfeed_1854 0 1 decap_w0
xfeed_1853 0 1 decap_w0
xfeed_1852 0 1 decap_w0
xfeed_1851 0 1 tie
xfeed_1850 0 1 decap_w0
xfeed_369 0 1 decap_w0
xfeed_368 0 1 decap_w0
xfeed_367 0 1 decap_w0
xfeed_366 0 1 decap_w0
xfeed_365 0 1 decap_w0
xfeed_364 0 1 decap_w0
xfeed_363 0 1 decap_w0
xfeed_362 0 1 decap_w0
xfeed_360 0 1 decap_w0
xsubckt_822_or2_x1 0 1 2103 1660 1654 or2_x1
xsubckt_433_or2_x1 0 1 317 684 462 or2_x1
xfeed_14049 0 1 tie
xfeed_14048 0 1 tie
xfeed_13519 0 1 decap_w0
xfeed_13518 0 1 decap_w0
xfeed_13517 0 1 decap_w0
xfeed_13516 0 1 decap_w0
xfeed_13515 0 1 decap_w0
xfeed_13514 0 1 decap_w0
xfeed_13513 0 1 decap_w0
xfeed_13512 0 1 decap_w0
xfeed_13511 0 1 decap_w0
xfeed_13510 0 1 decap_w0
xfeed_7319 0 1 decap_w0
xfeed_7318 0 1 tie
xfeed_7317 0 1 decap_w0
xfeed_7316 0 1 decap_w0
xfeed_7315 0 1 decap_w0
xfeed_7314 0 1 decap_w0
xfeed_7313 0 1 decap_w0
xfeed_7312 0 1 decap_w0
xfeed_7311 0 1 decap_w0
xfeed_3009 0 1 decap_w0
xfeed_3008 0 1 decap_w0
xfeed_3007 0 1 decap_w0
xfeed_3006 0 1 decap_w0
xfeed_3005 0 1 decap_w0
xfeed_3004 0 1 decap_w0
xfeed_3003 0 1 tie
xfeed_3002 0 1 decap_w0
xfeed_3001 0 1 decap_w0
xfeed_3000 0 1 decap_w0
xsubckt_780_or2_x1 0 1 2094 1692 1691 or2_x1
xsubckt_175_or3_x1 0 1 583 1920 2055 1921 or3_x1
xsubckt_124_nand2_x0 0 1 644 660 646 nand2_x0
xsubckt_1501_nand4_x0 0 1 1095 1996 1128 1098 1097 nand4_x0
xfeed_14054 0 1 tie
xfeed_14053 0 1 tie
xfeed_14052 0 1 tie
xfeed_14051 0 1 tie
xfeed_14050 0 1 tie
xfeed_2399 0 1 decap_w0
xfeed_2398 0 1 decap_w0
xfeed_2397 0 1 decap_w0
xfeed_2396 0 1 decap_w0
xfeed_2395 0 1 decap_w0
xfeed_2393 0 1 decap_w0
xfeed_2392 0 1 decap_w0
xfeed_2391 0 1 decap_w0
xfeed_2390 0 1 decap_w0
xfeed_1869 0 1 decap_w0
xfeed_1868 0 1 decap_w0
xfeed_1867 0 1 decap_w0
xfeed_1866 0 1 decap_w0
xfeed_1865 0 1 decap_w0
xfeed_1864 0 1 decap_w0
xfeed_1863 0 1 decap_w0
xfeed_1862 0 1 decap_w0
xfeed_1861 0 1 decap_w0
xfeed_1860 0 1 decap_w0
xfeed_379 0 1 decap_w0
xfeed_378 0 1 decap_w0
xfeed_377 0 1 decap_w0
xfeed_376 0 1 decap_w0
xfeed_375 0 1 decap_w0
xfeed_374 0 1 decap_w0
xfeed_373 0 1 decap_w0
xfeed_372 0 1 decap_w0
xfeed_371 0 1 decap_w0
xfeed_370 0 1 decap_w0
xsubckt_1068_nand4_x0 0 1 1475 650 637 633 525 nand4_x0
xsubckt_1329_or2_x1 0 1 1257 1261 1258 or2_x1
xsubckt_1716_or2_x1 0 1 878 696 1116 or2_x1
xfeed_14056 0 1 tie
xfeed_14055 0 1 tie
xfeed_13529 0 1 decap_w0
xfeed_13528 0 1 decap_w0
xfeed_13527 0 1 decap_w0
xfeed_13526 0 1 decap_w0
xfeed_13525 0 1 decap_w0
xfeed_13524 0 1 decap_w0
xfeed_13523 0 1 decap_w0
xfeed_13522 0 1 decap_w0
xfeed_13521 0 1 decap_w0
xfeed_13520 0 1 decap_w0
xfeed_7329 0 1 decap_w0
xfeed_7328 0 1 decap_w0
xfeed_7327 0 1 decap_w0
xfeed_7326 0 1 decap_w0
xfeed_7325 0 1 decap_w0
xfeed_7324 0 1 decap_w0
xfeed_7323 0 1 decap_w0
xfeed_7322 0 1 decap_w0
xfeed_7321 0 1 decap_w0
xfeed_7320 0 1 decap_w0
xfeed_3019 0 1 decap_w0
xfeed_3018 0 1 decap_w0
xfeed_3017 0 1 decap_w0
xfeed_3016 0 1 decap_w0
xfeed_3015 0 1 tie
xfeed_3014 0 1 decap_w0
xfeed_3013 0 1 decap_w0
xfeed_3012 0 1 decap_w0
xfeed_3011 0 1 decap_w0
xfeed_3010 0 1 decap_w0
xsubckt_1073_and2_x1 0 1 1470 1576 1531 and2_x1
xsubckt_788_or2_x1 0 1 2093 1690 1684 or2_x1
xsubckt_1596_and2_x1 0 1 998 1001 999 and2_x1
xfeed_14061 0 1 tie
xfeed_1879 0 1 decap_w0
xfeed_1878 0 1 decap_w0
xfeed_1877 0 1 decap_w0
xfeed_1876 0 1 decap_w0
xfeed_1875 0 1 decap_w0
xfeed_1874 0 1 decap_w0
xfeed_1873 0 1 decap_w0
xfeed_1872 0 1 decap_w0
xfeed_1871 0 1 decap_w0
xfeed_1870 0 1 decap_w0
xfeed_389 0 1 decap_w0
xfeed_388 0 1 decap_w0
xfeed_387 0 1 decap_w0
xfeed_386 0 1 decap_w0
xfeed_385 0 1 decap_w0
xfeed_384 0 1 decap_w0
xfeed_383 0 1 decap_w0
xfeed_382 0 1 decap_w0
xfeed_381 0 1 decap_w0
xfeed_380 0 1 decap_w0
xsubckt_521_and4_x1 0 1 231 545 542 514 513 and4_x1
xsubckt_1289_or2_x1 0 1 1293 1299 1294 or2_x1
xsubckt_1335_and21nor_x0 0 1 1252 748 478 1317 and21nor_x0
xsubckt_1644_mux2_x1 0 1 950 956 951 964 mux2_x1
xfeed_14068 0 1 tie
xfeed_14067 0 1 tie
xfeed_14066 0 1 tie
xfeed_14065 0 1 tie
xfeed_14064 0 1 tie
xfeed_14063 0 1 tie
xfeed_14062 0 1 tie
xfeed_13539 0 1 decap_w0
xfeed_13538 0 1 decap_w0
xfeed_13537 0 1 decap_w0
xfeed_13536 0 1 decap_w0
xfeed_13535 0 1 decap_w0
xfeed_13534 0 1 decap_w0
xfeed_13533 0 1 decap_w0
xfeed_13532 0 1 decap_w0
xfeed_13531 0 1 decap_w0
xfeed_13530 0 1 decap_w0
xfeed_7339 0 1 decap_w0
xfeed_7338 0 1 decap_w0
xfeed_7337 0 1 decap_w0
xfeed_7336 0 1 decap_w0
xfeed_7335 0 1 decap_w0
xfeed_7334 0 1 decap_w0
xfeed_7333 0 1 tie
xfeed_7332 0 1 decap_w0
xfeed_7331 0 1 decap_w0
xfeed_7330 0 1 decap_w0
xfeed_6800 0 1 decap_w0
xfeed_3029 0 1 tie
xfeed_3028 0 1 decap_w0
xfeed_3027 0 1 decap_w0
xfeed_3026 0 1 decap_w0
xfeed_3025 0 1 decap_w0
xfeed_3024 0 1 decap_w0
xfeed_3023 0 1 decap_w0
xfeed_3022 0 1 tie
xfeed_3020 0 1 decap_w0
xsubckt_1117_mux2_x1 0 1 1840 1998 1989 1438 mux2_x1
xsubckt_900_nexor2_x0 0 1 1587 1595 1588 nexor2_x0
xsubckt_108_and3_x1 0 1 667 679 674 670 and3_x1
xsubckt_1364_and4_x1 0 1 1225 435 1670 1227 1226 and4_x1
xsubckt_1404_nand3_x0 0 1 1188 2069 666 657 nand3_x0
xsubckt_1478_and3_x1 0 1 1118 498 211 1763 and3_x1
xsubckt_1668_nand4_x0 0 1 926 2001 1128 1098 1097 nand4_x0
xfeed_6809 0 1 decap_w0
xfeed_6808 0 1 decap_w0
xfeed_6807 0 1 decap_w0
xfeed_6806 0 1 tie
xfeed_6805 0 1 decap_w0
xfeed_6804 0 1 decap_w0
xfeed_6803 0 1 decap_w0
xfeed_6802 0 1 decap_w0
xfeed_6801 0 1 decap_w0
xfeed_1889 0 1 decap_w0
xfeed_1888 0 1 decap_w0
xfeed_1887 0 1 decap_w0
xfeed_1886 0 1 tie
xfeed_1885 0 1 decap_w0
xfeed_1884 0 1 decap_w0
xfeed_1883 0 1 decap_w0
xfeed_1882 0 1 decap_w0
xfeed_1881 0 1 decap_w0
xfeed_1880 0 1 decap_w0
xfeed_399 0 1 decap_w0
xfeed_398 0 1 decap_w0
xfeed_397 0 1 decap_w0
xfeed_396 0 1 decap_w0
xfeed_395 0 1 decap_w0
xfeed_394 0 1 decap_w0
xfeed_393 0 1 decap_w0
xfeed_392 0 1 decap_w0
xfeed_391 0 1 decap_w0
xfeed_390 0 1 decap_w0
xsubckt_111_or21nand_x0 0 1 657 782 730 1995 or21nand_x0
xsubckt_1574_or21nand_x0 0 1 1020 1023 1122 100 or21nand_x0
xsubckt_1578_nand4_x0 0 1 1016 1998 1128 1098 1097 nand4_x0
xfeed_14079 0 1 tie
xfeed_14077 0 1 tie
xfeed_14076 0 1 tie
xfeed_14075 0 1 tie
xfeed_14074 0 1 tie
xfeed_14073 0 1 tie
xfeed_14072 0 1 tie
xfeed_14071 0 1 tie
xfeed_14070 0 1 tie
xfeed_13549 0 1 decap_w0
xfeed_13548 0 1 decap_w0
xfeed_13547 0 1 decap_w0
xfeed_13546 0 1 decap_w0
xfeed_13545 0 1 decap_w0
xfeed_13544 0 1 decap_w0
xfeed_13543 0 1 decap_w0
xfeed_13542 0 1 decap_w0
xfeed_13541 0 1 decap_w0
xfeed_13540 0 1 decap_w0
xfeed_7346 0 1 decap_w0
xfeed_7345 0 1 decap_w0
xfeed_7344 0 1 decap_w0
xfeed_7343 0 1 decap_w0
xfeed_7342 0 1 decap_w0
xfeed_7341 0 1 decap_w0
xfeed_7340 0 1 decap_w0
xfeed_3039 0 1 decap_w0
xfeed_3038 0 1 decap_w0
xfeed_3037 0 1 decap_w0
xfeed_3036 0 1 decap_w0
xfeed_3035 0 1 decap_w0
xfeed_3034 0 1 decap_w0
xfeed_3033 0 1 decap_w0
xfeed_3032 0 1 decap_w0
xfeed_3031 0 1 decap_w0
xfeed_3030 0 1 decap_w0
xfeed_2507 0 1 decap_w0
xfeed_2506 0 1 decap_w0
xfeed_2505 0 1 decap_w0
xfeed_2504 0 1 decap_w0
xfeed_2503 0 1 decap_w0
xfeed_2502 0 1 tie
xfeed_2501 0 1 decap_w0
xfeed_2500 0 1 decap_w0
xcmpt_abc_11867_new_n430_hfns_0 0 1 670 668 buf_x4
xcmpt_abc_11867_new_n430_hfns_1 0 1 669 668 buf_x4
xcmpt_abc_11867_new_n430_hfns_2 0 1 668 671 buf_x4
xfeed_7349 0 1 decap_w0
xfeed_7348 0 1 tie
xfeed_7347 0 1 decap_w0
xfeed_6819 0 1 decap_w0
xfeed_6818 0 1 decap_w0
xfeed_6817 0 1 tie
xfeed_6816 0 1 decap_w0
xfeed_6815 0 1 decap_w0
xfeed_6814 0 1 decap_w0
xfeed_6813 0 1 tie
xfeed_6812 0 1 decap_w0
xfeed_6811 0 1 decap_w0
xfeed_6810 0 1 decap_w0
xfeed_2509 0 1 decap_w0
xfeed_2508 0 1 decap_w0
xfeed_1899 0 1 decap_w0
xfeed_1898 0 1 decap_w0
xfeed_1897 0 1 decap_w0
xfeed_1896 0 1 decap_w0
xfeed_1895 0 1 decap_w0
xfeed_1894 0 1 decap_w0
xfeed_1893 0 1 decap_w0
xfeed_1892 0 1 decap_w0
xfeed_1891 0 1 decap_w0
xfeed_1890 0 1 decap_w0
xsubckt_364_nand2_x0 0 1 385 652 622 nand2_x0
xfeed_14089 0 1 tie
xfeed_14088 0 1 tie
xfeed_14087 0 1 tie
xfeed_14086 0 1 tie
xfeed_14085 0 1 tie
xfeed_14083 0 1 tie
xfeed_14080 0 1 tie
xfeed_13559 0 1 decap_w0
xfeed_13558 0 1 decap_w0
xfeed_13557 0 1 decap_w0
xfeed_13556 0 1 decap_w0
xfeed_13555 0 1 decap_w0
xfeed_13554 0 1 tie
xfeed_13552 0 1 decap_w0
xfeed_13551 0 1 decap_w0
xfeed_13550 0 1 decap_w0
xfeed_7353 0 1 decap_w0
xfeed_7352 0 1 decap_w0
xfeed_7351 0 1 decap_w0
xfeed_7350 0 1 decap_w0
xfeed_3049 0 1 decap_w0
xfeed_3048 0 1 decap_w0
xfeed_3047 0 1 decap_w0
xfeed_3046 0 1 tie
xfeed_3045 0 1 decap_w0
xfeed_3044 0 1 decap_w0
xfeed_3043 0 1 decap_w0
xfeed_3042 0 1 decap_w0
xfeed_3041 0 1 decap_w0
xfeed_3040 0 1 decap_w0
xfeed_2514 0 1 decap_w0
xfeed_2513 0 1 decap_w0
xfeed_2512 0 1 decap_w0
xfeed_2511 0 1 decap_w0
xfeed_2510 0 1 decap_w0
xsubckt_1273_or21nand_x0 0 1 1308 1981 479 1316 or21nand_x0
xsubckt_996_and2_x1 0 1 1533 737 1575 and2_x1
xsubckt_918_and2_x1 0 1 1579 175 1620 and2_x1
xsubckt_856_and4_x1 0 1 1625 780 682 674 670 and4_x1
xsubckt_174_nor3_x0 0 1 584 1920 2055 1921 nor3_x0
xsubckt_613_nand3_x0 0 1 144 2019 184 177 nand3_x0
xsubckt_1651_and3_x1 0 1 943 1070 961 959 and3_x1
xsubckt_1920_dff_x1 0 1 2063 1828 45 dff_x1
xfeed_7359 0 1 decap_w0
xfeed_7358 0 1 decap_w0
xfeed_7357 0 1 tie
xfeed_7356 0 1 decap_w0
xfeed_7355 0 1 decap_w0
xfeed_7354 0 1 decap_w0
xfeed_6829 0 1 decap_w0
xfeed_6828 0 1 decap_w0
xfeed_6827 0 1 decap_w0
xfeed_6826 0 1 decap_w0
xfeed_6825 0 1 decap_w0
xfeed_6824 0 1 tie
xfeed_6823 0 1 decap_w0
xfeed_6822 0 1 decap_w0
xfeed_6821 0 1 decap_w0
xfeed_6820 0 1 decap_w0
xfeed_2519 0 1 decap_w0
xfeed_2518 0 1 decap_w0
xfeed_2517 0 1 decap_w0
xfeed_2516 0 1 decap_w0
xfeed_2515 0 1 decap_w0
xsubckt_1395_nand2_x0 0 1 1196 1203 1198 nand2_x0
xsubckt_1774_or21nand_x0 0 1 820 823 824 832 or21nand_x0
xsubckt_1922_dff_x1 0 1 2061 1826 35 dff_x1
xsubckt_1924_dff_x1 0 1 2059 1824 38 dff_x1
xsubckt_1926_dff_x1 0 1 2073 1822 38 dff_x1
xfeed_14097 0 1 tie
xfeed_14096 0 1 tie
xfeed_14095 0 1 tie
xfeed_14094 0 1 tie
xfeed_14093 0 1 tie
xfeed_14092 0 1 tie
xfeed_14091 0 1 tie
xfeed_14090 0 1 tie
xfeed_13569 0 1 decap_w0
xfeed_13568 0 1 decap_w0
xfeed_13567 0 1 decap_w0
xfeed_13566 0 1 decap_w0
xfeed_13565 0 1 decap_w0
xfeed_13564 0 1 decap_w0
xfeed_13563 0 1 decap_w0
xfeed_13562 0 1 decap_w0
xfeed_13561 0 1 decap_w0
xfeed_13560 0 1 decap_w0
xfeed_7360 0 1 decap_w0
xfeed_3059 0 1 decap_w0
xfeed_3058 0 1 decap_w0
xfeed_3057 0 1 decap_w0
xfeed_3056 0 1 decap_w0
xfeed_3055 0 1 decap_w0
xfeed_3054 0 1 decap_w0
xfeed_3053 0 1 decap_w0
xfeed_3052 0 1 decap_w0
xfeed_3051 0 1 decap_w0
xfeed_3050 0 1 decap_w0
xfeed_2521 0 1 decap_w0
xfeed_2520 0 1 decap_w0
xsubckt_1150_and2_x1 0 1 1410 777 1625 and2_x1
xsubckt_1010_and4_x1 0 1 1519 1531 1528 1524 1520 and4_x1
xsubckt_712_and3_x1 0 1 1752 498 462 399 and3_x1
xsubckt_1735_and21nor_x0 0 1 859 1070 870 1073 and21nor_x0
xsubckt_1809_mux2_x1 0 1 1793 2050 833 773 mux2_x1
xsubckt_1880_dff_x1 0 1 1934 1859 67 dff_x1
xsubckt_1882_dff_x1 0 1 1949 1857 77 dff_x1
xsubckt_1884_dff_x1 0 1 1920 1855 77 dff_x1
xsubckt_1928_dff_x1 0 1 2071 1820 64 dff_x1
xfeed_7369 0 1 decap_w0
xfeed_7368 0 1 decap_w0
xfeed_7367 0 1 decap_w0
xfeed_7366 0 1 decap_w0
xfeed_7365 0 1 decap_w0
xfeed_7364 0 1 decap_w0
xfeed_7363 0 1 decap_w0
xfeed_7362 0 1 decap_w0
xfeed_7361 0 1 decap_w0
xfeed_6839 0 1 decap_w0
xfeed_6838 0 1 decap_w0
xfeed_6837 0 1 decap_w0
xfeed_6836 0 1 decap_w0
xfeed_6835 0 1 decap_w0
xfeed_6834 0 1 decap_w0
xfeed_6833 0 1 decap_w0
xfeed_6832 0 1 decap_w0
xfeed_6831 0 1 tie
xfeed_6830 0 1 decap_w0
xfeed_2529 0 1 decap_w0
xfeed_2528 0 1 decap_w0
xfeed_2527 0 1 tie
xfeed_2526 0 1 decap_w0
xfeed_2525 0 1 decap_w0
xfeed_2524 0 1 decap_w0
xfeed_2523 0 1 decap_w0
xfeed_2522 0 1 decap_w0
xfeed_509 0 1 decap_w0
xfeed_508 0 1 decap_w0
xfeed_507 0 1 decap_w0
xfeed_506 0 1 decap_w0
xfeed_505 0 1 decap_w0
xfeed_504 0 1 decap_w0
xfeed_503 0 1 decap_w0
xfeed_502 0 1 decap_w0
xfeed_501 0 1 decap_w0
xfeed_500 0 1 tie
xsubckt_1886_dff_x1 0 1 1948 1853 77 dff_x1
xsubckt_1888_dff_x1 0 1 1931 1851 77 dff_x1
xfeed_13579 0 1 decap_w0
xfeed_13578 0 1 decap_w0
xfeed_13577 0 1 decap_w0
xfeed_13576 0 1 decap_w0
xfeed_13575 0 1 decap_w0
xfeed_13574 0 1 decap_w0
xfeed_13573 0 1 decap_w0
xfeed_13572 0 1 decap_w0
xfeed_13571 0 1 decap_w0
xfeed_13570 0 1 decap_w0
xfeed_3067 0 1 decap_w0
xfeed_3066 0 1 decap_w0
xfeed_3065 0 1 decap_w0
xfeed_3064 0 1 decap_w0
xfeed_3063 0 1 decap_w0
xfeed_3062 0 1 decap_w0
xfeed_3061 0 1 decap_w0
xfeed_3060 0 1 decap_w0
xsubckt_1146_and2_x1 0 1 1413 1435 1414 and2_x1
xsubckt_1032_and3_x1 0 1 1503 645 637 633 and3_x1
xsubckt_906_nexor2_x0 0 1 1582 1585 1583 nexor2_x0
xsubckt_594_or2_x1 0 1 161 734 212 or2_x1
xsubckt_1464_nand3_x0 0 1 1132 587 579 476 nand3_x0
xsubckt_1669_and2_x1 0 1 925 927 926 and2_x1
xfeed_7379 0 1 decap_w0
xfeed_7378 0 1 decap_w0
xfeed_7377 0 1 decap_w0
xfeed_7376 0 1 decap_w0
xfeed_7375 0 1 decap_w0
xfeed_7374 0 1 decap_w0
xfeed_7373 0 1 decap_w0
xfeed_7372 0 1 decap_w0
xfeed_7371 0 1 decap_w0
xfeed_6849 0 1 decap_w0
xfeed_6848 0 1 decap_w0
xfeed_6846 0 1 decap_w0
xfeed_6845 0 1 decap_w0
xfeed_6844 0 1 decap_w0
xfeed_6843 0 1 decap_w0
xfeed_6842 0 1 decap_w0
xfeed_6840 0 1 decap_w0
xfeed_3069 0 1 decap_w0
xfeed_3068 0 1 decap_w0
xfeed_2539 0 1 decap_w0
xfeed_2538 0 1 decap_w0
xfeed_2537 0 1 decap_w0
xfeed_2536 0 1 decap_w0
xfeed_2535 0 1 decap_w0
xfeed_2534 0 1 decap_w0
xfeed_2533 0 1 decap_w0
xfeed_2532 0 1 decap_w0
xfeed_2531 0 1 decap_w0
xfeed_2530 0 1 decap_w0
xfeed_519 0 1 tie
xfeed_518 0 1 decap_w0
xfeed_517 0 1 decap_w0
xfeed_516 0 1 decap_w0
xfeed_515 0 1 decap_w0
xfeed_514 0 1 decap_w0
xfeed_513 0 1 decap_w0
xfeed_512 0 1 tie
xfeed_511 0 1 decap_w0
xfeed_510 0 1 decap_w0
xsubckt_1180_mux2_x1 0 1 1382 1383 2003 484 mux2_x1
xsubckt_1106_nand3_x0 0 1 1442 663 503 430 nand3_x0
xsubckt_285_and2_x1 0 1 463 466 464 and2_x1
xsubckt_580_and4_x1 0 1 175 187 185 180 179 and4_x1
xsubckt_1284_nand3_x0 0 1 1298 2063 666 657 nand3_x0
xfeed_13589 0 1 decap_w0
xfeed_13588 0 1 decap_w0
xfeed_13587 0 1 decap_w0
xfeed_13586 0 1 decap_w0
xfeed_13585 0 1 decap_w0
xfeed_13584 0 1 decap_w0
xfeed_13583 0 1 decap_w0
xfeed_13582 0 1 decap_w0
xfeed_13581 0 1 decap_w0
xfeed_13580 0 1 decap_w0
xfeed_3074 0 1 decap_w0
xfeed_3073 0 1 decap_w0
xfeed_3072 0 1 decap_w0
xfeed_3071 0 1 decap_w0
xfeed_3070 0 1 decap_w0
xsubckt_1028_and3_x1 0 1 1506 638 632 1545 and3_x1
xsubckt_708_or21nand_x0 0 1 1756 421 608 617 or21nand_x0
xsubckt_322_nand4_x0 0 1 426 643 622 533 524 nand4_x0
xsubckt_1637_nand2_x0 0 1 957 961 959 nand2_x0
xfeed_7389 0 1 decap_w0
xfeed_7388 0 1 decap_w0
xfeed_7387 0 1 decap_w0
xfeed_7386 0 1 decap_w0
xfeed_7385 0 1 decap_w0
xfeed_7384 0 1 decap_w0
xfeed_7383 0 1 decap_w0
xfeed_7382 0 1 decap_w0
xfeed_7381 0 1 decap_w0
xfeed_7380 0 1 decap_w0
xfeed_6859 0 1 decap_w0
xfeed_6858 0 1 decap_w0
xfeed_6857 0 1 decap_w0
xfeed_6856 0 1 decap_w0
xfeed_6855 0 1 decap_w0
xfeed_6854 0 1 decap_w0
xfeed_6853 0 1 decap_w0
xfeed_6852 0 1 decap_w0
xfeed_6851 0 1 decap_w0
xfeed_3079 0 1 decap_w0
xfeed_3078 0 1 decap_w0
xfeed_3077 0 1 decap_w0
xfeed_3076 0 1 decap_w0
xfeed_3075 0 1 decap_w0
xfeed_2549 0 1 decap_w0
xfeed_2548 0 1 decap_w0
xfeed_2547 0 1 decap_w0
xfeed_2546 0 1 decap_w0
xfeed_2545 0 1 decap_w0
xfeed_2544 0 1 decap_w0
xfeed_2543 0 1 decap_w0
xfeed_2542 0 1 decap_w0
xfeed_2541 0 1 decap_w0
xfeed_2540 0 1 decap_w0
xfeed_529 0 1 decap_w0
xfeed_528 0 1 decap_w0
xfeed_527 0 1 decap_w0
xfeed_526 0 1 tie
xfeed_525 0 1 decap_w0
xfeed_524 0 1 decap_w0
xfeed_523 0 1 decap_w0
xfeed_522 0 1 decap_w0
xfeed_521 0 1 decap_w0
xfeed_520 0 1 decap_w0
xsubckt_1176_mux2_x1 0 1 1386 1389 484 1392 mux2_x1
xsubckt_611_or21nand_x0 0 1 2081 146 153 206 or21nand_x0
xsubckt_1457_nand2_x0 0 1 1139 756 548 nand2_x0
xfeed_13599 0 1 decap_w0
xfeed_13598 0 1 decap_w0
xfeed_13597 0 1 decap_w0
xfeed_13596 0 1 decap_w0
xfeed_13595 0 1 decap_w0
xfeed_13594 0 1 decap_w0
xfeed_13593 0 1 decap_w0
xfeed_13592 0 1 decap_w0
xfeed_13591 0 1 decap_w0
xfeed_13590 0 1 decap_w0
xfeed_8009 0 1 decap_w0
xfeed_8008 0 1 decap_w0
xfeed_8007 0 1 decap_w0
xfeed_8006 0 1 decap_w0
xfeed_8005 0 1 decap_w0
xfeed_8004 0 1 decap_w0
xfeed_8003 0 1 decap_w0
xfeed_8002 0 1 decap_w0
xfeed_8001 0 1 decap_w0
xfeed_8000 0 1 decap_w0
xfeed_3081 0 1 decap_w0
xfeed_3080 0 1 decap_w0
xsubckt_1_inv_x0 0 1 785 1986 inv_x0
xsubckt_3_inv_x0 0 1 783 2012 inv_x0
xsubckt_115_and2_x1 0 1 653 659 654 and2_x1
xsubckt_1367_nand2_x0 0 1 1222 1229 1224 nand2_x0
xsubckt_1407_and2_x1 0 1 1185 1191 1186 and2_x1
xfeed_7399 0 1 decap_w0
xfeed_7398 0 1 decap_w0
xfeed_7397 0 1 decap_w0
xfeed_7396 0 1 decap_w0
xfeed_7395 0 1 decap_w0
xfeed_7394 0 1 decap_w0
xfeed_7393 0 1 decap_w0
xfeed_7392 0 1 decap_w0
xfeed_7391 0 1 decap_w0
xfeed_7390 0 1 decap_w0
xfeed_6869 0 1 tie
xfeed_6868 0 1 decap_w0
xfeed_6867 0 1 decap_w0
xfeed_6866 0 1 decap_w0
xfeed_6865 0 1 decap_w0
xfeed_6864 0 1 decap_w0
xfeed_6862 0 1 tie
xfeed_6861 0 1 decap_w0
xfeed_6860 0 1 decap_w0
xfeed_3089 0 1 decap_w0
xfeed_3088 0 1 decap_w0
xfeed_3087 0 1 decap_w0
xfeed_3086 0 1 decap_w0
xfeed_3085 0 1 decap_w0
xfeed_3084 0 1 decap_w0
xfeed_3083 0 1 decap_w0
xfeed_3082 0 1 tie
xfeed_2559 0 1 decap_w0
xfeed_2558 0 1 decap_w0
xfeed_2557 0 1 decap_w0
xfeed_2556 0 1 decap_w0
xfeed_2555 0 1 decap_w0
xfeed_2554 0 1 decap_w0
xfeed_2553 0 1 decap_w0
xfeed_2552 0 1 decap_w0
xfeed_2551 0 1 decap_w0
xfeed_2550 0 1 decap_w0
xfeed_539 0 1 decap_w0
xfeed_538 0 1 decap_w0
xfeed_537 0 1 decap_w0
xfeed_536 0 1 decap_w0
xfeed_535 0 1 decap_w0
xfeed_534 0 1 decap_w0
xfeed_533 0 1 decap_w0
xfeed_532 0 1 decap_w0
xfeed_531 0 1 decap_w0
xfeed_530 0 1 decap_w0
xsubckt_5_inv_x0 0 1 781 1959 inv_x0
xsubckt_7_inv_x0 0 1 779 1934 inv_x0
xsubckt_9_inv_x0 0 1 777 1955 inv_x0
xsubckt_493_nand3_x0 0 1 258 610 556 418 nand3_x0
xsubckt_1393_and2_x1 0 1 1198 1202 1199 and2_x1
xfeed_8019 0 1 decap_w0
xfeed_8018 0 1 decap_w0
xfeed_8017 0 1 decap_w0
xfeed_8016 0 1 decap_w0
xfeed_8015 0 1 decap_w0
xfeed_8014 0 1 decap_w0
xfeed_8013 0 1 decap_w0
xfeed_8012 0 1 decap_w0
xfeed_8011 0 1 decap_w0
xfeed_8010 0 1 decap_w0
xsubckt_981_and2_x1 0 1 1546 1550 1547 and2_x1
xsubckt_796_nor2_x0 0 1 1676 1758 1677 nor2_x0
xsubckt_1372_or21nand_x0 0 1 1805 1230 1220 1218 or21nand_x0
xsubckt_1440_nand2_x0 0 1 1155 775 1975 nand2_x0
xfeed_6879 0 1 decap_w0
xfeed_6878 0 1 decap_w0
xfeed_6877 0 1 decap_w0
xfeed_6876 0 1 decap_w0
xfeed_6875 0 1 decap_w0
xfeed_6874 0 1 decap_w0
xfeed_6873 0 1 decap_w0
xfeed_6872 0 1 decap_w0
xfeed_6871 0 1 decap_w0
xfeed_6870 0 1 decap_w0
xfeed_3099 0 1 decap_w0
xfeed_3098 0 1 decap_w0
xfeed_3097 0 1 decap_w0
xfeed_3096 0 1 decap_w0
xfeed_3095 0 1 decap_w0
xfeed_3094 0 1 decap_w0
xfeed_3093 0 1 decap_w0
xfeed_3092 0 1 decap_w0
xfeed_3091 0 1 decap_w0
xfeed_3090 0 1 decap_w0
xfeed_2569 0 1 decap_w0
xfeed_2568 0 1 decap_w0
xfeed_2567 0 1 tie
xfeed_2566 0 1 decap_w0
xfeed_2565 0 1 decap_w0
xfeed_2564 0 1 decap_w0
xfeed_2563 0 1 decap_w0
xfeed_2562 0 1 decap_w0
xfeed_2561 0 1 decap_w0
xfeed_2560 0 1 decap_w0
xfeed_549 0 1 decap_w0
xfeed_548 0 1 decap_w0
xfeed_547 0 1 decap_w0
xfeed_546 0 1 decap_w0
xfeed_545 0 1 decap_w0
xfeed_544 0 1 tie
xfeed_543 0 1 decap_w0
xfeed_542 0 1 decap_w0
xfeed_541 0 1 decap_w0
xfeed_540 0 1 decap_w0
xsubckt_1029_and21nor_x0 0 1 1505 783 659 624 and21nor_x0
xsubckt_756_nand2_x0 0 1 2097 1718 1712 nand2_x0
xsubckt_392_and4_x1 0 1 357 533 524 518 360 and4_x1
xfeed_8029 0 1 decap_w0
xfeed_8028 0 1 decap_w0
xfeed_8027 0 1 decap_w0
xfeed_8026 0 1 decap_w0
xfeed_8025 0 1 decap_w0
xfeed_8024 0 1 decap_w0
xfeed_8023 0 1 decap_w0
xfeed_8022 0 1 decap_w0
xfeed_8021 0 1 decap_w0
xfeed_8020 0 1 decap_w0
xsubckt_1606_and4_x1 0 1 988 1999 1128 1098 1097 and4_x1
xsubckt_1632_and3_x1 0 1 962 1973 681 595 and3_x1
xfeed_6889 0 1 decap_w0
xfeed_6887 0 1 decap_w0
xfeed_6886 0 1 decap_w0
xfeed_6885 0 1 decap_w0
xfeed_6884 0 1 decap_w0
xfeed_6883 0 1 decap_w0
xfeed_6882 0 1 decap_w0
xfeed_6881 0 1 decap_w0
xfeed_6880 0 1 decap_w0
xfeed_2579 0 1 tie
xfeed_2578 0 1 decap_w0
xfeed_2577 0 1 decap_w0
xfeed_2576 0 1 decap_w0
xfeed_2575 0 1 decap_w0
xfeed_2574 0 1 tie
xfeed_2573 0 1 decap_w0
xfeed_2572 0 1 decap_w0
xfeed_2571 0 1 decap_w0
xfeed_2570 0 1 decap_w0
xfeed_559 0 1 decap_w0
xfeed_558 0 1 decap_w0
xfeed_557 0 1 decap_w0
xfeed_556 0 1 tie
xfeed_555 0 1 decap_w0
xfeed_553 0 1 decap_w0
xfeed_552 0 1 decap_w0
xfeed_551 0 1 tie
xfeed_550 0 1 decap_w0
xsubckt_933_mux2_x1 0 1 1884 2024 1593 1578 mux2_x1
xfeed_13709 0 1 decap_w0
xfeed_13708 0 1 decap_w0
xfeed_13707 0 1 decap_w0
xfeed_13706 0 1 decap_w0
xfeed_13705 0 1 decap_w0
xfeed_13704 0 1 decap_w0
xfeed_13703 0 1 decap_w0
xfeed_13702 0 1 decap_w0
xfeed_13701 0 1 decap_w0
xfeed_13700 0 1 decap_w0
xfeed_8039 0 1 decap_w0
xfeed_8038 0 1 decap_w0
xfeed_8037 0 1 decap_w0
xfeed_8036 0 1 decap_w0
xfeed_8035 0 1 decap_w0
xfeed_8034 0 1 decap_w0
xfeed_8033 0 1 decap_w0
xfeed_8032 0 1 decap_w0
xfeed_8031 0 1 decap_w0
xfeed_8030 0 1 decap_w0
xfeed_7500 0 1 decap_w0
xsubckt_1076_nand3_x0 0 1 1468 623 519 1515 nand3_x0
xsubckt_292_nand4_x0 0 1 456 1929 715 680 599 nand4_x0
xsubckt_198_or21nand_x0 0 1 560 687 619 561 or21nand_x0
xsubckt_128_nand2_x0 0 1 640 785 2003 nand2_x0
xsubckt_396_nand2_x0 0 1 353 563 354 nand2_x0
xsubckt_1572_or21nand_x0 0 1 1022 1025 1118 762 or21nand_x0
xfeed_7509 0 1 tie
xfeed_7508 0 1 decap_w0
xfeed_7507 0 1 decap_w0
xfeed_7506 0 1 decap_w0
xfeed_7505 0 1 decap_w0
xfeed_7504 0 1 decap_w0
xfeed_7503 0 1 decap_w0
xfeed_7502 0 1 tie
xfeed_7501 0 1 decap_w0
xfeed_6899 0 1 decap_w0
xfeed_6898 0 1 decap_w0
xfeed_6897 0 1 decap_w0
xfeed_6896 0 1 decap_w0
xfeed_6895 0 1 tie
xfeed_6894 0 1 decap_w0
xfeed_6893 0 1 decap_w0
xfeed_6892 0 1 decap_w0
xfeed_6891 0 1 decap_w0
xfeed_6890 0 1 decap_w0
xfeed_2589 0 1 decap_w0
xfeed_2588 0 1 decap_w0
xfeed_2587 0 1 decap_w0
xfeed_2586 0 1 tie
xfeed_2585 0 1 decap_w0
xfeed_2584 0 1 decap_w0
xfeed_2583 0 1 decap_w0
xfeed_2582 0 1 decap_w0
xfeed_2581 0 1 decap_w0
xfeed_2580 0 1 decap_w0
xfeed_569 0 1 decap_w0
xfeed_568 0 1 decap_w0
xfeed_567 0 1 decap_w0
xfeed_566 0 1 decap_w0
xfeed_565 0 1 tie
xfeed_564 0 1 decap_w0
xfeed_563 0 1 decap_w0
xfeed_562 0 1 decap_w0
xfeed_561 0 1 decap_w0
xfeed_560 0 1 decap_w0
xsubckt_1229_and21nor_x0 0 1 1335 576 1342 1336 and21nor_x0
xsubckt_999_nand4_x0 0 1 1530 645 637 633 525 nand4_x0
xsubckt_929_mux2_x1 0 1 1888 2028 1612 1578 mux2_x1
xsubckt_1368_or21nand_x0 0 1 1221 1223 1235 1244 or21nand_x0
xfeed_13719 0 1 decap_w0
xfeed_13718 0 1 decap_w0
xfeed_13717 0 1 decap_w0
xfeed_13716 0 1 decap_w0
xfeed_13715 0 1 decap_w0
xfeed_13714 0 1 decap_w0
xfeed_13713 0 1 decap_w0
xfeed_13712 0 1 decap_w0
xfeed_13711 0 1 decap_w0
xfeed_13710 0 1 decap_w0
xfeed_8046 0 1 decap_w0
xfeed_8045 0 1 decap_w0
xfeed_8044 0 1 decap_w0
xfeed_8043 0 1 decap_w0
xfeed_8042 0 1 decap_w0
xfeed_8041 0 1 decap_w0
xfeed_8040 0 1 tie
xfeed_3207 0 1 tie
xfeed_3206 0 1 decap_w0
xfeed_3205 0 1 decap_w0
xfeed_3204 0 1 decap_w0
xfeed_3203 0 1 decap_w0
xfeed_3202 0 1 decap_w0
xfeed_3201 0 1 decap_w0
xfeed_3200 0 1 decap_w0
xsubckt_1087_and3_x1 0 1 1458 1531 1465 1459 and3_x1
xsubckt_13_inv_x0 0 1 769 2053 inv_x0
xsubckt_11_inv_x0 0 1 771 10 inv_x0
xfeed_8049 0 1 decap_w0
xfeed_8048 0 1 decap_w0
xfeed_8047 0 1 decap_w0
xfeed_7519 0 1 decap_w0
xfeed_7518 0 1 decap_w0
xfeed_7517 0 1 decap_w0
xfeed_7516 0 1 tie
xfeed_7515 0 1 decap_w0
xfeed_7514 0 1 decap_w0
xfeed_7513 0 1 decap_w0
xfeed_7512 0 1 decap_w0
xfeed_7511 0 1 decap_w0
xfeed_7510 0 1 decap_w0
xfeed_3209 0 1 decap_w0
xfeed_3208 0 1 decap_w0
xfeed_2599 0 1 decap_w0
xfeed_2598 0 1 decap_w0
xfeed_2597 0 1 decap_w0
xfeed_2596 0 1 decap_w0
xfeed_2595 0 1 decap_w0
xfeed_2594 0 1 decap_w0
xfeed_2593 0 1 tie
xfeed_2592 0 1 decap_w0
xfeed_2591 0 1 decap_w0
xfeed_2590 0 1 decap_w0
xfeed_576 0 1 decap_w0
xfeed_575 0 1 decap_w0
xfeed_574 0 1 decap_w0
xfeed_573 0 1 decap_w0
xfeed_572 0 1 decap_w0
xfeed_571 0 1 decap_w0
xfeed_570 0 1 decap_w0
xsubckt_1145_nand4_x0 0 1 1414 679 673 669 1415 nand4_x0
xsubckt_1069_nand2_x0 0 1 1474 1530 1475 nand2_x0
xsubckt_19_inv_x0 0 1 763 2049 inv_x0
xsubckt_17_inv_x0 0 1 765 2051 inv_x0
xsubckt_15_inv_x0 0 1 767 1964 inv_x0
xsubckt_561_and4_x1 0 1 194 537 503 325 200 and4_x1
xsubckt_1298_or2_x1 0 1 1285 1289 1286 or2_x1
xsubckt_1412_nand2_x0 0 1 1180 1917 1183 nand2_x0
xfeed_13729 0 1 decap_w0
xfeed_13728 0 1 decap_w0
xfeed_13727 0 1 decap_w0
xfeed_13726 0 1 decap_w0
xfeed_13725 0 1 decap_w0
xfeed_13724 0 1 decap_w0
xfeed_13723 0 1 decap_w0
xfeed_13722 0 1 decap_w0
xfeed_13721 0 1 decap_w0
xfeed_13720 0 1 decap_w0
xfeed_8053 0 1 decap_w0
xfeed_8052 0 1 tie
xfeed_8051 0 1 decap_w0
xfeed_8050 0 1 decap_w0
xfeed_3214 0 1 decap_w0
xfeed_3213 0 1 decap_w0
xfeed_3212 0 1 decap_w0
xfeed_3211 0 1 decap_w0
xfeed_3210 0 1 decap_w0
xfeed_579 0 1 decap_w0
xfeed_578 0 1 decap_w0
xfeed_577 0 1 decap_w0
xsubckt_1171_nor3_x0 0 1 1391 1934 1963 1955 nor3_x0
xsubckt_1157_mux2_x1 0 1 1834 1404 1985 1405 mux2_x1
xsubckt_728_nand2_x0 0 1 1736 2003 1746 nand2_x0
xsubckt_1772_or21nand_x0 0 1 822 939 938 835 or21nand_x0
xfeed_8059 0 1 tie
xfeed_8058 0 1 decap_w0
xfeed_8057 0 1 decap_w0
xfeed_8056 0 1 decap_w0
xfeed_8055 0 1 decap_w0
xfeed_8054 0 1 decap_w0
xfeed_7529 0 1 decap_w0
xfeed_7528 0 1 decap_w0
xfeed_7527 0 1 decap_w0
xfeed_7526 0 1 decap_w0
xfeed_7525 0 1 decap_w0
xfeed_7524 0 1 decap_w0
xfeed_7523 0 1 tie
xfeed_7522 0 1 decap_w0
xfeed_7521 0 1 decap_w0
xfeed_7520 0 1 decap_w0
xfeed_3219 0 1 decap_w0
xfeed_3218 0 1 decap_w0
xfeed_3217 0 1 decap_w0
xfeed_3216 0 1 decap_w0
xfeed_3215 0 1 decap_w0
xfeed_583 0 1 decap_w0
xfeed_582 0 1 decap_w0
xfeed_581 0 1 decap_w0
xfeed_580 0 1 decap_w0
xsubckt_548_nand2_x0 0 1 206 600 209 nand2_x0
xfeed_13739 0 1 decap_w0
xfeed_13738 0 1 decap_w0
xfeed_13737 0 1 decap_w0
xfeed_13736 0 1 decap_w0
xfeed_13735 0 1 decap_w0
xfeed_13734 0 1 decap_w0
xfeed_13733 0 1 decap_w0
xfeed_13732 0 1 decap_w0
xfeed_13731 0 1 tie
xfeed_13730 0 1 decap_w0
xfeed_8060 0 1 decap_w0
xfeed_3221 0 1 tie
xfeed_3220 0 1 decap_w0
xfeed_589 0 1 decap_w0
xfeed_588 0 1 decap_w0
xfeed_587 0 1 decap_w0
xfeed_586 0 1 decap_w0
xfeed_585 0 1 decap_w0
xfeed_584 0 1 decap_w0
xsubckt_1065_mux2_x1 0 1 1852 1478 1932 1576 mux2_x1
xsubckt_755_nor3_x0 0 1 1712 1717 1716 1713 nor3_x0
xsubckt_711_nand2_x0 0 1 1753 498 462 nand2_x0
xsubckt_458_nand2_x0 0 1 292 368 356 nand2_x0
xsubckt_491_and3_x1 0 1 260 616 556 418 and3_x1
xsubckt_606_or21nand_x0 0 1 150 1965 436 167 or21nand_x0
xsubckt_1588_mux2_x1 0 1 1006 1009 1012 1020 mux2_x1
xfeed_8069 0 1 decap_w0
xfeed_8068 0 1 decap_w0
xfeed_8067 0 1 decap_w0
xfeed_8066 0 1 tie
xfeed_8065 0 1 decap_w0
xfeed_8064 0 1 decap_w0
xfeed_8063 0 1 decap_w0
xfeed_8062 0 1 decap_w0
xfeed_8061 0 1 decap_w0
xfeed_7539 0 1 decap_w0
xfeed_7538 0 1 decap_w0
xfeed_7537 0 1 decap_w0
xfeed_7536 0 1 decap_w0
xfeed_7535 0 1 decap_w0
xfeed_7534 0 1 tie
xfeed_7533 0 1 decap_w0
xfeed_7532 0 1 decap_w0
xfeed_7531 0 1 decap_w0
xfeed_7530 0 1 decap_w0
xfeed_3228 0 1 decap_w0
xfeed_3227 0 1 decap_w0
xfeed_3226 0 1 decap_w0
xfeed_3225 0 1 decap_w0
xfeed_3224 0 1 decap_w0
xfeed_3223 0 1 decap_w0
xfeed_3222 0 1 decap_w0
xfeed_590 0 1 decap_w0
xsubckt_899_nexor2_x0 0 1 1588 760 1592 nexor2_x0
xsubckt_354_nand4_x0 0 1 394 1917 771 680 405 nand4_x0
xfeed_13749 0 1 decap_w0
xfeed_13748 0 1 tie
xfeed_13747 0 1 decap_w0
xfeed_13746 0 1 decap_w0
xfeed_13745 0 1 decap_w0
xfeed_13744 0 1 decap_w0
xfeed_13743 0 1 tie
xfeed_13742 0 1 decap_w0
xfeed_13741 0 1 decap_w0
xfeed_13740 0 1 decap_w0
xfeed_599 0 1 decap_w0
xfeed_598 0 1 decap_w0
xfeed_597 0 1 decap_w0
xfeed_596 0 1 decap_w0
xfeed_595 0 1 decap_w0
xfeed_594 0 1 decap_w0
xfeed_593 0 1 decap_w0
xfeed_592 0 1 decap_w0
xfeed_591 0 1 decap_w0
xsubckt_1256_and3_x1 0 1 1324 1332 1327 1325 and3_x1
xsubckt_373_and4_x1 0 1 376 532 530 518 384 and4_x1
xsubckt_598_or21nand_x0 0 1 2082 158 169 206 or21nand_x0
xsubckt_1475_nand4_x0 0 1 1121 1768 1360 1124 1123 nand4_x0
xfeed_8079 0 1 decap_w0
xfeed_8078 0 1 decap_w0
xfeed_8077 0 1 tie
xfeed_8076 0 1 decap_w0
xfeed_8075 0 1 decap_w0
xfeed_8074 0 1 decap_w0
xfeed_8073 0 1 decap_w0
xfeed_8072 0 1 decap_w0
xfeed_8071 0 1 decap_w0
xfeed_8070 0 1 tie
xfeed_7549 0 1 decap_w0
xfeed_7548 0 1 decap_w0
xfeed_7547 0 1 decap_w0
xfeed_7546 0 1 decap_w0
xfeed_7545 0 1 decap_w0
xfeed_7544 0 1 decap_w0
xfeed_7543 0 1 decap_w0
xfeed_7542 0 1 decap_w0
xfeed_7541 0 1 tie
xfeed_7540 0 1 decap_w0
xfeed_3239 0 1 decap_w0
xfeed_3238 0 1 decap_w0
xfeed_3237 0 1 decap_w0
xfeed_3236 0 1 tie
xfeed_3235 0 1 decap_w0
xfeed_3234 0 1 decap_w0
xfeed_3233 0 1 decap_w0
xfeed_3232 0 1 decap_w0
xfeed_3231 0 1 decap_w0
xfeed_2709 0 1 decap_w0
xfeed_2708 0 1 decap_w0
xfeed_2707 0 1 decap_w0
xfeed_2706 0 1 decap_w0
xfeed_2705 0 1 decap_w0
xfeed_2704 0 1 decap_w0
xfeed_2703 0 1 decap_w0
xfeed_2702 0 1 decap_w0
xfeed_2701 0 1 decap_w0
xfeed_2700 0 1 decap_w0
xsubckt_1204_and2_x1 0 1 1360 193 1769 and2_x1
xsubckt_162_nor2_x0 0 1 599 1927 1928 nor2_x0
xsubckt_435_and2_x1 0 1 315 317 316 and2_x1
xsubckt_1399_nand2_x0 0 1 1803 1204 1193 nand2_x0
xsubckt_1742_nand2_x0 0 1 852 1082 1077 nand2_x0
xsubckt_1931_dff_x1 0 1 2068 1817 64 dff_x1
xsubckt_1933_dff_x1 0 1 2066 1815 58 dff_x1
xfeed_13759 0 1 decap_w0
xfeed_13758 0 1 decap_w0
xfeed_13757 0 1 decap_w0
xfeed_13756 0 1 decap_w0
xfeed_13755 0 1 decap_w0
xfeed_13754 0 1 decap_w0
xfeed_13753 0 1 decap_w0
xfeed_13752 0 1 decap_w0
xfeed_13751 0 1 decap_w0
xfeed_13750 0 1 decap_w0
xsubckt_866_and2_x1 0 1 1616 1962 1617 and2_x1
xsubckt_317_and3_x1 0 1 431 463 453 432 and3_x1
xsubckt_607_nor2_x0 0 1 149 733 212 nor2_x0
xsubckt_1891_dff_x1 0 1 1939 1848 54 dff_x1
xsubckt_1935_dff_x1 0 1 1981 1813 51 dff_x1
xsubckt_1937_dff_x1 0 1 1973 1811 41 dff_x1
xsubckt_1939_dff_x1 0 1 1971 1809 38 dff_x1
xfeed_8089 0 1 decap_w0
xfeed_8088 0 1 decap_w0
xfeed_8087 0 1 decap_w0
xfeed_8085 0 1 decap_w0
xfeed_8084 0 1 decap_w0
xfeed_8083 0 1 decap_w0
xfeed_8082 0 1 decap_w0
xfeed_8081 0 1 decap_w0
xfeed_8080 0 1 decap_w0
xfeed_7559 0 1 decap_w0
xfeed_7558 0 1 decap_w0
xfeed_7557 0 1 decap_w0
xfeed_7556 0 1 decap_w0
xfeed_7555 0 1 decap_w0
xfeed_7554 0 1 decap_w0
xfeed_7553 0 1 decap_w0
xfeed_7552 0 1 decap_w0
xfeed_7551 0 1 decap_w0
xfeed_7550 0 1 decap_w0
xfeed_3249 0 1 decap_w0
xfeed_3248 0 1 decap_w0
xfeed_3247 0 1 decap_w0
xfeed_3246 0 1 decap_w0
xfeed_3245 0 1 decap_w0
xfeed_3244 0 1 decap_w0
xfeed_3243 0 1 decap_w0
xfeed_3242 0 1 decap_w0
xfeed_3241 0 1 decap_w0
xfeed_3240 0 1 decap_w0
xfeed_2719 0 1 decap_w0
xfeed_2718 0 1 decap_w0
xfeed_2717 0 1 decap_w0
xfeed_2716 0 1 tie
xfeed_2714 0 1 decap_w0
xfeed_2713 0 1 decap_w0
xfeed_2712 0 1 decap_w0
xfeed_2711 0 1 decap_w0
xfeed_2710 0 1 decap_w0
xsubckt_914_mux2_x1 0 1 1901 1599 2041 1580 mux2_x1
xsubckt_277_and4_x1 0 1 471 492 486 477 472 and4_x1
xsubckt_257_nand3_x0 0 1 494 714 1928 589 nand3_x0
xsubckt_600_nand3_x0 0 1 156 2020 184 177 nand3_x0
xsubckt_1893_dff_x1 0 1 2010 2002 64 dff_x1
xsubckt_1895_dff_x1 0 1 2008 2000 64 dff_x1
xsubckt_1897_dff_x1 0 1 2006 1998 58 dff_x1
xfeed_13769 0 1 decap_w0
xfeed_13768 0 1 decap_w0
xfeed_13767 0 1 decap_w0
xfeed_13766 0 1 decap_w0
xfeed_13765 0 1 decap_w0
xfeed_13764 0 1 decap_w0
xfeed_13763 0 1 decap_w0
xfeed_13762 0 1 decap_w0
xfeed_13761 0 1 decap_w0
xfeed_13760 0 1 decap_w0
xsubckt_1234_mux2_x1 0 1 1827 2097 2062 1334 mux2_x1
xsubckt_774_and2_x1 0 1 1696 2047 1748 and2_x1
xsubckt_649_or2_x1 0 1 110 729 212 or2_x1
xsubckt_167_nand3_x0 0 1 591 714 616 613 nand3_x0
xsubckt_397_or21nand_x0 0 1 352 438 420 614 or21nand_x0
xsubckt_420_nand3_x0 0 1 329 680 558 447 nand3_x0
xsubckt_1721_nand3_x0 0 1 873 1982 678 595 nand3_x0
xsubckt_1899_dff_x1 0 1 2004 1996 38 dff_x1
xfeed_8099 0 1 decap_w0
xfeed_8098 0 1 decap_w0
xfeed_8097 0 1 decap_w0
xfeed_8096 0 1 decap_w0
xfeed_8095 0 1 decap_w0
xfeed_8094 0 1 decap_w0
xfeed_8093 0 1 decap_w0
xfeed_8092 0 1 decap_w0
xfeed_8091 0 1 decap_w0
xfeed_8090 0 1 decap_w0
xfeed_7569 0 1 decap_w0
xfeed_7568 0 1 decap_w0
xfeed_7567 0 1 decap_w0
xfeed_7566 0 1 decap_w0
xfeed_7565 0 1 decap_w0
xfeed_7564 0 1 decap_w0
xfeed_7563 0 1 decap_w0
xfeed_7562 0 1 decap_w0
xfeed_7561 0 1 decap_w0
xfeed_7560 0 1 decap_w0
xfeed_3259 0 1 decap_w0
xfeed_3258 0 1 decap_w0
xfeed_3256 0 1 decap_w0
xfeed_3255 0 1 decap_w0
xfeed_3254 0 1 decap_w0
xfeed_3253 0 1 decap_w0
xfeed_3252 0 1 decap_w0
xfeed_3251 0 1 decap_w0
xfeed_3250 0 1 decap_w0
xfeed_2729 0 1 decap_w0
xfeed_2728 0 1 decap_w0
xfeed_2727 0 1 decap_w0
xfeed_2726 0 1 decap_w0
xfeed_2725 0 1 decap_w0
xfeed_2724 0 1 decap_w0
xfeed_2723 0 1 decap_w0
xfeed_2722 0 1 decap_w0
xfeed_2721 0 1 decap_w0
xfeed_2720 0 1 decap_w0
xfeed_709 0 1 tie
xfeed_708 0 1 decap_w0
xfeed_707 0 1 decap_w0
xfeed_706 0 1 decap_w0
xfeed_705 0 1 decap_w0
xfeed_703 0 1 decap_w0
xfeed_702 0 1 decap_w0
xfeed_701 0 1 decap_w0
xfeed_700 0 1 decap_w0
xsubckt_1517_and3_x1 0 1 1079 1961 682 490 and3_x1
xfeed_13779 0 1 decap_w0
xfeed_13778 0 1 decap_w0
xfeed_13777 0 1 decap_w0
xfeed_13776 0 1 decap_w0
xfeed_13775 0 1 decap_w0
xfeed_13774 0 1 decap_w0
xfeed_13773 0 1 decap_w0
xfeed_13772 0 1 decap_w0
xfeed_13771 0 1 decap_w0
xfeed_13770 0 1 decap_w0
xfeed_7579 0 1 decap_w0
xfeed_7578 0 1 tie
xfeed_7577 0 1 decap_w0
xfeed_7576 0 1 decap_w0
xfeed_7575 0 1 decap_w0
xfeed_7574 0 1 decap_w0
xfeed_7573 0 1 decap_w0
xfeed_7572 0 1 decap_w0
xfeed_7571 0 1 decap_w0
xfeed_7570 0 1 decap_w0
xfeed_3268 0 1 decap_w0
xfeed_3267 0 1 decap_w0
xfeed_3266 0 1 decap_w0
xfeed_3265 0 1 decap_w0
xfeed_3264 0 1 decap_w0
xfeed_3262 0 1 decap_w0
xfeed_3261 0 1 decap_w0
xfeed_3260 0 1 decap_w0
xfeed_2739 0 1 decap_w0
xfeed_2738 0 1 decap_w0
xfeed_2737 0 1 decap_w0
xfeed_2736 0 1 decap_w0
xfeed_2735 0 1 decap_w0
xfeed_2734 0 1 decap_w0
xfeed_2733 0 1 decap_w0
xfeed_2732 0 1 decap_w0
xfeed_2731 0 1 decap_w0
xfeed_2730 0 1 decap_w0
xfeed_716 0 1 decap_w0
xfeed_715 0 1 decap_w0
xfeed_714 0 1 decap_w0
xfeed_713 0 1 decap_w0
xfeed_712 0 1 decap_w0
xfeed_711 0 1 decap_w0
xfeed_710 0 1 decap_w0
xsubckt_859_and21nor_x0 0 1 1622 544 447 617 and21nor_x0
xsubckt_605_or21nand_x0 0 1 151 2052 601 163 or21nand_x0
xsubckt_1311_and4_x1 0 1 1273 1302 1293 1285 1275 and4_x1
xfeed_13789 0 1 decap_w0
xfeed_13788 0 1 decap_w0
xfeed_13787 0 1 decap_w0
xfeed_13786 0 1 decap_w0
xfeed_13785 0 1 decap_w0
xfeed_13784 0 1 decap_w0
xfeed_13783 0 1 decap_w0
xfeed_13782 0 1 decap_w0
xfeed_13781 0 1 decap_w0
xfeed_13780 0 1 decap_w0
xfeed_719 0 1 tie
xfeed_718 0 1 decap_w0
xfeed_717 0 1 decap_w0
xsubckt_590_and2_x1 0 1 165 435 166 and2_x1
xsubckt_1570_or21nand_x0 0 1 1024 1642 1116 691 or21nand_x0
xsubckt_1628_and21nor_x0 0 1 966 967 1117 2050 and21nor_x0
xfeed_7589 0 1 decap_w0
xfeed_7588 0 1 decap_w0
xfeed_7587 0 1 decap_w0
xfeed_7586 0 1 decap_w0
xfeed_7585 0 1 decap_w0
xfeed_7584 0 1 decap_w0
xfeed_7583 0 1 decap_w0
xfeed_7582 0 1 decap_w0
xfeed_7581 0 1 decap_w0
xfeed_7580 0 1 decap_w0
xfeed_3279 0 1 decap_w0
xfeed_3277 0 1 decap_w0
xfeed_3276 0 1 decap_w0
xfeed_3275 0 1 decap_w0
xfeed_3274 0 1 decap_w0
xfeed_3273 0 1 decap_w0
xfeed_3271 0 1 decap_w0
xfeed_3270 0 1 decap_w0
xfeed_2749 0 1 decap_w0
xfeed_2748 0 1 decap_w0
xfeed_2747 0 1 decap_w0
xfeed_2746 0 1 decap_w0
xfeed_2745 0 1 decap_w0
xfeed_2744 0 1 decap_w0
xfeed_2743 0 1 decap_w0
xfeed_2742 0 1 decap_w0
xfeed_2741 0 1 decap_w0
xfeed_2740 0 1 decap_w0
xfeed_723 0 1 decap_w0
xfeed_722 0 1 decap_w0
xfeed_721 0 1 decap_w0
xfeed_720 0 1 decap_w0
xsubckt_1003_nand3_x0 0 1 1526 532 360 1527 nand3_x0
xsubckt_196_or21nand_x0 0 1 562 778 572 564 or21nand_x0
xsubckt_497_nand3_x0 0 1 254 568 556 405 nand3_x0
xsubckt_512_and2_x1 0 1 239 388 240 and2_x1
xfeed_13799 0 1 decap_w0
xfeed_13798 0 1 decap_w0
xfeed_13797 0 1 decap_w0
xfeed_13796 0 1 decap_w0
xfeed_13795 0 1 decap_w0
xfeed_13794 0 1 decap_w0
xfeed_13793 0 1 decap_w0
xfeed_13792 0 1 decap_w0
xfeed_13791 0 1 decap_w0
xfeed_13790 0 1 decap_w0
xfeed_8200 0 1 decap_w0
xfeed_729 0 1 decap_w0
xfeed_728 0 1 decap_w0
xfeed_727 0 1 decap_w0
xfeed_726 0 1 decap_w0
xfeed_725 0 1 decap_w0
xfeed_724 0 1 decap_w0
xsubckt_96_mux2_x1 0 1 691 718 717 773 mux2_x1
xsubckt_143_nand2_x0 0 1 625 785 1996 nand2_x0
xfeed_8209 0 1 decap_w0
xfeed_8208 0 1 decap_w0
xfeed_8207 0 1 decap_w0
xfeed_8206 0 1 decap_w0
xfeed_8205 0 1 decap_w0
xfeed_8204 0 1 decap_w0
xfeed_8203 0 1 decap_w0
xfeed_8202 0 1 decap_w0
xfeed_8201 0 1 decap_w0
xfeed_7599 0 1 decap_w0
xfeed_7598 0 1 decap_w0
xfeed_7597 0 1 decap_w0
xfeed_7596 0 1 decap_w0
xfeed_7595 0 1 decap_w0
xfeed_7594 0 1 decap_w0
xfeed_7593 0 1 decap_w0
xfeed_7592 0 1 decap_w0
xfeed_7591 0 1 decap_w0
xfeed_7590 0 1 decap_w0
xfeed_3289 0 1 decap_w0
xfeed_3287 0 1 decap_w0
xfeed_3286 0 1 decap_w0
xfeed_3285 0 1 decap_w0
xfeed_3284 0 1 decap_w0
xfeed_3283 0 1 decap_w0
xfeed_3281 0 1 decap_w0
xfeed_3280 0 1 decap_w0
xfeed_2759 0 1 decap_w0
xfeed_2758 0 1 decap_w0
xfeed_2757 0 1 decap_w0
xfeed_2756 0 1 tie
xfeed_2755 0 1 decap_w0
xfeed_2754 0 1 decap_w0
xfeed_2753 0 1 decap_w0
xfeed_2752 0 1 tie
xfeed_2751 0 1 decap_w0
xfeed_2750 0 1 decap_w0
xfeed_730 0 1 decap_w0
xsubckt_468_and3_x1 0 1 282 285 284 283 and3_x1
xsubckt_1354_nand2_x0 0 1 1234 1241 1236 nand2_x0
xfeed_10109 0 1 decap_w0
xfeed_10108 0 1 decap_w0
xfeed_10107 0 1 decap_w0
xfeed_10106 0 1 decap_w0
xfeed_10105 0 1 decap_w0
xfeed_10104 0 1 decap_w0
xfeed_10103 0 1 decap_w0
xfeed_10102 0 1 decap_w0
xfeed_10101 0 1 decap_w0
xfeed_738 0 1 decap_w0
xfeed_737 0 1 decap_w0
xfeed_736 0 1 decap_w0
xfeed_735 0 1 decap_w0
xfeed_734 0 1 decap_w0
xfeed_733 0 1 tie
xfeed_732 0 1 decap_w0
xfeed_731 0 1 decap_w0
xsubckt_1230_and21nor_x0 0 1 1334 775 1352 1335 and21nor_x0
xsubckt_1174_nand2_x0 0 1 1388 1391 1390 nand2_x0
xsubckt_380_and3_x1 0 1 369 638 632 530 and3_x1
xsubckt_1770_or21nand_x0 0 1 824 831 829 827 or21nand_x0
xfeed_8219 0 1 decap_w0
xfeed_8218 0 1 tie
xfeed_8217 0 1 decap_w0
xfeed_8216 0 1 decap_w0
xfeed_8215 0 1 decap_w0
xfeed_8214 0 1 decap_w0
xfeed_8213 0 1 decap_w0
xfeed_8212 0 1 decap_w0
xfeed_8211 0 1 tie
xfeed_8210 0 1 decap_w0
xfeed_3299 0 1 decap_w0
xfeed_3298 0 1 decap_w0
xfeed_3297 0 1 decap_w0
xfeed_3296 0 1 decap_w0
xfeed_3295 0 1 decap_w0
xfeed_3294 0 1 tie
xfeed_3293 0 1 decap_w0
xfeed_3292 0 1 decap_w0
xfeed_3291 0 1 decap_w0
xfeed_3290 0 1 decap_w0
xfeed_2769 0 1 decap_w0
xfeed_2768 0 1 decap_w0
xfeed_2767 0 1 decap_w0
xfeed_2766 0 1 decap_w0
xfeed_2765 0 1 decap_w0
xfeed_2764 0 1 decap_w0
xfeed_2763 0 1 decap_w0
xfeed_2762 0 1 decap_w0
xfeed_2761 0 1 decap_w0
xfeed_2760 0 1 decap_w0
xsubckt_390_nand3_x0 0 1 359 660 651 646 nand3_x0
xfeed_10119 0 1 decap_w0
xfeed_10118 0 1 decap_w0
xfeed_10117 0 1 decap_w0
xfeed_10116 0 1 decap_w0
xfeed_10115 0 1 decap_w0
xfeed_10114 0 1 decap_w0
xfeed_10113 0 1 decap_w0
xfeed_10112 0 1 decap_w0
xfeed_10111 0 1 decap_w0
xfeed_10110 0 1 decap_w0
xfeed_749 0 1 decap_w0
xfeed_748 0 1 decap_w0
xfeed_747 0 1 decap_w0
xfeed_746 0 1 decap_w0
xfeed_745 0 1 tie
xfeed_744 0 1 decap_w0
xfeed_743 0 1 decap_w0
xfeed_742 0 1 decap_w0
xfeed_741 0 1 decap_w0
xfeed_740 0 1 decap_w0
xsubckt_1330_and21nor_x0 0 1 1256 1257 1266 1273 and21nor_x0
xfeed_8229 0 1 decap_w0
xfeed_8228 0 1 decap_w0
xfeed_8227 0 1 decap_w0
xfeed_8226 0 1 decap_w0
xfeed_8225 0 1 decap_w0
xfeed_8224 0 1 decap_w0
xfeed_8223 0 1 decap_w0
xfeed_8222 0 1 tie
xfeed_8221 0 1 decap_w0
xfeed_8220 0 1 decap_w0
xfeed_2779 0 1 decap_w0
xfeed_2778 0 1 decap_w0
xfeed_2777 0 1 decap_w0
xfeed_2776 0 1 decap_w0
xfeed_2775 0 1 decap_w0
xfeed_2774 0 1 decap_w0
xfeed_2773 0 1 decap_w0
xfeed_2772 0 1 decap_w0
xfeed_2771 0 1 decap_w0
xfeed_2770 0 1 decap_w0
xsubckt_1126_and21nor_x0 0 1 1431 1432 1436 1437 and21nor_x0
xsubckt_846_or2_x1 0 1 2100 1639 1633 or2_x1
xsubckt_1527_and21nor_x0 0 1 1066 1069 1073 1094 and21nor_x0
xsubckt_1666_or21nand_x0 0 1 928 931 1122 141 or21nand_x0
xfeed_13909 0 1 tie
xfeed_13908 0 1 tie
xfeed_13907 0 1 tie
xfeed_13905 0 1 tie
xfeed_13904 0 1 tie
xfeed_13902 0 1 tie
xfeed_10129 0 1 decap_w0
xfeed_10128 0 1 decap_w0
xfeed_10127 0 1 decap_w0
xfeed_10126 0 1 decap_w0
xfeed_10125 0 1 decap_w0
xfeed_10124 0 1 decap_w0
xfeed_10123 0 1 decap_w0
xfeed_10122 0 1 decap_w0
xfeed_10121 0 1 decap_w0
xfeed_10120 0 1 decap_w0
xfeed_759 0 1 decap_w0
xfeed_758 0 1 decap_w0
xfeed_757 0 1 decap_w0
xfeed_756 0 1 decap_w0
xfeed_755 0 1 decap_w0
xfeed_754 0 1 decap_w0
xfeed_753 0 1 decap_w0
xfeed_752 0 1 tie
xfeed_751 0 1 decap_w0
xfeed_750 0 1 decap_w0
xsubckt_1265_or21nand_x0 0 1 1315 1982 479 1316 or21nand_x0
xsubckt_1053_and3_x1 0 1 1488 653 623 519 and3_x1
xsubckt_20_inv_x0 0 1 762 2048 inv_x0
xsubckt_1410_and3_x1 0 1 1182 1207 1196 1184 and3_x1
xfeed_8239 0 1 decap_w0
xfeed_8238 0 1 decap_w0
xfeed_8237 0 1 decap_w0
xfeed_8235 0 1 decap_w0
xfeed_8234 0 1 decap_w0
xfeed_8233 0 1 decap_w0
xfeed_8232 0 1 decap_w0
xfeed_8231 0 1 decap_w0
xfeed_8230 0 1 decap_w0
xfeed_7709 0 1 decap_w0
xfeed_7708 0 1 decap_w0
xfeed_7707 0 1 decap_w0
xfeed_7706 0 1 decap_w0
xfeed_7705 0 1 decap_w0
xfeed_7704 0 1 decap_w0
xfeed_7703 0 1 decap_w0
xfeed_7702 0 1 decap_w0
xfeed_7701 0 1 decap_w0
xfeed_7700 0 1 decap_w0
xfeed_2788 0 1 decap_w0
xfeed_2787 0 1 decap_w0
xfeed_2786 0 1 decap_w0
xfeed_2785 0 1 decap_w0
xfeed_2784 0 1 decap_w0
xfeed_2782 0 1 tie
xfeed_2781 0 1 decap_w0
xfeed_2780 0 1 decap_w0
xsubckt_1063_nand3_x0 0 1 1479 643 313 1554 nand3_x0
xsubckt_22_inv_x0 0 1 760 2047 inv_x0
xsubckt_24_inv_x0 0 1 758 1957 inv_x0
xsubckt_26_inv_x0 0 1 756 1947 inv_x0
xsubckt_1339_nor2_x0 0 1 1248 1252 1249 nor2_x0
xfeed_13919 0 1 tie
xfeed_13915 0 1 tie
xfeed_13913 0 1 tie
xfeed_13912 0 1 tie
xfeed_13911 0 1 tie
xfeed_13910 0 1 tie
xfeed_10139 0 1 decap_w0
xfeed_10138 0 1 decap_w0
xfeed_10137 0 1 decap_w0
xfeed_10136 0 1 decap_w0
xfeed_10135 0 1 decap_w0
xfeed_10134 0 1 decap_w0
xfeed_10133 0 1 decap_w0
xfeed_10132 0 1 tie
xfeed_10131 0 1 decap_w0
xfeed_10130 0 1 decap_w0
xfeed_769 0 1 decap_w0
xfeed_768 0 1 decap_w0
xfeed_767 0 1 decap_w0
xfeed_766 0 1 decap_w0
xfeed_765 0 1 decap_w0
xfeed_763 0 1 decap_w0
xfeed_762 0 1 decap_w0
xfeed_761 0 1 decap_w0
xfeed_760 0 1 decap_w0
xsubckt_861_and21nor_x0 0 1 1620 775 1623 1621 and21nor_x0
xsubckt_289_nand3_x0 0 1 459 1929 715 599 nand3_x0
xsubckt_188_and3_x1 0 1 570 1925 711 571 and3_x1
xsubckt_28_inv_x0 0 1 754 1981 inv_x0
xsubckt_523_and4_x1 0 1 229 448 444 317 316 and4_x1
xsubckt_1646_mux2_x1 0 1 948 991 950 1142 mux2_x1
xfeed_8249 0 1 decap_w0
xfeed_8248 0 1 decap_w0
xfeed_8247 0 1 decap_w0
xfeed_8246 0 1 decap_w0
xfeed_8245 0 1 decap_w0
xfeed_8244 0 1 decap_w0
xfeed_8243 0 1 decap_w0
xfeed_8242 0 1 decap_w0
xfeed_8241 0 1 decap_w0
xfeed_8240 0 1 decap_w0
xfeed_7719 0 1 decap_w0
xfeed_7718 0 1 decap_w0
xfeed_7717 0 1 decap_w0
xfeed_7716 0 1 decap_w0
xfeed_7715 0 1 tie
xfeed_7714 0 1 decap_w0
xfeed_7713 0 1 decap_w0
xfeed_7712 0 1 decap_w0
xfeed_7711 0 1 tie
xfeed_7710 0 1 decap_w0
xfeed_3409 0 1 decap_w0
xfeed_3408 0 1 decap_w0
xfeed_3407 0 1 decap_w0
xfeed_3406 0 1 decap_w0
xfeed_3405 0 1 decap_w0
xfeed_3404 0 1 decap_w0
xfeed_3403 0 1 decap_w0
xfeed_3402 0 1 decap_w0
xfeed_3401 0 1 decap_w0
xfeed_3400 0 1 decap_w0
xfeed_2799 0 1 decap_w0
xfeed_2798 0 1 decap_w0
xfeed_2797 0 1 decap_w0
xfeed_2796 0 1 tie
xfeed_2795 0 1 decap_w0
xfeed_2794 0 1 decap_w0
xfeed_2793 0 1 decap_w0
xfeed_2792 0 1 decap_w0
xfeed_2791 0 1 decap_w0
xfeed_2790 0 1 decap_w0
xsubckt_1119_mux2_x1 0 1 1838 1996 1987 1438 mux2_x1
xsubckt_431_and4_x1 0 1 318 469 431 332 320 and4_x1
xsubckt_1630_and21nor_x0 0 1 964 965 1121 128 and21nor_x0
xfeed_13929 0 1 tie
xfeed_13928 0 1 tie
xfeed_13927 0 1 tie
xfeed_13925 0 1 tie
xfeed_13924 0 1 tie
xfeed_13923 0 1 tie
xfeed_13921 0 1 tie
xfeed_13920 0 1 tie
xfeed_10149 0 1 tie
xfeed_10148 0 1 decap_w0
xfeed_10147 0 1 decap_w0
xfeed_10146 0 1 decap_w0
xfeed_10145 0 1 decap_w0
xfeed_10144 0 1 decap_w0
xfeed_10143 0 1 decap_w0
xfeed_10142 0 1 decap_w0
xfeed_10141 0 1 decap_w0
xfeed_10140 0 1 decap_w0
xfeed_779 0 1 decap_w0
xfeed_778 0 1 decap_w0
xfeed_776 0 1 decap_w0
xfeed_775 0 1 decap_w0
xfeed_774 0 1 decap_w0
xfeed_773 0 1 decap_w0
xfeed_772 0 1 decap_w0
xfeed_771 0 1 decap_w0
xfeed_770 0 1 decap_w0
xfeed_8259 0 1 decap_w0
xfeed_8257 0 1 decap_w0
xfeed_8256 0 1 decap_w0
xfeed_8255 0 1 decap_w0
xfeed_8254 0 1 decap_w0
xfeed_8253 0 1 decap_w0
xfeed_8252 0 1 decap_w0
xfeed_8251 0 1 decap_w0
xfeed_8250 0 1 decap_w0
xfeed_7729 0 1 decap_w0
xfeed_7728 0 1 decap_w0
xfeed_7727 0 1 decap_w0
xfeed_7726 0 1 decap_w0
xfeed_7725 0 1 decap_w0
xfeed_7724 0 1 decap_w0
xfeed_7723 0 1 decap_w0
xfeed_7722 0 1 tie
xfeed_7721 0 1 decap_w0
xfeed_7720 0 1 decap_w0
xfeed_3419 0 1 decap_w0
xfeed_3418 0 1 decap_w0
xfeed_3417 0 1 decap_w0
xfeed_3416 0 1 decap_w0
xfeed_3415 0 1 decap_w0
xfeed_3414 0 1 decap_w0
xfeed_3413 0 1 decap_w0
xfeed_3412 0 1 tie
xfeed_3411 0 1 decap_w0
xfeed_3410 0 1 decap_w0
xfeed_13939 0 1 tie
xfeed_13938 0 1 tie
xfeed_13937 0 1 tie
xfeed_13936 0 1 tie
xfeed_13935 0 1 tie
xfeed_13934 0 1 tie
xfeed_13933 0 1 tie
xfeed_13932 0 1 tie
xfeed_13931 0 1 tie
xfeed_13930 0 1 tie
xfeed_10159 0 1 decap_w0
xfeed_10158 0 1 tie
xfeed_10157 0 1 decap_w0
xfeed_10156 0 1 decap_w0
xfeed_10155 0 1 decap_w0
xfeed_10154 0 1 decap_w0
xfeed_10153 0 1 decap_w0
xfeed_10152 0 1 decap_w0
xfeed_10151 0 1 decap_w0
xfeed_10150 0 1 decap_w0
xfeed_789 0 1 decap_w0
xfeed_788 0 1 tie
xfeed_787 0 1 decap_w0
xfeed_786 0 1 decap_w0
xfeed_785 0 1 decap_w0
xfeed_784 0 1 decap_w0
xfeed_783 0 1 tie
xfeed_782 0 1 decap_w0
xfeed_781 0 1 decap_w0
xfeed_780 0 1 decap_w0
xsubckt_810_and3_x1 0 1 1664 2071 680 490 and3_x1
xsubckt_1305_nand3_x0 0 1 1279 2061 666 657 nand3_x0
xfeed_8269 0 1 decap_w0
xfeed_8268 0 1 decap_w0
xfeed_8267 0 1 decap_w0
xfeed_8266 0 1 decap_w0
xfeed_8265 0 1 tie
xfeed_8264 0 1 decap_w0
xfeed_8263 0 1 decap_w0
xfeed_8262 0 1 decap_w0
xfeed_8261 0 1 decap_w0
xfeed_8260 0 1 decap_w0
xfeed_7739 0 1 decap_w0
xfeed_7738 0 1 decap_w0
xfeed_7737 0 1 tie
xfeed_7736 0 1 decap_w0
xfeed_7735 0 1 decap_w0
xfeed_7734 0 1 decap_w0
xfeed_7732 0 1 decap_w0
xfeed_7731 0 1 decap_w0
xfeed_7730 0 1 decap_w0
xfeed_3429 0 1 decap_w0
xfeed_3428 0 1 decap_w0
xfeed_3427 0 1 tie
xfeed_3426 0 1 decap_w0
xfeed_3425 0 1 decap_w0
xfeed_3424 0 1 decap_w0
xfeed_3423 0 1 decap_w0
xfeed_3422 0 1 decap_w0
xfeed_3421 0 1 decap_w0
xfeed_3420 0 1 decap_w0
xsubckt_1218_and3_x1 0 1 1346 1350 1349 1347 and3_x1
xsubckt_651_nor2_x0 0 1 108 763 109 nor2_x0
xsubckt_1940_dff_x1 0 1 1970 1808 38 dff_x1
xfeed_13949 0 1 tie
xfeed_13948 0 1 tie
xfeed_13947 0 1 tie
xfeed_13946 0 1 tie
xfeed_13945 0 1 tie
xfeed_13944 0 1 tie
xfeed_13943 0 1 tie
xfeed_13942 0 1 tie
xfeed_13941 0 1 tie
xfeed_13940 0 1 tie
xfeed_10169 0 1 decap_w0
xfeed_10168 0 1 decap_w0
xfeed_10167 0 1 decap_w0
xfeed_10166 0 1 decap_w0
xfeed_10164 0 1 decap_w0
xfeed_10163 0 1 decap_w0
xfeed_10162 0 1 decap_w0
xfeed_10161 0 1 decap_w0
xfeed_10160 0 1 decap_w0
xfeed_799 0 1 decap_w0
xfeed_798 0 1 decap_w0
xfeed_797 0 1 decap_w0
xfeed_796 0 1 decap_w0
xfeed_795 0 1 decap_w0
xfeed_794 0 1 decap_w0
xfeed_793 0 1 decap_w0
xfeed_792 0 1 decap_w0
xfeed_791 0 1 decap_w0
xfeed_790 0 1 decap_w0
xsubckt_1264_or21nand_x0 0 1 1316 1330 1321 1318 or21nand_x0
xsubckt_595_or21nand_x0 0 1 160 1982 450 411 or21nand_x0
xsubckt_1815_mux2_x1 0 1 1790 2047 798 773 mux2_x1
xsubckt_1942_dff_x1 0 1 1968 1806 38 dff_x1
xsubckt_1944_dff_x1 0 1 1980 1804 38 dff_x1
xsubckt_1946_dff_x1 0 1 1978 1802 58 dff_x1
xfeed_8279 0 1 tie
xfeed_8278 0 1 decap_w0
xfeed_8277 0 1 decap_w0
xfeed_8276 0 1 decap_w0
xfeed_8275 0 1 decap_w0
xfeed_8274 0 1 decap_w0
xfeed_8273 0 1 decap_w0
xfeed_8272 0 1 tie
xfeed_8271 0 1 decap_w0
xfeed_8270 0 1 decap_w0
xfeed_7749 0 1 decap_w0
xfeed_7748 0 1 decap_w0
xfeed_7747 0 1 decap_w0
xfeed_7746 0 1 decap_w0
xfeed_7745 0 1 decap_w0
xfeed_7744 0 1 decap_w0
xfeed_7743 0 1 decap_w0
xfeed_7742 0 1 tie
xfeed_7741 0 1 decap_w0
xfeed_7740 0 1 decap_w0
xfeed_3439 0 1 tie
xfeed_3438 0 1 decap_w0
xfeed_3437 0 1 decap_w0
xfeed_3436 0 1 decap_w0
xfeed_3435 0 1 decap_w0
xfeed_3434 0 1 tie
xfeed_3433 0 1 decap_w0
xfeed_3432 0 1 decap_w0
xfeed_3431 0 1 decap_w0
xfeed_3430 0 1 decap_w0
xfeed_2909 0 1 decap_w0
xfeed_2908 0 1 decap_w0
xfeed_2907 0 1 decap_w0
xfeed_2906 0 1 decap_w0
xfeed_2905 0 1 decap_w0
xfeed_2904 0 1 decap_w0
xfeed_2903 0 1 decap_w0
xfeed_2902 0 1 decap_w0
xfeed_2901 0 1 decap_w0
xfeed_2900 0 1 decap_w0
xsubckt_714_and3_x1 0 1 1750 1755 1754 1751 and3_x1
xsubckt_305_and2_x1 0 1 443 448 444 and2_x1
xsubckt_1948_dff_x1 0 1 1976 1800 58 dff_x1
xfeed_13959 0 1 tie
xfeed_13958 0 1 tie
xfeed_13957 0 1 tie
xfeed_13955 0 1 tie
xfeed_13954 0 1 tie
xfeed_13953 0 1 tie
xfeed_13952 0 1 tie
xfeed_13951 0 1 tie
xfeed_13950 0 1 tie
xfeed_10179 0 1 decap_w0
xfeed_10178 0 1 decap_w0
xfeed_10177 0 1 decap_w0
xfeed_10176 0 1 decap_w0
xfeed_10175 0 1 decap_w0
xfeed_10174 0 1 decap_w0
xfeed_10173 0 1 decap_w0
xfeed_10172 0 1 decap_w0
xfeed_10171 0 1 decap_w0
xfeed_10170 0 1 decap_w0
xsubckt_787_or3_x1 0 1 1684 1689 1688 1685 or3_x1
xsubckt_441_nor3_x0 0 1 309 428 331 311 nor3_x0
xfeed_8289 0 1 tie
xfeed_8288 0 1 decap_w0
xfeed_8287 0 1 decap_w0
xfeed_8286 0 1 decap_w0
xfeed_8285 0 1 decap_w0
xfeed_8284 0 1 decap_w0
xfeed_8283 0 1 decap_w0
xfeed_8282 0 1 decap_w0
xfeed_8281 0 1 decap_w0
xfeed_8280 0 1 decap_w0
xfeed_7759 0 1 decap_w0
xfeed_7758 0 1 tie
xfeed_7757 0 1 decap_w0
xfeed_7756 0 1 decap_w0
xfeed_7755 0 1 decap_w0
xfeed_7754 0 1 tie
xfeed_7753 0 1 decap_w0
xfeed_7752 0 1 decap_w0
xfeed_7751 0 1 decap_w0
xfeed_7750 0 1 decap_w0
xfeed_3449 0 1 tie
xfeed_3448 0 1 decap_w0
xfeed_3447 0 1 decap_w0
xfeed_3446 0 1 decap_w0
xfeed_3445 0 1 decap_w0
xfeed_3444 0 1 decap_w0
xfeed_3443 0 1 decap_w0
xfeed_3442 0 1 decap_w0
xfeed_3441 0 1 decap_w0
xfeed_2919 0 1 decap_w0
xfeed_2918 0 1 decap_w0
xfeed_2917 0 1 decap_w0
xfeed_2916 0 1 decap_w0
xfeed_2915 0 1 decap_w0
xfeed_2914 0 1 decap_w0
xfeed_2913 0 1 decap_w0
xfeed_2912 0 1 decap_w0
xfeed_2911 0 1 decap_w0
xfeed_2910 0 1 decap_w0
xsubckt_955_nand2_x0 0 1 1565 383 1567 nand2_x0
xsubckt_1325_and21nor_x0 0 1 1261 749 478 1317 and21nor_x0
xsubckt_1726_and21nor_x0 0 1 868 1104 873 871 and21nor_x0
xfeed_13969 0 1 tie
xfeed_13967 0 1 tie
xfeed_13966 0 1 tie
xfeed_13965 0 1 tie
xfeed_13964 0 1 tie
xfeed_13963 0 1 tie
xfeed_13962 0 1 tie
xfeed_13961 0 1 tie
xfeed_13960 0 1 tie
xfeed_10189 0 1 decap_w0
xfeed_10188 0 1 decap_w0
xfeed_10187 0 1 decap_w0
xfeed_10186 0 1 decap_w0
xfeed_10185 0 1 decap_w0
xfeed_10184 0 1 tie
xfeed_10183 0 1 decap_w0
xfeed_10182 0 1 decap_w0
xfeed_10181 0 1 decap_w0
xfeed_10180 0 1 decap_w0
xfeed_8299 0 1 decap_w0
xfeed_8298 0 1 decap_w0
xfeed_8297 0 1 decap_w0
xfeed_8296 0 1 decap_w0
xfeed_8295 0 1 decap_w0
xfeed_8294 0 1 decap_w0
xfeed_8293 0 1 decap_w0
xfeed_8292 0 1 decap_w0
xfeed_8291 0 1 decap_w0
xfeed_8290 0 1 decap_w0
xfeed_7769 0 1 decap_w0
xfeed_7768 0 1 tie
xfeed_7767 0 1 decap_w0
xfeed_7766 0 1 decap_w0
xfeed_7765 0 1 decap_w0
xfeed_7764 0 1 decap_w0
xfeed_7763 0 1 decap_w0
xfeed_7762 0 1 decap_w0
xfeed_7761 0 1 decap_w0
xfeed_7760 0 1 decap_w0
xfeed_3459 0 1 decap_w0
xfeed_3458 0 1 decap_w0
xfeed_3457 0 1 decap_w0
xfeed_3456 0 1 decap_w0
xfeed_3455 0 1 decap_w0
xfeed_3454 0 1 decap_w0
xfeed_3453 0 1 decap_w0
xfeed_3452 0 1 decap_w0
xfeed_3451 0 1 decap_w0
xfeed_3450 0 1 decap_w0
xfeed_2929 0 1 decap_w0
xfeed_2928 0 1 decap_w0
xfeed_2927 0 1 decap_w0
xfeed_2926 0 1 decap_w0
xfeed_2925 0 1 decap_w0
xfeed_2924 0 1 decap_w0
xfeed_2923 0 1 decap_w0
xfeed_2922 0 1 decap_w0
xfeed_2921 0 1 decap_w0
xfeed_2920 0 1 decap_w0
xsubckt_1351_and4_x1 0 1 1237 435 1682 1239 1238 and4_x1
xsubckt_1579_and2_x1 0 1 1015 1018 1016 and2_x1
xfeed_13978 0 1 tie
xfeed_13977 0 1 tie
xfeed_13976 0 1 tie
xfeed_13974 0 1 tie
xfeed_13973 0 1 tie
xfeed_13972 0 1 tie
xfeed_13971 0 1 tie
xfeed_13970 0 1 tie
xfeed_10199 0 1 decap_w0
xfeed_10198 0 1 decap_w0
xfeed_10197 0 1 decap_w0
xfeed_10196 0 1 decap_w0
xfeed_10195 0 1 decap_w0
xfeed_10194 0 1 decap_w0
xfeed_10193 0 1 decap_w0
xfeed_10192 0 1 decap_w0
xfeed_10191 0 1 tie
xfeed_10190 0 1 decap_w0
xfeed_909 0 1 decap_w0
xfeed_908 0 1 decap_w0
xfeed_907 0 1 decap_w0
xfeed_906 0 1 tie
xfeed_905 0 1 decap_w0
xfeed_904 0 1 decap_w0
xfeed_903 0 1 decap_w0
xfeed_902 0 1 decap_w0
xfeed_901 0 1 decap_w0
xfeed_900 0 1 decap_w0
xsubckt_1275_nand3_x0 0 1 1306 784 679 447 nand3_x0
xsubckt_1178_mux2_x1 0 1 1384 2053 781 1940 mux2_x1
xsubckt_195_and2_x1 0 1 563 573 565 and2_x1
xfeed_7779 0 1 decap_w0
xfeed_7778 0 1 decap_w0
xfeed_7777 0 1 decap_w0
xfeed_7776 0 1 decap_w0
xfeed_7775 0 1 decap_w0
xfeed_7774 0 1 decap_w0
xfeed_7773 0 1 decap_w0
xfeed_7772 0 1 decap_w0
xfeed_7771 0 1 decap_w0
xfeed_7770 0 1 decap_w0
xfeed_3469 0 1 decap_w0
xfeed_3468 0 1 tie
xfeed_3467 0 1 decap_w0
xfeed_3466 0 1 decap_w0
xfeed_3465 0 1 decap_w0
xfeed_3464 0 1 decap_w0
xfeed_3463 0 1 decap_w0
xfeed_3462 0 1 decap_w0
xfeed_3461 0 1 decap_w0
xfeed_3460 0 1 decap_w0
xfeed_2939 0 1 decap_w0
xfeed_2938 0 1 decap_w0
xfeed_2937 0 1 decap_w0
xfeed_2936 0 1 decap_w0
xfeed_2935 0 1 decap_w0
xfeed_2934 0 1 decap_w0
xfeed_2933 0 1 decap_w0
xfeed_2932 0 1 decap_w0
xfeed_2931 0 1 decap_w0
xfeed_2930 0 1 decap_w0
xfeed_13985 0 1 tie
xfeed_13984 0 1 tie
xfeed_13983 0 1 tie
xfeed_13981 0 1 tie
xfeed_13980 0 1 tie
xfeed_919 0 1 decap_w0
xfeed_918 0 1 tie
xfeed_917 0 1 decap_w0
xfeed_916 0 1 decap_w0
xfeed_915 0 1 decap_w0
xfeed_914 0 1 decap_w0
xfeed_913 0 1 tie
xfeed_912 0 1 decap_w0
xfeed_911 0 1 decap_w0
xfeed_910 0 1 decap_w0
xsubckt_1369_and3_x1 0 1 1220 1245 1234 1222 and3_x1
xsubckt_1664_or21nand_x0 0 1 930 933 1118 765 or21nand_x0
xfeed_13989 0 1 tie
xfeed_13988 0 1 tie
xfeed_13987 0 1 tie
xfeed_13986 0 1 tie
xfeed_7789 0 1 decap_w0
xfeed_7788 0 1 decap_w0
xfeed_7787 0 1 tie
xfeed_7786 0 1 decap_w0
xfeed_7785 0 1 decap_w0
xfeed_7784 0 1 decap_w0
xfeed_7783 0 1 decap_w0
xfeed_7782 0 1 decap_w0
xfeed_7781 0 1 decap_w0
xfeed_7780 0 1 decap_w0
xfeed_3479 0 1 decap_w0
xfeed_3478 0 1 decap_w0
xfeed_3477 0 1 decap_w0
xfeed_3476 0 1 decap_w0
xfeed_3475 0 1 tie
xfeed_3474 0 1 decap_w0
xfeed_3473 0 1 decap_w0
xfeed_3472 0 1 decap_w0
xfeed_3471 0 1 decap_w0
xfeed_3470 0 1 decap_w0
xfeed_2949 0 1 decap_w0
xfeed_2947 0 1 decap_w0
xfeed_2946 0 1 decap_w0
xfeed_2945 0 1 decap_w0
xfeed_2944 0 1 decap_w0
xfeed_2943 0 1 decap_w0
xfeed_2942 0 1 decap_w0
xfeed_2941 0 1 decap_w0
xfeed_2940 0 1 decap_w0
xsubckt_1317_and2_x1 0 1 1268 435 1269 and2_x1
xsubckt_1358_nand2_x0 0 1 1806 1242 1231 nand2_x0
xfeed_13992 0 1 tie
xfeed_13991 0 1 tie
xfeed_929 0 1 decap_w0
xfeed_928 0 1 decap_w0
xfeed_927 0 1 decap_w0
xfeed_926 0 1 decap_w0
xfeed_925 0 1 decap_w0
xfeed_924 0 1 decap_w0
xfeed_923 0 1 decap_w0
xfeed_922 0 1 decap_w0
xfeed_921 0 1 decap_w0
xfeed_920 0 1 decap_w0
xsubckt_1224_and21nor_x0 0 1 1340 499 495 609 and21nor_x0
xsubckt_306_nand3_x0 0 1 442 609 557 451 nand3_x0
xsubckt_1521_nand2_x0 0 1 1075 1082 1078 nand2_x0
xsubckt_1567_nor2_x0 0 1 1027 100 1122 nor2_x0
xfeed_13999 0 1 tie
xfeed_13998 0 1 tie
xfeed_13997 0 1 tie
xfeed_13996 0 1 tie
xfeed_13995 0 1 tie
xfeed_13994 0 1 tie
xfeed_13993 0 1 tie
xfeed_8409 0 1 decap_w0
xfeed_8408 0 1 decap_w0
xfeed_8407 0 1 decap_w0
xfeed_8406 0 1 decap_w0
xfeed_8405 0 1 decap_w0
xfeed_8404 0 1 tie
xfeed_8403 0 1 decap_w0
xfeed_8402 0 1 decap_w0
xfeed_8401 0 1 decap_w0
xfeed_8400 0 1 decap_w0
xfeed_7798 0 1 decap_w0
xfeed_7797 0 1 decap_w0
xfeed_7796 0 1 tie
xfeed_7795 0 1 decap_w0
xfeed_7794 0 1 decap_w0
xfeed_7793 0 1 decap_w0
xfeed_7792 0 1 decap_w0
xfeed_7791 0 1 decap_w0
xfeed_7790 0 1 decap_w0
xfeed_3489 0 1 decap_w0
xfeed_3488 0 1 decap_w0
xfeed_3487 0 1 decap_w0
xfeed_3486 0 1 decap_w0
xfeed_3485 0 1 decap_w0
xfeed_3484 0 1 decap_w0
xfeed_3483 0 1 decap_w0
xfeed_3482 0 1 decap_w0
xfeed_3481 0 1 decap_w0
xfeed_3480 0 1 decap_w0
xfeed_2959 0 1 tie
xfeed_2958 0 1 decap_w0
xfeed_2957 0 1 decap_w0
xfeed_2956 0 1 decap_w0
xfeed_2955 0 1 decap_w0
xfeed_2954 0 1 decap_w0
xfeed_2953 0 1 decap_w0
xfeed_2952 0 1 decap_w0
xfeed_2951 0 1 decap_w0
xfeed_2950 0 1 decap_w0
xsubckt_1695_nand3_x0 0 1 899 1981 679 595 nand3_x0
xfeed_10309 0 1 decap_w0
xfeed_10308 0 1 decap_w0
xfeed_10307 0 1 decap_w0
xfeed_10305 0 1 decap_w0
xfeed_10304 0 1 decap_w0
xfeed_10303 0 1 decap_w0
xfeed_10302 0 1 decap_w0
xfeed_10301 0 1 tie
xfeed_10300 0 1 decap_w0
xfeed_939 0 1 decap_w0
xfeed_938 0 1 decap_w0
xfeed_937 0 1 decap_w0
xfeed_936 0 1 decap_w0
xfeed_935 0 1 decap_w0
xfeed_934 0 1 decap_w0
xfeed_933 0 1 decap_w0
xfeed_932 0 1 decap_w0
xfeed_930 0 1 tie
xsubckt_1071_and4_x1 0 1 1472 652 532 526 1563 and4_x1
xsubckt_935_mux2_x1 0 1 1882 2022 1581 1578 mux2_x1
xsubckt_773_and3_x1 0 1 1697 1970 1749 1739 and3_x1
xfeed_8419 0 1 decap_w0
xfeed_8418 0 1 decap_w0
xfeed_8417 0 1 decap_w0
xfeed_8416 0 1 decap_w0
xfeed_8415 0 1 decap_w0
xfeed_8414 0 1 decap_w0
xfeed_8413 0 1 decap_w0
xfeed_8412 0 1 decap_w0
xfeed_8411 0 1 decap_w0
xfeed_8410 0 1 decap_w0
xfeed_4109 0 1 decap_w0
xfeed_4108 0 1 decap_w0
xfeed_4106 0 1 tie
xfeed_4105 0 1 decap_w0
xfeed_4104 0 1 decap_w0
xfeed_4103 0 1 decap_w0
xfeed_4102 0 1 decap_w0
xfeed_4101 0 1 decap_w0
xfeed_4100 0 1 decap_w0
xfeed_3499 0 1 decap_w0
xfeed_3498 0 1 decap_w0
xfeed_3497 0 1 decap_w0
xfeed_3496 0 1 decap_w0
xfeed_3495 0 1 decap_w0
xfeed_3494 0 1 decap_w0
xfeed_3493 0 1 decap_w0
xfeed_3492 0 1 decap_w0
xfeed_3491 0 1 decap_w0
xfeed_3490 0 1 decap_w0
xfeed_2969 0 1 decap_w0
xfeed_2968 0 1 decap_w0
xfeed_2967 0 1 decap_w0
xfeed_2966 0 1 decap_w0
xfeed_2965 0 1 decap_w0
xfeed_2964 0 1 decap_w0
xfeed_2963 0 1 decap_w0
xfeed_2962 0 1 decap_w0
xfeed_2961 0 1 decap_w0
xfeed_2960 0 1 decap_w0
xsubckt_809_and2_x1 0 1 1665 2051 1740 and2_x1
xsubckt_721_and2_x1 0 1 1743 600 1745 and2_x1
xsubckt_567_nand2_x0 0 1 188 663 191 nand2_x0
xsubckt_1704_mux2_x1 0 1 890 895 891 901 mux2_x1
xfeed_10319 0 1 decap_w0
xfeed_10318 0 1 decap_w0
xfeed_10317 0 1 decap_w0
xfeed_10316 0 1 decap_w0
xfeed_10315 0 1 decap_w0
xfeed_10314 0 1 decap_w0
xfeed_10313 0 1 decap_w0
xfeed_10312 0 1 decap_w0
xfeed_10311 0 1 tie
xfeed_10310 0 1 decap_w0
xfeed_949 0 1 decap_w0
xfeed_948 0 1 decap_w0
xfeed_947 0 1 decap_w0
xfeed_946 0 1 decap_w0
xfeed_945 0 1 decap_w0
xfeed_944 0 1 decap_w0
xfeed_943 0 1 decap_w0
xfeed_942 0 1 decap_w0
xfeed_941 0 1 decap_w0
xfeed_940 0 1 tie
xsubckt_1094_or3_x1 0 1 1453 642 312 1454 or3_x1
xsubckt_1067_and4_x1 0 1 1476 661 651 529 528 and4_x1
xsubckt_730_nand2_x0 0 1 1734 1736 1735 nand2_x0
xsubckt_1424_and4_x1 0 1 1169 1207 1196 1184 1171 and4_x1
xsubckt_1564_and2_x1 0 1 1030 1033 1031 and2_x1
xfeed_8429 0 1 decap_w0
xfeed_8428 0 1 decap_w0
xfeed_8427 0 1 decap_w0
xfeed_8426 0 1 decap_w0
xfeed_8425 0 1 decap_w0
xfeed_8424 0 1 decap_w0
xfeed_8423 0 1 decap_w0
xfeed_8422 0 1 decap_w0
xfeed_8421 0 1 tie
xfeed_8420 0 1 decap_w0
xfeed_4119 0 1 decap_w0
xfeed_4118 0 1 tie
xfeed_4116 0 1 decap_w0
xfeed_4115 0 1 decap_w0
xfeed_4114 0 1 decap_w0
xfeed_4113 0 1 tie
xfeed_4112 0 1 decap_w0
xfeed_4111 0 1 decap_w0
xfeed_4110 0 1 decap_w0
xfeed_2979 0 1 decap_w0
xfeed_2978 0 1 decap_w0
xfeed_2977 0 1 decap_w0
xfeed_2976 0 1 decap_w0
xfeed_2974 0 1 tie
xfeed_2973 0 1 decap_w0
xfeed_2972 0 1 decap_w0
xfeed_2971 0 1 decap_w0
xfeed_2970 0 1 decap_w0
xsubckt_31_inv_x0 0 1 751 1972 inv_x0
xsubckt_33_inv_x0 0 1 749 1970 inv_x0
xsubckt_119_nand2_x0 0 1 649 660 651 nand2_x0
xsubckt_640_nand2_x0 0 1 119 121 120 nand2_x0
xsubckt_1498_and4_x1 0 1 1098 1380 1354 1348 1339 and4_x1
xfeed_10329 0 1 decap_w0
xfeed_10328 0 1 decap_w0
xfeed_10327 0 1 decap_w0
xfeed_10326 0 1 decap_w0
xfeed_10325 0 1 decap_w0
xfeed_10324 0 1 decap_w0
xfeed_10323 0 1 decap_w0
xfeed_10322 0 1 decap_w0
xfeed_10321 0 1 decap_w0
xfeed_10320 0 1 decap_w0
xfeed_959 0 1 decap_w0
xfeed_958 0 1 decap_w0
xfeed_957 0 1 decap_w0
xfeed_955 0 1 decap_w0
xfeed_954 0 1 decap_w0
xfeed_953 0 1 decap_w0
xfeed_952 0 1 decap_w0
xfeed_951 0 1 decap_w0
xfeed_950 0 1 decap_w0
xsubckt_994_or21nand_x0 0 1 1534 1576 1541 1535 or21nand_x0
xsubckt_677_and3_x1 0 1 1785 89 88 85 and3_x1
xsubckt_268_and2_x1 0 1 480 483 481 and2_x1
xsubckt_35_inv_x0 0 1 747 2073 inv_x0
xsubckt_37_inv_x0 0 1 745 2071 inv_x0
xsubckt_39_inv_x0 0 1 743 2069 inv_x0
xfeed_8439 0 1 decap_w0
xfeed_8438 0 1 decap_w0
xfeed_8437 0 1 decap_w0
xfeed_8436 0 1 decap_w0
xfeed_8435 0 1 decap_w0
xfeed_8434 0 1 decap_w0
xfeed_8433 0 1 decap_w0
xfeed_8432 0 1 decap_w0
xfeed_8431 0 1 decap_w0
xfeed_8430 0 1 decap_w0
xfeed_7909 0 1 decap_w0
xfeed_7908 0 1 decap_w0
xfeed_7907 0 1 decap_w0
xfeed_7906 0 1 decap_w0
xfeed_7905 0 1 decap_w0
xfeed_7904 0 1 decap_w0
xfeed_7903 0 1 decap_w0
xfeed_7902 0 1 decap_w0
xfeed_7901 0 1 decap_w0
xfeed_7900 0 1 decap_w0
xfeed_4129 0 1 decap_w0
xfeed_4128 0 1 decap_w0
xfeed_4127 0 1 decap_w0
xfeed_4126 0 1 decap_w0
xfeed_4125 0 1 tie
xfeed_4124 0 1 decap_w0
xfeed_4123 0 1 decap_w0
xfeed_4122 0 1 decap_w0
xfeed_4121 0 1 decap_w0
xfeed_4120 0 1 decap_w0
xfeed_2989 0 1 decap_w0
xfeed_2988 0 1 decap_w0
xfeed_2987 0 1 decap_w0
xfeed_2986 0 1 decap_w0
xfeed_2985 0 1 decap_w0
xfeed_2984 0 1 decap_w0
xfeed_2983 0 1 decap_w0
xfeed_2982 0 1 decap_w0
xfeed_2981 0 1 decap_w0
xfeed_2980 0 1 decap_w0
xsubckt_102_and2_x1 0 1 688 1916 771 and2_x1
xsubckt_511_and3_x1 0 1 240 373 336 241 and3_x1
xsubckt_593_or21nand_x0 0 1 162 2053 601 163 or21nand_x0
xsubckt_1761_nexor2_x0 0 1 833 936 835 nexor2_x0
xfeed_10339 0 1 tie
xfeed_10338 0 1 decap_w0
xfeed_10337 0 1 decap_w0
xfeed_10336 0 1 decap_w0
xfeed_10335 0 1 decap_w0
xfeed_10334 0 1 decap_w0
xfeed_10333 0 1 decap_w0
xfeed_10332 0 1 decap_w0
xfeed_10331 0 1 decap_w0
xfeed_10330 0 1 decap_w0
xfeed_969 0 1 decap_w0
xfeed_968 0 1 tie
xfeed_967 0 1 decap_w0
xfeed_966 0 1 decap_w0
xfeed_965 0 1 decap_w0
xfeed_964 0 1 decap_w0
xfeed_963 0 1 decap_w0
xfeed_962 0 1 decap_w0
xfeed_961 0 1 decap_w0
xfeed_960 0 1 tie
xsubckt_1058_or21nand_x0 0 1 1484 532 1532 1485 or21nand_x0
xsubckt_224_mux2_x1 0 1 527 1989 1998 1986 mux2_x1
xsubckt_507_and3_x1 0 1 244 248 247 245 and3_x1
xsubckt_1380_and2_x1 0 1 1210 1216 1211 and2_x1
xsubckt_1403_nand2_x0 0 1 1189 2049 479 nand2_x0
xsubckt_1459_or21nand_x0 0 1 1137 2013 1140 1138 or21nand_x0
xsubckt_1667_nand3_x0 0 1 927 1974 680 595 nand3_x0
xfeed_8449 0 1 decap_w0
xfeed_8448 0 1 decap_w0
xfeed_8447 0 1 decap_w0
xfeed_8446 0 1 decap_w0
xfeed_8445 0 1 decap_w0
xfeed_8444 0 1 decap_w0
xfeed_8443 0 1 decap_w0
xfeed_8442 0 1 decap_w0
xfeed_8441 0 1 decap_w0
xfeed_8440 0 1 decap_w0
xfeed_7919 0 1 tie
xfeed_7918 0 1 decap_w0
xfeed_7917 0 1 decap_w0
xfeed_7916 0 1 decap_w0
xfeed_7915 0 1 tie
xfeed_7914 0 1 decap_w0
xfeed_7913 0 1 decap_w0
xfeed_7912 0 1 decap_w0
xfeed_7911 0 1 decap_w0
xfeed_7910 0 1 tie
xfeed_4139 0 1 decap_w0
xfeed_4138 0 1 decap_w0
xfeed_4137 0 1 decap_w0
xfeed_4136 0 1 decap_w0
xfeed_4135 0 1 decap_w0
xfeed_4134 0 1 decap_w0
xfeed_4133 0 1 decap_w0
xfeed_4132 0 1 tie
xfeed_4131 0 1 decap_w0
xfeed_4130 0 1 decap_w0
xfeed_3609 0 1 decap_w0
xfeed_3608 0 1 decap_w0
xfeed_3607 0 1 decap_w0
xfeed_3606 0 1 decap_w0
xfeed_3605 0 1 decap_w0
xfeed_3604 0 1 decap_w0
xfeed_3603 0 1 decap_w0
xfeed_3602 0 1 decap_w0
xfeed_3601 0 1 decap_w0
xfeed_3600 0 1 decap_w0
xfeed_2998 0 1 tie
xfeed_2997 0 1 decap_w0
xfeed_2996 0 1 decap_w0
xfeed_2995 0 1 decap_w0
xfeed_2994 0 1 decap_w0
xfeed_2993 0 1 decap_w0
xfeed_2992 0 1 decap_w0
xfeed_2991 0 1 tie
xfeed_2990 0 1 decap_w0
xsubckt_276_nand3_x0 0 1 472 678 490 473 nand3_x0
xsubckt_1711_and3_x1 0 1 883 1070 899 898 and3_x1
xfeed_10349 0 1 decap_w0
xfeed_10348 0 1 decap_w0
xfeed_10347 0 1 decap_w0
xfeed_10346 0 1 decap_w0
xfeed_10345 0 1 decap_w0
xfeed_10344 0 1 decap_w0
xfeed_10343 0 1 decap_w0
xfeed_10342 0 1 decap_w0
xfeed_10341 0 1 decap_w0
xfeed_10340 0 1 decap_w0
xfeed_2999 0 1 decap_w0
xfeed_979 0 1 decap_w0
xfeed_978 0 1 decap_w0
xfeed_977 0 1 decap_w0
xfeed_976 0 1 decap_w0
xfeed_975 0 1 tie
xfeed_974 0 1 decap_w0
xfeed_973 0 1 decap_w0
xfeed_972 0 1 decap_w0
xfeed_971 0 1 decap_w0
xfeed_970 0 1 decap_w0
xsubckt_1158_or21nand_x0 0 1 1403 1407 1409 1960 or21nand_x0
xsubckt_850_and3_x1 0 1 1629 2066 682 490 and3_x1
xsubckt_301_and4_x1 0 1 447 1929 715 1927 713 and4_x1
xfeed_8459 0 1 decap_w0
xfeed_8458 0 1 decap_w0
xfeed_8457 0 1 decap_w0
xfeed_8456 0 1 decap_w0
xfeed_8455 0 1 decap_w0
xfeed_8454 0 1 decap_w0
xfeed_8453 0 1 decap_w0
xfeed_8452 0 1 decap_w0
xfeed_8451 0 1 decap_w0
xfeed_8450 0 1 decap_w0
xfeed_7929 0 1 decap_w0
xfeed_7928 0 1 decap_w0
xfeed_7927 0 1 decap_w0
xfeed_7926 0 1 decap_w0
xfeed_7925 0 1 decap_w0
xfeed_7924 0 1 decap_w0
xfeed_7923 0 1 tie
xfeed_7922 0 1 decap_w0
xfeed_7921 0 1 decap_w0
xfeed_4148 0 1 decap_w0
xfeed_4147 0 1 decap_w0
xfeed_4146 0 1 decap_w0
xfeed_4145 0 1 decap_w0
xfeed_4144 0 1 tie
xfeed_4143 0 1 decap_w0
xfeed_4142 0 1 decap_w0
xfeed_4141 0 1 decap_w0
xfeed_4140 0 1 decap_w0
xfeed_3619 0 1 decap_w0
xfeed_3618 0 1 decap_w0
xfeed_3617 0 1 decap_w0
xfeed_3616 0 1 decap_w0
xfeed_3615 0 1 decap_w0
xfeed_3614 0 1 decap_w0
xfeed_3613 0 1 decap_w0
xfeed_3612 0 1 decap_w0
xfeed_3610 0 1 decap_w0
xsubckt_1462_or21nand_x0 0 1 1134 1136 1135 1745 or21nand_x0
xfeed_10359 0 1 decap_w0
xfeed_10358 0 1 decap_w0
xfeed_10357 0 1 decap_w0
xfeed_10356 0 1 decap_w0
xfeed_10355 0 1 decap_w0
xfeed_10354 0 1 decap_w0
xfeed_10353 0 1 decap_w0
xfeed_10352 0 1 decap_w0
xfeed_10351 0 1 decap_w0
xfeed_10350 0 1 decap_w0
xfeed_989 0 1 decap_w0
xfeed_988 0 1 decap_w0
xfeed_987 0 1 decap_w0
xfeed_986 0 1 decap_w0
xfeed_985 0 1 decap_w0
xfeed_984 0 1 decap_w0
xfeed_983 0 1 decap_w0
xfeed_982 0 1 tie
xfeed_981 0 1 decap_w0
xfeed_980 0 1 decap_w0
xsubckt_920_mux2_x1 0 1 1896 1612 2036 1579 mux2_x1
xsubckt_1729_and2_x1 0 1 865 1101 866 and2_x1
xsubckt_1951_dff_x1 0 1 2055 1797 45 dff_x1
xsubckt_1953_dff_x1 0 1 2052 1795 45 dff_x1
xfeed_8469 0 1 decap_w0
xfeed_8468 0 1 decap_w0
xfeed_8467 0 1 decap_w0
xfeed_8466 0 1 decap_w0
xfeed_8465 0 1 tie
xfeed_8464 0 1 tie
xfeed_8463 0 1 decap_w0
xfeed_8462 0 1 decap_w0
xfeed_8461 0 1 decap_w0
xfeed_8460 0 1 decap_w0
xfeed_7939 0 1 decap_w0
xfeed_7938 0 1 decap_w0
xfeed_7937 0 1 decap_w0
xfeed_7936 0 1 decap_w0
xfeed_7935 0 1 tie
xfeed_7934 0 1 decap_w0
xfeed_7933 0 1 decap_w0
xfeed_7932 0 1 decap_w0
xfeed_7931 0 1 decap_w0
xfeed_7930 0 1 tie
xfeed_4159 0 1 decap_w0
xfeed_4158 0 1 decap_w0
xfeed_4157 0 1 decap_w0
xfeed_4156 0 1 decap_w0
xfeed_4155 0 1 decap_w0
xfeed_4154 0 1 decap_w0
xfeed_4153 0 1 decap_w0
xfeed_4152 0 1 decap_w0
xfeed_4151 0 1 decap_w0
xfeed_4150 0 1 decap_w0
xfeed_3629 0 1 decap_w0
xfeed_3628 0 1 decap_w0
xfeed_3627 0 1 tie
xfeed_3626 0 1 decap_w0
xfeed_3625 0 1 decap_w0
xfeed_3624 0 1 decap_w0
xfeed_3623 0 1 decap_w0
xfeed_3622 0 1 decap_w0
xfeed_3621 0 1 decap_w0
xfeed_3620 0 1 decap_w0
xsubckt_1200_or2_x1 0 1 1364 1367 1365 or2_x1
xsubckt_1161_or21nand_x0 0 1 1400 780 606 494 or21nand_x0
xsubckt_319_and3_x1 0 1 429 609 598 557 and3_x1
xsubckt_179_nand2_x0 0 1 579 616 581 nand2_x0
xsubckt_609_nor2_x0 0 1 147 149 148 nor2_x0
xsubckt_1794_nexor2_x0 0 1 800 817 813 nexor2_x0
xsubckt_1955_dff_x1 0 1 2050 1793 35 dff_x1
xsubckt_1957_dff_x1 0 1 2048 1791 35 dff_x1
xsubckt_1959_dff_x1 0 1 2046 1789 35 dff_x1
xdiode_9 0 1 610 diode_w1
xdiode_8 0 1 610 diode_w1
xdiode_7 0 1 610 diode_w1
xdiode_6 0 1 609 diode_w1
xdiode_5 0 1 609 diode_w1
xdiode_4 0 1 609 diode_w1
xdiode_3 0 1 608 diode_w1
xdiode_2 0 1 608 diode_w1
xdiode_1 0 1 608 diode_w1
xdiode_0 0 1 608 diode_w1
xfeed_10369 0 1 decap_w0
xfeed_10368 0 1 decap_w0
xfeed_10367 0 1 decap_w0
xfeed_10366 0 1 decap_w0
xfeed_10365 0 1 decap_w0
xfeed_10364 0 1 decap_w0
xfeed_10363 0 1 decap_w0
xfeed_10362 0 1 decap_w0
xfeed_10361 0 1 decap_w0
xfeed_10360 0 1 decap_w0
xfeed_999 0 1 decap_w0
xfeed_998 0 1 decap_w0
xfeed_997 0 1 decap_w0
xfeed_996 0 1 decap_w0
xfeed_995 0 1 decap_w0
xfeed_994 0 1 decap_w0
xfeed_993 0 1 decap_w0
xfeed_992 0 1 decap_w0
xfeed_990 0 1 decap_w0
xsubckt_1240_mux2_x1 0 1 1821 2091 2072 1334 mux2_x1
xsubckt_1022_nand3_x0 0 1 1511 1526 1525 1512 nand3_x0
xsubckt_916_mux2_x1 0 1 1899 1586 2039 1580 mux2_x1
xsubckt_689_or21nand_x0 0 1 1774 1985 436 167 or21nand_x0
xsubckt_663_or2_x1 0 1 97 762 109 or2_x1
xsubckt_661_or2_x1 0 1 99 728 212 or2_x1
xsubckt_149_and21nor_x0 0 1 619 663 628 620 and21nor_x0
xsubckt_1643_nand2_x0 0 1 951 1101 953 nand2_x0
xsubckt_1662_or21nand_x0 0 1 932 1663 1116 694 or21nand_x0
xsubckt_1776_nexor2_x0 0 1 818 977 972 nexor2_x0
xfeed_8479 0 1 decap_w0
xfeed_8478 0 1 decap_w0
xfeed_8477 0 1 decap_w0
xfeed_8476 0 1 tie
xfeed_8475 0 1 decap_w0
xfeed_8474 0 1 decap_w0
xfeed_8473 0 1 decap_w0
xfeed_8472 0 1 decap_w0
xfeed_8471 0 1 decap_w0
xfeed_8470 0 1 decap_w0
xfeed_7949 0 1 decap_w0
xfeed_7948 0 1 decap_w0
xfeed_7947 0 1 decap_w0
xfeed_7946 0 1 decap_w0
xfeed_7945 0 1 decap_w0
xfeed_7944 0 1 decap_w0
xfeed_7943 0 1 decap_w0
xfeed_7942 0 1 decap_w0
xfeed_7941 0 1 decap_w0
xfeed_7940 0 1 tie
xfeed_4169 0 1 decap_w0
xfeed_4168 0 1 decap_w0
xfeed_4167 0 1 decap_w0
xfeed_4166 0 1 decap_w0
xfeed_4165 0 1 decap_w0
xfeed_4164 0 1 decap_w0
xfeed_4163 0 1 decap_w0
xfeed_4162 0 1 decap_w0
xfeed_4161 0 1 decap_w0
xfeed_4160 0 1 decap_w0
xfeed_3639 0 1 decap_w0
xfeed_3638 0 1 decap_w0
xfeed_3637 0 1 decap_w0
xfeed_3636 0 1 decap_w0
xfeed_3635 0 1 decap_w0
xfeed_3634 0 1 tie
xfeed_3633 0 1 decap_w0
xfeed_3632 0 1 decap_w0
xfeed_3631 0 1 decap_w0
xfeed_3630 0 1 decap_w0
xsubckt_1236_mux2_x1 0 1 1825 2095 2060 1334 mux2_x1
xsubckt_1188_and2_x1 0 1 1376 456 1380 and2_x1
xsubckt_191_and4_x1 0 1 567 716 1924 599 568 and4_x1
xsubckt_1597_and3_x1 0 1 997 1005 1001 999 and3_x1
xsubckt_1767_nexor2_x0 0 1 827 840 836 nexor2_x0
xfeed_10379 0 1 decap_w0
xfeed_10378 0 1 decap_w0
xfeed_10377 0 1 decap_w0
xfeed_10376 0 1 tie
xfeed_10375 0 1 decap_w0
xfeed_10374 0 1 decap_w0
xfeed_10372 0 1 decap_w0
xfeed_10371 0 1 decap_w0
xfeed_10370 0 1 decap_w0
xsubckt_700_or21nand_x0 0 1 1764 609 490 451 or21nand_x0
xsubckt_187_and4_x1 0 1 571 1929 1924 1927 1928 and4_x1
xsubckt_1405_and4_x1 0 1 1187 435 1649 1189 1188 and4_x1
xsubckt_1463_nand2_x0 0 1 1133 755 1134 nand2_x0
xsubckt_1758_nexor2_x0 0 1 836 915 909 nexor2_x0
xfeed_8489 0 1 decap_w0
xfeed_8488 0 1 decap_w0
xfeed_8487 0 1 decap_w0
xfeed_8486 0 1 decap_w0
xfeed_8485 0 1 decap_w0
xfeed_8484 0 1 decap_w0
xfeed_8483 0 1 decap_w0
xfeed_8482 0 1 decap_w0
xfeed_8481 0 1 decap_w0
xfeed_8480 0 1 tie
xfeed_7959 0 1 tie
xfeed_7958 0 1 decap_w0
xfeed_7957 0 1 decap_w0
xfeed_7956 0 1 decap_w0
xfeed_7955 0 1 decap_w0
xfeed_7954 0 1 decap_w0
xfeed_7953 0 1 decap_w0
xfeed_7952 0 1 decap_w0
xfeed_7951 0 1 decap_w0
xfeed_7950 0 1 decap_w0
xfeed_4179 0 1 decap_w0
xfeed_4178 0 1 decap_w0
xfeed_4177 0 1 decap_w0
xfeed_4176 0 1 decap_w0
xfeed_4175 0 1 decap_w0
xfeed_4174 0 1 decap_w0
xfeed_4173 0 1 decap_w0
xfeed_4172 0 1 decap_w0
xfeed_4170 0 1 decap_w0
xfeed_3649 0 1 decap_w0
xfeed_3648 0 1 decap_w0
xfeed_3647 0 1 decap_w0
xfeed_3645 0 1 decap_w0
xfeed_3644 0 1 decap_w0
xfeed_3643 0 1 decap_w0
xfeed_3642 0 1 decap_w0
xfeed_3641 0 1 tie
xfeed_3640 0 1 decap_w0
xsubckt_1105_nand2_x0 0 1 1443 503 430 nand2_x0
xsubckt_1373_nand2_x0 0 1 1217 775 1980 nand2_x0
xsubckt_1712_nand3_x0 0 1 882 1070 899 898 nand3_x0
xfeed_10389 0 1 decap_w0
xfeed_10388 0 1 decap_w0
xfeed_10387 0 1 decap_w0
xfeed_10386 0 1 decap_w0
xfeed_10385 0 1 decap_w0
xfeed_10384 0 1 decap_w0
xfeed_10382 0 1 decap_w0
xfeed_10381 0 1 decap_w0
xfeed_10380 0 1 decap_w0
xsubckt_1453_and2_x1 0 1 1143 547 1745 and2_x1
xfeed_9109 0 1 decap_w0
xfeed_9108 0 1 decap_w0
xfeed_9107 0 1 decap_w0
xfeed_9106 0 1 decap_w0
xfeed_9105 0 1 decap_w0
xfeed_9104 0 1 decap_w0
xfeed_9103 0 1 decap_w0
xfeed_9102 0 1 tie
xfeed_9101 0 1 decap_w0
xfeed_9100 0 1 decap_w0
xfeed_8499 0 1 decap_w0
xfeed_8498 0 1 decap_w0
xfeed_8497 0 1 decap_w0
xfeed_8496 0 1 decap_w0
xfeed_8495 0 1 decap_w0
xfeed_8494 0 1 decap_w0
xfeed_8493 0 1 decap_w0
xfeed_8492 0 1 tie
xfeed_8490 0 1 decap_w0
xfeed_7969 0 1 decap_w0
xfeed_7968 0 1 decap_w0
xfeed_7967 0 1 decap_w0
xfeed_7966 0 1 decap_w0
xfeed_7965 0 1 decap_w0
xfeed_7964 0 1 decap_w0
xfeed_7963 0 1 decap_w0
xfeed_7962 0 1 decap_w0
xfeed_7961 0 1 decap_w0
xfeed_7960 0 1 decap_w0
xfeed_4189 0 1 decap_w0
xfeed_4188 0 1 decap_w0
xfeed_4187 0 1 decap_w0
xfeed_4186 0 1 decap_w0
xfeed_4185 0 1 decap_w0
xfeed_4184 0 1 decap_w0
xfeed_4183 0 1 decap_w0
xfeed_4182 0 1 decap_w0
xfeed_4181 0 1 decap_w0
xfeed_4180 0 1 decap_w0
xfeed_3659 0 1 decap_w0
xfeed_3657 0 1 decap_w0
xfeed_3656 0 1 tie
xfeed_3654 0 1 decap_w0
xfeed_3653 0 1 decap_w0
xfeed_3651 0 1 decap_w0
xfeed_3650 0 1 decap_w0
xsubckt_762_nand2_x0 0 1 1706 1708 1707 nand2_x0
xsubckt_157_and2_x1 0 1 604 1929 715 and2_x1
xfeed_11009 0 1 decap_w0
xfeed_11008 0 1 decap_w0
xfeed_11007 0 1 tie
xfeed_11006 0 1 decap_w0
xfeed_11005 0 1 decap_w0
xfeed_11004 0 1 decap_w0
xfeed_11003 0 1 decap_w0
xfeed_11002 0 1 decap_w0
xfeed_11001 0 1 decap_w0
xfeed_11000 0 1 tie
xfeed_10398 0 1 decap_w0
xfeed_10397 0 1 decap_w0
xfeed_10396 0 1 decap_w0
xfeed_10395 0 1 decap_w0
xfeed_10394 0 1 decap_w0
xfeed_10393 0 1 decap_w0
xfeed_10392 0 1 tie
xfeed_10391 0 1 decap_w0
xfeed_10390 0 1 decap_w0
xfeed_9119 0 1 decap_w0
xfeed_9118 0 1 decap_w0
xfeed_9117 0 1 decap_w0
xfeed_9116 0 1 decap_w0
xfeed_9115 0 1 tie
xfeed_9114 0 1 decap_w0
xfeed_9113 0 1 decap_w0
xfeed_9112 0 1 decap_w0
xfeed_9111 0 1 decap_w0
xfeed_9110 0 1 tie
xfeed_7977 0 1 decap_w0
xfeed_7976 0 1 decap_w0
xfeed_7975 0 1 decap_w0
xfeed_7974 0 1 decap_w0
xfeed_7973 0 1 decap_w0
xfeed_7972 0 1 decap_w0
xfeed_7971 0 1 decap_w0
xfeed_7970 0 1 decap_w0
xfeed_4199 0 1 decap_w0
xfeed_4198 0 1 decap_w0
xfeed_4197 0 1 decap_w0
xfeed_4196 0 1 decap_w0
xfeed_4195 0 1 decap_w0
xfeed_4194 0 1 decap_w0
xfeed_4193 0 1 decap_w0
xfeed_4192 0 1 tie
xfeed_4191 0 1 decap_w0
xfeed_4190 0 1 decap_w0
xfeed_3668 0 1 tie
xfeed_3667 0 1 decap_w0
xfeed_3666 0 1 decap_w0
xfeed_3665 0 1 decap_w0
xfeed_3664 0 1 decap_w0
xfeed_3663 0 1 decap_w0
xfeed_3662 0 1 decap_w0
xfeed_3661 0 1 tie
xfeed_3660 0 1 decap_w0
xsubckt_813_or4_x1 0 1 1661 1666 1665 1664 1662 or4_x1
xsubckt_668_nand3_x0 0 1 93 2015 184 177 nand3_x0
xsubckt_98_mux2_x1 0 1 690 720 719 774 mux2_x1
xsubckt_1561_or21nand_x0 0 1 1033 1035 1036 1075 or21nand_x0
xsubckt_1619_and21nor_x0 0 1 975 1070 986 1073 and21nor_x0
xfeed_11019 0 1 decap_w0
xfeed_11018 0 1 decap_w0
xfeed_11017 0 1 decap_w0
xfeed_11016 0 1 decap_w0
xfeed_11015 0 1 decap_w0
xfeed_11014 0 1 decap_w0
xfeed_11013 0 1 decap_w0
xfeed_11012 0 1 decap_w0
xfeed_11011 0 1 decap_w0
xfeed_11010 0 1 decap_w0
xfeed_7979 0 1 decap_w0
xfeed_7978 0 1 decap_w0
xsubckt_1121_and21nor_x0 0 1 1436 666 608 495 and21nor_x0
xsubckt_831_and3_x1 0 1 1646 1977 1749 1739 and3_x1
xsubckt_688_or21nand_x0 0 1 1775 2046 601 163 or21nand_x0
xfeed_9129 0 1 decap_w0
xfeed_9128 0 1 decap_w0
xfeed_9127 0 1 decap_w0
xfeed_9126 0 1 decap_w0
xfeed_9125 0 1 decap_w0
xfeed_9124 0 1 decap_w0
xfeed_9123 0 1 decap_w0
xfeed_9122 0 1 decap_w0
xfeed_9121 0 1 decap_w0
xfeed_9120 0 1 decap_w0
xfeed_7984 0 1 tie
xfeed_7983 0 1 decap_w0
xfeed_7982 0 1 decap_w0
xfeed_7981 0 1 decap_w0
xfeed_7980 0 1 decap_w0
xfeed_3679 0 1 decap_w0
xfeed_3678 0 1 decap_w0
xfeed_3677 0 1 decap_w0
xfeed_3676 0 1 decap_w0
xfeed_3675 0 1 tie
xfeed_3674 0 1 decap_w0
xfeed_3673 0 1 decap_w0
xfeed_3672 0 1 decap_w0
xfeed_3671 0 1 decap_w0
xfeed_3670 0 1 decap_w0
xsubckt_1125_and4_x1 0 1 1432 682 674 670 1433 and4_x1
xsubckt_791_and4_x1 0 1 1681 537 198 1769 1682 and4_x1
xsubckt_398_nand3_x0 0 1 351 563 354 352 nand3_x0
xsubckt_496_and2_x1 0 1 255 259 256 and2_x1
xsubckt_591_or21nand_x0 0 1 164 2013 436 167 or21nand_x0
xsubckt_1719_and21nor_x0 0 1 875 876 1121 168 and21nor_x0
xfeed_11029 0 1 decap_w0
xfeed_11028 0 1 decap_w0
xfeed_11027 0 1 decap_w0
xfeed_11026 0 1 decap_w0
xfeed_11025 0 1 decap_w0
xfeed_11024 0 1 decap_w0
xfeed_11023 0 1 decap_w0
xfeed_11022 0 1 tie
xfeed_11021 0 1 decap_w0
xfeed_11020 0 1 decap_w0
xfeed_7989 0 1 decap_w0
xfeed_7988 0 1 decap_w0
xfeed_7987 0 1 decap_w0
xfeed_7986 0 1 decap_w0
xfeed_7985 0 1 decap_w0
xsubckt_901_mux2_x1 0 1 1586 1587 1997 445 mux2_x1
xsubckt_1622_and2_x1 0 1 972 974 973 and2_x1
xsubckt_1658_nexor2_x0 0 1 936 947 941 nexor2_x0
xfeed_9139 0 1 decap_w0
xfeed_9138 0 1 decap_w0
xfeed_9137 0 1 decap_w0
xfeed_9136 0 1 decap_w0
xfeed_9135 0 1 decap_w0
xfeed_9134 0 1 decap_w0
xfeed_9133 0 1 decap_w0
xfeed_9132 0 1 decap_w0
xfeed_9131 0 1 decap_w0
xfeed_9130 0 1 decap_w0
xfeed_8609 0 1 decap_w0
xfeed_8607 0 1 decap_w0
xfeed_8606 0 1 decap_w0
xfeed_8605 0 1 decap_w0
xfeed_8604 0 1 decap_w0
xfeed_8603 0 1 decap_w0
xfeed_8602 0 1 tie
xfeed_8601 0 1 decap_w0
xfeed_8600 0 1 decap_w0
xfeed_7991 0 1 decap_w0
xfeed_7990 0 1 decap_w0
xfeed_3689 0 1 decap_w0
xfeed_3688 0 1 decap_w0
xfeed_3687 0 1 tie
xfeed_3686 0 1 decap_w0
xfeed_3685 0 1 decap_w0
xfeed_3684 0 1 decap_w0
xfeed_3683 0 1 decap_w0
xfeed_3682 0 1 decap_w0
xfeed_3681 0 1 decap_w0
xfeed_3680 0 1 decap_w0
xsubckt_1173_and2_x1 0 1 1389 1391 1390 and2_x1
xsubckt_849_and2_x1 0 1 1630 2046 1740 and2_x1
xsubckt_326_and2_x1 0 1 422 424 423 and2_x1
xfeed_11039 0 1 decap_w0
xfeed_11038 0 1 decap_w0
xfeed_11037 0 1 decap_w0
xfeed_11036 0 1 decap_w0
xfeed_11035 0 1 decap_w0
xfeed_11034 0 1 decap_w0
xfeed_11033 0 1 decap_w0
xfeed_11032 0 1 decap_w0
xfeed_11031 0 1 decap_w0
xfeed_11030 0 1 decap_w0
xfeed_10509 0 1 decap_w0
xfeed_10508 0 1 decap_w0
xfeed_10507 0 1 decap_w0
xfeed_10506 0 1 decap_w0
xfeed_10505 0 1 decap_w0
xfeed_10504 0 1 decap_w0
xfeed_10503 0 1 decap_w0
xfeed_10502 0 1 decap_w0
xfeed_10500 0 1 decap_w0
xfeed_7999 0 1 decap_w0
xfeed_7998 0 1 decap_w0
xfeed_7997 0 1 decap_w0
xfeed_7996 0 1 decap_w0
xfeed_7995 0 1 decap_w0
xfeed_7994 0 1 decap_w0
xfeed_7993 0 1 decap_w0
xfeed_7992 0 1 decap_w0
xsubckt_291_nand3_x0 0 1 457 687 616 460 nand3_x0
xsubckt_1361_or2_x1 0 1 1228 695 1323 or2_x1
xfeed_9149 0 1 decap_w0
xfeed_9148 0 1 decap_w0
xfeed_9147 0 1 decap_w0
xfeed_9146 0 1 decap_w0
xfeed_9145 0 1 decap_w0
xfeed_9144 0 1 decap_w0
xfeed_9143 0 1 decap_w0
xfeed_9142 0 1 tie
xfeed_9141 0 1 decap_w0
xfeed_9140 0 1 decap_w0
xfeed_8619 0 1 decap_w0
xfeed_8618 0 1 decap_w0
xfeed_8617 0 1 decap_w0
xfeed_8616 0 1 tie
xfeed_8615 0 1 decap_w0
xfeed_8614 0 1 decap_w0
xfeed_8613 0 1 decap_w0
xfeed_8612 0 1 decap_w0
xfeed_8611 0 1 decap_w0
xfeed_8610 0 1 decap_w0
xfeed_4309 0 1 decap_w0
xfeed_4308 0 1 decap_w0
xfeed_4307 0 1 decap_w0
xfeed_4306 0 1 decap_w0
xfeed_4305 0 1 decap_w0
xfeed_4304 0 1 decap_w0
xfeed_4303 0 1 decap_w0
xfeed_4302 0 1 tie
xfeed_4301 0 1 decap_w0
xfeed_4300 0 1 decap_w0
xfeed_3698 0 1 tie
xfeed_3697 0 1 decap_w0
xfeed_3696 0 1 decap_w0
xfeed_3695 0 1 decap_w0
xfeed_3694 0 1 decap_w0
xfeed_3693 0 1 decap_w0
xfeed_3691 0 1 tie
xfeed_3690 0 1 decap_w0
xsubckt_998_nand3_x0 0 1 1531 643 313 1532 nand3_x0
xsubckt_40_inv_x0 0 1 742 2068 inv_x0
xsubckt_630_nand4_x0 0 1 128 133 132 131 130 nand4_x0
xfeed_11049 0 1 tie
xfeed_11048 0 1 decap_w0
xfeed_11047 0 1 decap_w0
xfeed_11046 0 1 decap_w0
xfeed_11045 0 1 decap_w0
xfeed_11044 0 1 decap_w0
xfeed_11043 0 1 decap_w0
xfeed_11042 0 1 decap_w0
xfeed_11041 0 1 decap_w0
xfeed_11040 0 1 decap_w0
xfeed_10519 0 1 decap_w0
xfeed_10518 0 1 decap_w0
xfeed_10517 0 1 tie
xfeed_10516 0 1 decap_w0
xfeed_10515 0 1 decap_w0
xfeed_10514 0 1 decap_w0
xfeed_10513 0 1 decap_w0
xfeed_10512 0 1 decap_w0
xfeed_10511 0 1 decap_w0
xfeed_10510 0 1 decap_w0
xfeed_3699 0 1 decap_w0
xsubckt_879_mux2_x1 0 1 1911 2019 1605 1619 mux2_x1
xsubckt_46_inv_x0 0 1 736 1942 inv_x0
xsubckt_44_inv_x0 0 1 738 1944 inv_x0
xsubckt_42_inv_x0 0 1 740 2066 inv_x0
xsubckt_554_nand2_x0 0 1 1914 207 201 nand2_x0
xsubckt_1657_or21nand_x0 0 1 937 947 946 943 or21nand_x0
xfeed_9159 0 1 decap_w0
xfeed_9158 0 1 decap_w0
xfeed_9157 0 1 decap_w0
xfeed_9156 0 1 decap_w0
xfeed_9155 0 1 decap_w0
xfeed_9154 0 1 decap_w0
xfeed_9153 0 1 decap_w0
xfeed_9152 0 1 decap_w0
xfeed_9151 0 1 decap_w0
xfeed_9150 0 1 decap_w0
xfeed_8629 0 1 decap_w0
xfeed_8628 0 1 decap_w0
xfeed_8627 0 1 decap_w0
xfeed_8626 0 1 decap_w0
xfeed_8625 0 1 tie
xfeed_8624 0 1 decap_w0
xfeed_8623 0 1 decap_w0
xfeed_8622 0 1 decap_w0
xfeed_8621 0 1 decap_w0
xfeed_8620 0 1 tie
xfeed_4319 0 1 decap_w0
xfeed_4318 0 1 decap_w0
xfeed_4317 0 1 tie
xfeed_4316 0 1 decap_w0
xfeed_4315 0 1 decap_w0
xfeed_4314 0 1 decap_w0
xfeed_4313 0 1 decap_w0
xfeed_4312 0 1 decap_w0
xfeed_4311 0 1 decap_w0
xfeed_4310 0 1 decap_w0
xsubckt_803_nand3_x0 0 1 1670 2072 679 490 nand3_x0
xsubckt_186_or21nand_x0 0 1 572 574 597 676 or21nand_x0
xsubckt_48_inv_x0 0 1 734 1968 inv_x0
xsubckt_525_and4_x1 0 1 227 461 457 419 416 and4_x1
xsubckt_1560_or21nand_x0 0 1 1034 1067 1046 1072 or21nand_x0
xsubckt_1675_nand2_x0 0 1 919 1101 921 nand2_x0
xfeed_11059 0 1 decap_w0
xfeed_11058 0 1 decap_w0
xfeed_11057 0 1 decap_w0
xfeed_11056 0 1 decap_w0
xfeed_11055 0 1 decap_w0
xfeed_11054 0 1 decap_w0
xfeed_11053 0 1 decap_w0
xfeed_11052 0 1 decap_w0
xfeed_11051 0 1 decap_w0
xfeed_11050 0 1 decap_w0
xfeed_10529 0 1 decap_w0
xfeed_10528 0 1 decap_w0
xfeed_10527 0 1 decap_w0
xfeed_10526 0 1 decap_w0
xfeed_10525 0 1 decap_w0
xfeed_10524 0 1 decap_w0
xfeed_10523 0 1 decap_w0
xfeed_10522 0 1 decap_w0
xfeed_10521 0 1 decap_w0
xfeed_10520 0 1 decap_w0
xsubckt_891_nand3_x0 0 1 1595 1962 2048 1598 nand3_x0
xsubckt_852_and21nor_x0 0 1 1627 740 600 1745 and21nor_x0
xsubckt_270_nand4_x0 0 1 478 714 1928 678 589 nand4_x0
xsubckt_1556_mux2_x1 0 1 1038 1041 1044 1052 mux2_x1
xsubckt_1757_or21nand_x0 0 1 837 915 914 911 or21nand_x0
xfeed_9169 0 1 decap_w0
xfeed_9168 0 1 decap_w0
xfeed_9167 0 1 decap_w0
xfeed_9166 0 1 decap_w0
xfeed_9165 0 1 decap_w0
xfeed_9164 0 1 decap_w0
xfeed_9163 0 1 decap_w0
xfeed_9162 0 1 tie
xfeed_9161 0 1 decap_w0
xfeed_9160 0 1 decap_w0
xfeed_8639 0 1 decap_w0
xfeed_8638 0 1 decap_w0
xfeed_8637 0 1 decap_w0
xfeed_8636 0 1 decap_w0
xfeed_8635 0 1 decap_w0
xfeed_8634 0 1 decap_w0
xfeed_8633 0 1 decap_w0
xfeed_8632 0 1 decap_w0
xfeed_8631 0 1 decap_w0
xfeed_8630 0 1 tie
xfeed_4329 0 1 tie
xfeed_4328 0 1 decap_w0
xfeed_4327 0 1 decap_w0
xfeed_4326 0 1 decap_w0
xfeed_4325 0 1 decap_w0
xfeed_4324 0 1 decap_w0
xfeed_4323 0 1 decap_w0
xfeed_4322 0 1 tie
xfeed_4321 0 1 decap_w0
xfeed_4320 0 1 decap_w0
xsubckt_982_and3_x1 0 1 1545 661 527 521 and3_x1
xsubckt_904_and3_x1 0 1 1584 1962 767 761 and3_x1
xsubckt_1495_nand2_x0 0 1 1101 1105 1103 nand2_x0
xfeed_11069 0 1 decap_w0
xfeed_11068 0 1 decap_w0
xfeed_11067 0 1 decap_w0
xfeed_11066 0 1 decap_w0
xfeed_11065 0 1 decap_w0
xfeed_11064 0 1 decap_w0
xfeed_11063 0 1 decap_w0
xfeed_11062 0 1 decap_w0
xfeed_11061 0 1 tie
xfeed_11060 0 1 decap_w0
xfeed_10539 0 1 decap_w0
xfeed_10538 0 1 decap_w0
xfeed_10537 0 1 decap_w0
xfeed_10536 0 1 decap_w0
xfeed_10535 0 1 decap_w0
xfeed_10534 0 1 decap_w0
xfeed_10533 0 1 decap_w0
xfeed_10532 0 1 decap_w0
xfeed_10531 0 1 decap_w0
xfeed_10530 0 1 decap_w0
xsubckt_890_and3_x1 0 1 1596 1962 2048 1598 and3_x1
xfeed_9179 0 1 decap_w0
xfeed_9178 0 1 decap_w0
xfeed_9177 0 1 decap_w0
xfeed_9176 0 1 decap_w0
xfeed_9175 0 1 decap_w0
xfeed_9174 0 1 tie
xfeed_9173 0 1 decap_w0
xfeed_9172 0 1 decap_w0
xfeed_9171 0 1 decap_w0
xfeed_9170 0 1 decap_w0
xfeed_8649 0 1 decap_w0
xfeed_8648 0 1 decap_w0
xfeed_8647 0 1 decap_w0
xfeed_8646 0 1 decap_w0
xfeed_8645 0 1 tie
xfeed_8644 0 1 decap_w0
xfeed_8643 0 1 decap_w0
xfeed_8642 0 1 decap_w0
xfeed_8641 0 1 decap_w0
xfeed_8640 0 1 decap_w0
xfeed_4339 0 1 decap_w0
xfeed_4338 0 1 decap_w0
xfeed_4337 0 1 decap_w0
xfeed_4336 0 1 decap_w0
xfeed_4335 0 1 decap_w0
xfeed_4334 0 1 decap_w0
xfeed_4333 0 1 tie
xfeed_4332 0 1 decap_w0
xfeed_4331 0 1 decap_w0
xfeed_4330 0 1 decap_w0
xfeed_3809 0 1 decap_w0
xfeed_3808 0 1 decap_w0
xfeed_3807 0 1 decap_w0
xfeed_3806 0 1 decap_w0
xfeed_3805 0 1 decap_w0
xfeed_3804 0 1 tie
xfeed_3803 0 1 decap_w0
xfeed_3802 0 1 decap_w0
xfeed_3801 0 1 decap_w0
xfeed_3800 0 1 decap_w0
xsubckt_1760_or21nand_x0 0 1 834 907 840 838 or21nand_x0
xfeed_11079 0 1 decap_w0
xfeed_11078 0 1 decap_w0
xfeed_11077 0 1 decap_w0
xfeed_11076 0 1 decap_w0
xfeed_11075 0 1 decap_w0
xfeed_11074 0 1 decap_w0
xfeed_11073 0 1 decap_w0
xfeed_11072 0 1 decap_w0
xfeed_11071 0 1 decap_w0
xfeed_11070 0 1 decap_w0
xfeed_10546 0 1 decap_w0
xfeed_10545 0 1 tie
xfeed_10544 0 1 decap_w0
xfeed_10543 0 1 decap_w0
xfeed_10542 0 1 decap_w0
xfeed_10541 0 1 decap_w0
xfeed_10540 0 1 decap_w0
xsubckt_653_nor2_x0 0 1 106 114 108 nor2_x0
xsubckt_347_and21nor_x0 0 1 401 402 558 567 and21nor_x0
xsubckt_1960_dff_x1 0 1 2054 1788 35 dff_x1
xfeed_10549 0 1 decap_w0
xfeed_10548 0 1 decap_w0
xfeed_10547 0 1 tie
xfeed_9189 0 1 decap_w0
xfeed_9188 0 1 decap_w0
xfeed_9187 0 1 decap_w0
xfeed_9186 0 1 decap_w0
xfeed_9185 0 1 decap_w0
xfeed_9184 0 1 decap_w0
xfeed_9183 0 1 decap_w0
xfeed_9182 0 1 decap_w0
xfeed_9181 0 1 decap_w0
xfeed_9180 0 1 decap_w0
xfeed_8659 0 1 decap_w0
xfeed_8658 0 1 decap_w0
xfeed_8657 0 1 decap_w0
xfeed_8656 0 1 decap_w0
xfeed_8655 0 1 tie
xfeed_8654 0 1 decap_w0
xfeed_8653 0 1 decap_w0
xfeed_8652 0 1 decap_w0
xfeed_8651 0 1 decap_w0
xfeed_8650 0 1 decap_w0
xfeed_4349 0 1 decap_w0
xfeed_4348 0 1 decap_w0
xfeed_4347 0 1 tie
xfeed_4346 0 1 decap_w0
xfeed_4345 0 1 decap_w0
xfeed_4344 0 1 decap_w0
xfeed_4343 0 1 decap_w0
xfeed_4342 0 1 decap_w0
xfeed_4340 0 1 tie
xfeed_3819 0 1 decap_w0
xfeed_3818 0 1 decap_w0
xfeed_3817 0 1 decap_w0
xfeed_3816 0 1 decap_w0
xfeed_3815 0 1 decap_w0
xfeed_3814 0 1 decap_w0
xfeed_3813 0 1 decap_w0
xfeed_3812 0 1 decap_w0
xfeed_3811 0 1 tie
xfeed_3810 0 1 decap_w0
xsubckt_1120_nand2_x0 0 1 1437 1960 548 nand2_x0
xsubckt_848_and21nor_x0 0 1 1631 689 1755 1754 and21nor_x0
xsubckt_1817_mux2_x1 0 1 1788 2054 820 775 mux2_x1
xfeed_11089 0 1 decap_w0
xfeed_11088 0 1 decap_w0
xfeed_11087 0 1 decap_w0
xfeed_11086 0 1 decap_w0
xfeed_11085 0 1 decap_w0
xfeed_11084 0 1 decap_w0
xfeed_11083 0 1 decap_w0
xfeed_11082 0 1 decap_w0
xfeed_11081 0 1 decap_w0
xfeed_11080 0 1 decap_w0
xfeed_10553 0 1 decap_w0
xfeed_10552 0 1 decap_w0
xfeed_10551 0 1 decap_w0
xfeed_10550 0 1 decap_w0
xsubckt_1723_nand4_x0 0 1 871 2003 1128 1098 1097 nand4_x0
xfeed_10559 0 1 decap_w0
xfeed_10558 0 1 decap_w0
xfeed_10557 0 1 decap_w0
xfeed_10556 0 1 decap_w0
xfeed_10555 0 1 decap_w0
xfeed_10554 0 1 tie
xfeed_9199 0 1 decap_w0
xfeed_9198 0 1 decap_w0
xfeed_9197 0 1 decap_w0
xfeed_9196 0 1 tie
xfeed_9195 0 1 decap_w0
xfeed_9194 0 1 decap_w0
xfeed_9193 0 1 decap_w0
xfeed_9192 0 1 decap_w0
xfeed_9191 0 1 decap_w0
xfeed_9190 0 1 decap_w0
xfeed_8669 0 1 decap_w0
xfeed_8668 0 1 decap_w0
xfeed_8667 0 1 decap_w0
xfeed_8666 0 1 decap_w0
xfeed_8665 0 1 decap_w0
xfeed_8664 0 1 decap_w0
xfeed_8663 0 1 decap_w0
xfeed_8662 0 1 decap_w0
xfeed_8661 0 1 decap_w0
xfeed_8660 0 1 decap_w0
xfeed_4359 0 1 decap_w0
xfeed_4358 0 1 decap_w0
xfeed_4357 0 1 decap_w0
xfeed_4356 0 1 decap_w0
xfeed_4355 0 1 decap_w0
xfeed_4353 0 1 decap_w0
xfeed_4352 0 1 decap_w0
xfeed_4351 0 1 decap_w0
xfeed_3829 0 1 decap_w0
xfeed_3828 0 1 tie
xfeed_3827 0 1 decap_w0
xfeed_3826 0 1 decap_w0
xfeed_3825 0 1 decap_w0
xfeed_3824 0 1 decap_w0
xfeed_3823 0 1 decap_w0
xfeed_3822 0 1 decap_w0
xfeed_3821 0 1 tie
xfeed_3820 0 1 decap_w0
xsubckt_949_nand4_x0 0 1 1570 660 654 529 528 nand4_x0
xsubckt_242_nand4_x0 0 1 509 1925 711 571 557 nand4_x0
xfeed_11099 0 1 decap_w0
xfeed_11098 0 1 decap_w0
xfeed_11097 0 1 decap_w0
xfeed_11096 0 1 tie
xfeed_11095 0 1 decap_w0
xfeed_11094 0 1 decap_w0
xfeed_11093 0 1 decap_w0
xfeed_11092 0 1 decap_w0
xfeed_11091 0 1 tie
xfeed_11090 0 1 decap_w0
xfeed_10560 0 1 decap_w0
xsubckt_1062_and2_x1 0 1 1480 1484 1481 and2_x1
xsubckt_864_mux2_x1 0 1 1913 2021 1618 1619 mux2_x1
xsubckt_287_or2_x1 0 1 461 554 462 or2_x1
xsubckt_215_and2_x1 0 1 539 560 540 and2_x1
xsubckt_166_nand2_x0 0 1 592 616 595 nand2_x0
xsubckt_1568_or2_x1 0 1 1026 691 1116 or2_x1
xsubckt_1810_nand2_x0 0 1 789 773 2049 nand2_x0
xfeed_10569 0 1 decap_w0
xfeed_10568 0 1 decap_w0
xfeed_10567 0 1 decap_w0
xfeed_10566 0 1 decap_w0
xfeed_10565 0 1 decap_w0
xfeed_10564 0 1 decap_w0
xfeed_10563 0 1 decap_w0
xfeed_10562 0 1 decap_w0
xfeed_10561 0 1 decap_w0
xfeed_8677 0 1 decap_w0
xfeed_8676 0 1 decap_w0
xfeed_8675 0 1 decap_w0
xfeed_8674 0 1 decap_w0
xfeed_8673 0 1 tie
xfeed_8672 0 1 decap_w0
xfeed_8671 0 1 decap_w0
xfeed_8670 0 1 decap_w0
xfeed_4369 0 1 tie
xfeed_4368 0 1 decap_w0
xfeed_4367 0 1 decap_w0
xfeed_4366 0 1 decap_w0
xfeed_4365 0 1 decap_w0
xfeed_4364 0 1 decap_w0
xfeed_4363 0 1 decap_w0
xfeed_4362 0 1 decap_w0
xfeed_4361 0 1 decap_w0
xfeed_4360 0 1 tie
xfeed_3838 0 1 decap_w0
xfeed_3837 0 1 decap_w0
xfeed_3836 0 1 decap_w0
xfeed_3835 0 1 decap_w0
xfeed_3834 0 1 decap_w0
xfeed_3833 0 1 decap_w0
xfeed_3832 0 1 decap_w0
xfeed_3831 0 1 decap_w0
xfeed_3830 0 1 decap_w0
xsubckt_510_and4_x1 0 1 241 319 265 261 242 and4_x1
xfeed_8679 0 1 decap_w0
xfeed_8678 0 1 decap_w0
xfeed_3839 0 1 decap_w0
xsubckt_1197_nand2_x0 0 1 1367 198 1368 nand2_x0
xsubckt_946_nand2_x0 0 1 1572 1941 1575 nand2_x0
xsubckt_941_and4_x1 0 1 1576 1917 680 673 670 and4_x1
xsubckt_123_and2_x1 0 1 645 660 646 and2_x1
xsubckt_1467_and3_x1 0 1 1129 537 458 1130 and3_x1
xfeed_10579 0 1 decap_w0
xfeed_10578 0 1 decap_w0
xfeed_10577 0 1 decap_w0
xfeed_10576 0 1 decap_w0
xfeed_10575 0 1 decap_w0
xfeed_10574 0 1 decap_w0
xfeed_10573 0 1 decap_w0
xfeed_10572 0 1 tie
xfeed_10571 0 1 decap_w0
xfeed_10570 0 1 decap_w0
xfeed_8684 0 1 decap_w0
xfeed_8683 0 1 decap_w0
xfeed_8682 0 1 decap_w0
xfeed_8681 0 1 decap_w0
xfeed_8680 0 1 tie
xfeed_4379 0 1 decap_w0
xfeed_4378 0 1 decap_w0
xfeed_4377 0 1 decap_w0
xfeed_4376 0 1 decap_w0
xfeed_4375 0 1 decap_w0
xfeed_4374 0 1 tie
xfeed_4373 0 1 decap_w0
xfeed_4372 0 1 decap_w0
xfeed_4371 0 1 decap_w0
xfeed_4370 0 1 decap_w0
xfeed_3845 0 1 tie
xfeed_3844 0 1 decap_w0
xfeed_3843 0 1 decap_w0
xfeed_3842 0 1 decap_w0
xfeed_3841 0 1 decap_w0
xfeed_3840 0 1 tie
xsubckt_1360_nand2_x0 0 1 1229 1967 1316 nand2_x0
xsubckt_1450_nand2_x0 0 1 1145 1917 1147 nand2_x0
xsubckt_1455_or21nand_x0 0 1 1141 1933 548 1744 or21nand_x0
xsubckt_1525_nor4_x0 0 1 1071 208 1082 1080 1079 nor4_x0
xfeed_8689 0 1 decap_w0
xfeed_8688 0 1 decap_w0
xfeed_8687 0 1 decap_w0
xfeed_8686 0 1 decap_w0
xfeed_8685 0 1 decap_w0
xfeed_3849 0 1 decap_w0
xfeed_3848 0 1 decap_w0
xfeed_3847 0 1 decap_w0
xfeed_3846 0 1 decap_w0
xsubckt_440_and3_x1 0 1 310 643 532 385 and3_x1
xfeed_10589 0 1 decap_w0
xfeed_10588 0 1 decap_w0
xfeed_10587 0 1 decap_w0
xfeed_10586 0 1 decap_w0
xfeed_10585 0 1 decap_w0
xfeed_10584 0 1 decap_w0
xfeed_10583 0 1 decap_w0
xfeed_10582 0 1 decap_w0
xfeed_10581 0 1 decap_w0
xfeed_10580 0 1 decap_w0
xfeed_9309 0 1 decap_w0
xfeed_9308 0 1 decap_w0
xfeed_9307 0 1 decap_w0
xfeed_9306 0 1 decap_w0
xfeed_9305 0 1 decap_w0
xfeed_9304 0 1 decap_w0
xfeed_9303 0 1 tie
xfeed_9302 0 1 decap_w0
xfeed_9301 0 1 decap_w0
xfeed_9300 0 1 decap_w0
xfeed_8691 0 1 decap_w0
xfeed_8690 0 1 decap_w0
xfeed_4389 0 1 decap_w0
xfeed_4388 0 1 decap_w0
xfeed_4387 0 1 decap_w0
xfeed_4386 0 1 decap_w0
xfeed_4385 0 1 decap_w0
xfeed_4384 0 1 decap_w0
xfeed_4383 0 1 decap_w0
xfeed_4382 0 1 decap_w0
xfeed_4381 0 1 decap_w0
xfeed_4380 0 1 decap_w0
xfeed_3852 0 1 tie
xfeed_3851 0 1 decap_w0
xfeed_3850 0 1 decap_w0
xsubckt_1573_nor2_x0 0 1 1021 1027 1022 nor2_x0
xfeed_11209 0 1 decap_w0
xfeed_11208 0 1 decap_w0
xfeed_11207 0 1 decap_w0
xfeed_11206 0 1 decap_w0
xfeed_11205 0 1 decap_w0
xfeed_11204 0 1 decap_w0
xfeed_11203 0 1 decap_w0
xfeed_11202 0 1 tie
xfeed_11201 0 1 decap_w0
xfeed_11200 0 1 decap_w0
xfeed_8699 0 1 decap_w0
xfeed_8698 0 1 decap_w0
xfeed_8697 0 1 tie
xfeed_8696 0 1 decap_w0
xfeed_8695 0 1 decap_w0
xfeed_8694 0 1 decap_w0
xfeed_8693 0 1 decap_w0
xfeed_8692 0 1 tie
xfeed_3859 0 1 decap_w0
xfeed_3858 0 1 decap_w0
xfeed_3856 0 1 decap_w0
xfeed_3855 0 1 decap_w0
xfeed_3854 0 1 decap_w0
xfeed_3853 0 1 decap_w0
xsubckt_835_nand3_x0 0 1 1642 2068 682 490 nand3_x0
xsubckt_318_nand2_x0 0 1 430 609 598 nand2_x0
xsubckt_273_xor2_x0 0 1 475 2055 1961 xor2_x0
xsubckt_228_nand2_x0 0 1 523 1986 1988 nand2_x0
xsubckt_462_and2_x1 0 1 288 609 581 and2_x1
xsubckt_1516_and21nor_x0 0 1 1080 737 547 1745 and21nor_x0
xfeed_10599 0 1 decap_w0
xfeed_10598 0 1 decap_w0
xfeed_10597 0 1 decap_w0
xfeed_10596 0 1 decap_w0
xfeed_10595 0 1 decap_w0
xfeed_10594 0 1 tie
xfeed_10593 0 1 decap_w0
xfeed_10592 0 1 decap_w0
xfeed_10591 0 1 decap_w0
xfeed_10590 0 1 tie
xfeed_9319 0 1 decap_w0
xfeed_9318 0 1 decap_w0
xfeed_9317 0 1 tie
xfeed_9316 0 1 decap_w0
xfeed_9315 0 1 decap_w0
xfeed_9314 0 1 decap_w0
xfeed_9313 0 1 decap_w0
xfeed_9312 0 1 decap_w0
xfeed_9311 0 1 decap_w0
xfeed_9310 0 1 tie
xfeed_5009 0 1 decap_w0
xfeed_5008 0 1 decap_w0
xfeed_5007 0 1 decap_w0
xfeed_5006 0 1 decap_w0
xfeed_5005 0 1 decap_w0
xfeed_5004 0 1 decap_w0
xfeed_5003 0 1 decap_w0
xfeed_5002 0 1 tie
xfeed_5001 0 1 decap_w0
xfeed_5000 0 1 decap_w0
xfeed_4398 0 1 decap_w0
xfeed_4397 0 1 decap_w0
xfeed_4396 0 1 decap_w0
xfeed_4395 0 1 decap_w0
xfeed_4394 0 1 tie
xfeed_4393 0 1 decap_w0
xfeed_4391 0 1 decap_w0
xfeed_4390 0 1 decap_w0
xsubckt_867_and3_x1 0 1 1615 2052 1962 1617 and3_x1
xsubckt_1425_nand4_x0 0 1 1168 1207 1196 1184 1171 nand4_x0
xsubckt_1439_nand2_x0 0 1 1800 1166 1156 nand2_x0
xfeed_11219 0 1 decap_w0
xfeed_11218 0 1 decap_w0
xfeed_11217 0 1 decap_w0
xfeed_11216 0 1 decap_w0
xfeed_11215 0 1 decap_w0
xfeed_11214 0 1 decap_w0
xfeed_11213 0 1 decap_w0
xfeed_11212 0 1 decap_w0
xfeed_11211 0 1 tie
xfeed_11210 0 1 decap_w0
xfeed_3869 0 1 decap_w0
xfeed_3868 0 1 decap_w0
xfeed_3867 0 1 decap_w0
xfeed_3866 0 1 decap_w0
xfeed_3865 0 1 decap_w0
xfeed_3864 0 1 decap_w0
xfeed_3863 0 1 decap_w0
xfeed_3862 0 1 decap_w0
xfeed_3861 0 1 decap_w0
xfeed_3860 0 1 decap_w0
xsubckt_876_nexor2_x0 0 1 1607 765 1611 nexor2_x0
xsubckt_701_and3_x1 0 1 1763 484 435 1764 and3_x1
xsubckt_1349_nand2_x0 0 1 1239 2053 479 nand2_x0
xsubckt_1755_or21nand_x0 0 1 839 879 845 843 or21nand_x0
xspare_buffer_0 0 1 82 83 buf_x4
xspare_buffer_3 0 1 22 23 buf_x4
xspare_buffer_4 0 1 81 82 buf_x4
xspare_buffer_7 0 1 21 22 buf_x4
xspare_buffer_8 0 1 68 82 buf_x4
xfeed_9329 0 1 decap_w0
xfeed_9328 0 1 decap_w0
xfeed_9327 0 1 decap_w0
xfeed_9326 0 1 decap_w0
xfeed_9325 0 1 decap_w0
xfeed_9324 0 1 tie
xfeed_9323 0 1 decap_w0
xfeed_9322 0 1 decap_w0
xfeed_9321 0 1 decap_w0
xfeed_9320 0 1 decap_w0
xfeed_5019 0 1 decap_w0
xfeed_5018 0 1 decap_w0
xfeed_5017 0 1 decap_w0
xfeed_5016 0 1 decap_w0
xfeed_5015 0 1 decap_w0
xfeed_5014 0 1 decap_w0
xfeed_5013 0 1 decap_w0
xfeed_5012 0 1 decap_w0
xfeed_5011 0 1 decap_w0
xfeed_5010 0 1 decap_w0
xsubckt_889_and2_x1 0 1 1597 1962 1598 and2_x1
xfeed_11229 0 1 decap_w0
xfeed_11228 0 1 tie
xfeed_11227 0 1 decap_w0
xfeed_11226 0 1 decap_w0
xfeed_11225 0 1 decap_w0
xfeed_11224 0 1 decap_w0
xfeed_11223 0 1 decap_w0
xfeed_11222 0 1 decap_w0
xfeed_11221 0 1 tie
xfeed_11220 0 1 decap_w0
xfeed_3879 0 1 decap_w0
xfeed_3878 0 1 decap_w0
xfeed_3877 0 1 decap_w0
xfeed_3876 0 1 decap_w0
xfeed_3875 0 1 decap_w0
xfeed_3874 0 1 tie
xfeed_3873 0 1 decap_w0
xfeed_3872 0 1 decap_w0
xfeed_3871 0 1 decap_w0
xfeed_3870 0 1 decap_w0
xsubckt_992_nand4_x0 0 1 1536 638 632 525 520 nand4_x0
xsubckt_937_mux2_x1 0 1 1881 438 1577 1983 mux2_x1
xsubckt_284_or21nand_x0 0 1 464 465 564 572 or21nand_x0
xsubckt_121_nand2_x0 0 1 647 785 2001 nand2_x0
xsubckt_1315_and21nor_x0 0 1 1270 750 478 1317 and21nor_x0
xsubckt_1332_nand2_x0 0 1 1254 1917 1255 nand2_x0
xsubckt_1416_or2_x1 0 1 1177 691 1323 or2_x1
xsubckt_1422_nand2_x0 0 1 1171 1178 1173 nand2_x0
xsubckt_1706_mux2_x1 0 1 888 928 890 1142 mux2_x1
xfeed_9339 0 1 decap_w0
xfeed_9338 0 1 tie
xfeed_9337 0 1 decap_w0
xfeed_9336 0 1 decap_w0
xfeed_9335 0 1 decap_w0
xfeed_9334 0 1 decap_w0
xfeed_9333 0 1 decap_w0
xfeed_9332 0 1 decap_w0
xfeed_9331 0 1 tie
xfeed_9330 0 1 decap_w0
xfeed_8809 0 1 decap_w0
xfeed_8808 0 1 decap_w0
xfeed_8807 0 1 decap_w0
xfeed_8806 0 1 decap_w0
xfeed_8805 0 1 decap_w0
xfeed_8804 0 1 decap_w0
xfeed_8803 0 1 decap_w0
xfeed_8802 0 1 decap_w0
xfeed_8801 0 1 decap_w0
xfeed_8800 0 1 decap_w0
xfeed_5029 0 1 decap_w0
xfeed_5028 0 1 decap_w0
xfeed_5027 0 1 decap_w0
xfeed_5026 0 1 decap_w0
xfeed_5025 0 1 decap_w0
xfeed_5024 0 1 decap_w0
xfeed_5023 0 1 decap_w0
xfeed_5022 0 1 decap_w0
xfeed_5021 0 1 decap_w0
xfeed_5020 0 1 decap_w0
xsubckt_738_nand2_x0 0 1 1727 1729 1728 nand2_x0
xsubckt_1418_nand3_x0 0 1 1175 2068 665 657 nand3_x0
xfeed_11239 0 1 decap_w0
xfeed_11238 0 1 decap_w0
xfeed_11237 0 1 decap_w0
xfeed_11236 0 1 decap_w0
xfeed_11235 0 1 decap_w0
xfeed_11234 0 1 decap_w0
xfeed_11233 0 1 decap_w0
xfeed_11232 0 1 decap_w0
xfeed_11231 0 1 decap_w0
xfeed_11230 0 1 decap_w0
xfeed_10700 0 1 decap_w0
xfeed_3889 0 1 decap_w0
xfeed_3888 0 1 tie
xfeed_3887 0 1 decap_w0
xfeed_3885 0 1 decap_w0
xfeed_3884 0 1 decap_w0
xfeed_3883 0 1 decap_w0
xfeed_3882 0 1 decap_w0
xfeed_3881 0 1 tie
xfeed_3880 0 1 decap_w0
xsubckt_53_inv_x0 0 1 729 1978 inv_x0
xsubckt_51_inv_x0 0 1 731 1979 inv_x0
xfeed_10709 0 1 decap_w0
xfeed_10708 0 1 decap_w0
xfeed_10707 0 1 decap_w0
xfeed_10706 0 1 decap_w0
xfeed_10705 0 1 decap_w0
xfeed_10704 0 1 decap_w0
xfeed_10703 0 1 decap_w0
xfeed_10702 0 1 decap_w0
xfeed_10701 0 1 decap_w0
xfeed_9348 0 1 decap_w0
xfeed_9347 0 1 decap_w0
xfeed_9346 0 1 decap_w0
xfeed_9345 0 1 decap_w0
xfeed_9344 0 1 decap_w0
xfeed_9343 0 1 tie
xfeed_9342 0 1 decap_w0
xfeed_9341 0 1 decap_w0
xfeed_9340 0 1 decap_w0
xfeed_8817 0 1 decap_w0
xfeed_8816 0 1 decap_w0
xfeed_8815 0 1 decap_w0
xfeed_8814 0 1 tie
xfeed_8813 0 1 decap_w0
xfeed_8812 0 1 decap_w0
xfeed_8811 0 1 decap_w0
xfeed_8810 0 1 decap_w0
xfeed_5039 0 1 decap_w0
xfeed_5038 0 1 decap_w0
xfeed_5037 0 1 decap_w0
xfeed_5036 0 1 decap_w0
xfeed_5035 0 1 decap_w0
xfeed_5034 0 1 decap_w0
xfeed_5033 0 1 decap_w0
xfeed_5032 0 1 decap_w0
xfeed_5031 0 1 decap_w0
xfeed_5030 0 1 tie
xfeed_4509 0 1 decap_w0
xfeed_4508 0 1 decap_w0
xfeed_4507 0 1 decap_w0
xfeed_4506 0 1 decap_w0
xfeed_4505 0 1 decap_w0
xfeed_4504 0 1 tie
xfeed_4503 0 1 decap_w0
xfeed_4502 0 1 decap_w0
xfeed_4501 0 1 decap_w0
xfeed_4500 0 1 decap_w0
xsubckt_230_mux2_x1 0 1 521 1988 1997 1986 mux2_x1
xsubckt_59_inv_x0 0 1 723 1933 inv_x0
xsubckt_57_inv_x0 0 1 725 1984 inv_x0
xsubckt_55_inv_x0 0 1 727 1976 inv_x0
xsubckt_454_nand4_x0 0 1 296 533 518 384 360 nand4_x0
xfeed_11246 0 1 decap_w0
xfeed_11245 0 1 decap_w0
xfeed_11244 0 1 decap_w0
xfeed_11243 0 1 decap_w0
xfeed_11242 0 1 decap_w0
xfeed_11241 0 1 decap_w0
xfeed_11240 0 1 tie
xfeed_8819 0 1 decap_w0
xfeed_8818 0 1 tie
xfeed_3898 0 1 decap_w0
xfeed_3897 0 1 decap_w0
xfeed_3896 0 1 decap_w0
xfeed_3895 0 1 decap_w0
xfeed_3894 0 1 decap_w0
xfeed_3892 0 1 decap_w0
xfeed_3891 0 1 decap_w0
xfeed_3890 0 1 decap_w0
xsubckt_763_nor3_x0 0 1 1705 1710 1709 1706 nor3_x0
xfeed_11249 0 1 decap_w0
xfeed_11248 0 1 decap_w0
xfeed_11247 0 1 decap_w0
xfeed_10719 0 1 decap_w0
xfeed_10718 0 1 decap_w0
xfeed_10717 0 1 decap_w0
xfeed_10716 0 1 decap_w0
xfeed_10715 0 1 decap_w0
xfeed_10714 0 1 decap_w0
xfeed_10713 0 1 decap_w0
xfeed_10712 0 1 decap_w0
xfeed_10711 0 1 decap_w0
xfeed_10710 0 1 decap_w0
xfeed_9359 0 1 decap_w0
xfeed_9358 0 1 decap_w0
xfeed_9357 0 1 decap_w0
xfeed_9356 0 1 decap_w0
xfeed_9354 0 1 decap_w0
xfeed_9353 0 1 tie
xfeed_9352 0 1 decap_w0
xfeed_9351 0 1 decap_w0
xfeed_9350 0 1 decap_w0
xfeed_8824 0 1 decap_w0
xfeed_8823 0 1 decap_w0
xfeed_8822 0 1 decap_w0
xfeed_8821 0 1 decap_w0
xfeed_8820 0 1 decap_w0
xfeed_5049 0 1 decap_w0
xfeed_5048 0 1 decap_w0
xfeed_5047 0 1 decap_w0
xfeed_5046 0 1 decap_w0
xfeed_5045 0 1 decap_w0
xfeed_5044 0 1 decap_w0
xfeed_5043 0 1 decap_w0
xfeed_5042 0 1 decap_w0
xfeed_5041 0 1 decap_w0
xfeed_5040 0 1 decap_w0
xfeed_4519 0 1 decap_w0
xfeed_4518 0 1 decap_w0
xfeed_4517 0 1 decap_w0
xfeed_4516 0 1 decap_w0
xfeed_4515 0 1 decap_w0
xfeed_4514 0 1 decap_w0
xfeed_4513 0 1 decap_w0
xfeed_4512 0 1 decap_w0
xfeed_4511 0 1 decap_w0
xfeed_4510 0 1 decap_w0
xsubckt_184_nand4_x0 0 1 574 714 1928 681 674 nand4_x0
xsubckt_451_nand2_x0 0 1 299 301 300 nand2_x0
xsubckt_509_and3_x1 0 1 242 259 256 243 and3_x1
xsubckt_1382_and2_x1 0 1 1208 1219 1210 and2_x1
xspare_feed_10 0 1 tie
xspare_feed_11 0 1 tie
xspare_feed_12 0 1 tie
xspare_feed_13 0 1 tie
xfeed_11253 0 1 tie
xfeed_11252 0 1 decap_w0
xfeed_11251 0 1 decap_w0
xfeed_11250 0 1 decap_w0
xfeed_8829 0 1 decap_w0
xfeed_8828 0 1 tie
xfeed_8827 0 1 decap_w0
xfeed_8826 0 1 decap_w0
xfeed_8825 0 1 decap_w0
xspare_feed_14 0 1 tie
xspare_feed_15 0 1 tie
xspare_feed_16 0 1 tie
xspare_feed_17 0 1 tie
xspare_feed_18 0 1 tie
xspare_feed_19 0 1 tie
xfeed_11259 0 1 decap_w0
xfeed_11258 0 1 decap_w0
xfeed_11257 0 1 decap_w0
xfeed_11256 0 1 decap_w0
xfeed_11255 0 1 decap_w0
xfeed_11254 0 1 decap_w0
xfeed_10729 0 1 decap_w0
xfeed_10728 0 1 tie
xfeed_10727 0 1 decap_w0
xfeed_10726 0 1 decap_w0
xfeed_10725 0 1 decap_w0
xfeed_10724 0 1 decap_w0
xfeed_10723 0 1 decap_w0
xfeed_10722 0 1 decap_w0
xfeed_10721 0 1 tie
xfeed_10720 0 1 decap_w0
xfeed_9369 0 1 decap_w0
xfeed_9368 0 1 decap_w0
xfeed_9367 0 1 decap_w0
xfeed_9366 0 1 decap_w0
xfeed_9365 0 1 tie
xfeed_9364 0 1 decap_w0
xfeed_9363 0 1 decap_w0
xfeed_9362 0 1 decap_w0
xfeed_9361 0 1 tie
xfeed_9360 0 1 decap_w0
xfeed_8831 0 1 decap_w0
xfeed_8830 0 1 decap_w0
xfeed_5059 0 1 decap_w0
xfeed_5058 0 1 decap_w0
xfeed_5057 0 1 decap_w0
xfeed_5056 0 1 decap_w0
xfeed_5055 0 1 decap_w0
xfeed_5054 0 1 decap_w0
xfeed_5053 0 1 decap_w0
xfeed_5052 0 1 decap_w0
xfeed_5051 0 1 decap_w0
xfeed_5050 0 1 decap_w0
xfeed_4529 0 1 decap_w0
xfeed_4528 0 1 decap_w0
xfeed_4527 0 1 decap_w0
xfeed_4526 0 1 decap_w0
xfeed_4525 0 1 decap_w0
xfeed_4524 0 1 tie
xfeed_4523 0 1 decap_w0
xfeed_4522 0 1 decap_w0
xfeed_4521 0 1 decap_w0
xfeed_4520 0 1 decap_w0
xsubckt_964_nand4_x0 0 1 1559 653 622 525 520 nand4_x0
xsubckt_271_nand2_x0 0 1 477 558 479 nand2_x0
xsubckt_134_mux2_x1 0 1 634 1993 2002 1986 mux2_x1
xspare_feed_20 0 1 tie
xfeed_11260 0 1 decap_w0
xfeed_8839 0 1 decap_w0
xfeed_8838 0 1 decap_w0
xfeed_8837 0 1 decap_w0
xfeed_8836 0 1 decap_w0
xfeed_8835 0 1 decap_w0
xfeed_8834 0 1 decap_w0
xfeed_8833 0 1 decap_w0
xfeed_8832 0 1 decap_w0
xsubckt_645_and21nor_x0 0 1 114 751 449 410 and21nor_x0
xsubckt_267_nand3_x0 0 1 481 687 609 489 nand3_x0
xspare_feed_21 0 1 tie
xspare_feed_22 0 1 tie
xspare_feed_23 0 1 tie
xspare_feed_24 0 1 tie
xspare_feed_25 0 1 tie
xspare_feed_26 0 1 tie
xspare_feed_27 0 1 tie
xspare_feed_28 0 1 tie
xspare_feed_29 0 1 tie
xfeed_11269 0 1 decap_w0
xfeed_11268 0 1 decap_w0
xfeed_11267 0 1 tie
xfeed_11266 0 1 decap_w0
xfeed_11265 0 1 decap_w0
xfeed_11264 0 1 decap_w0
xfeed_11263 0 1 decap_w0
xfeed_11262 0 1 decap_w0
xfeed_11261 0 1 decap_w0
xfeed_10739 0 1 decap_w0
xfeed_10738 0 1 decap_w0
xfeed_10737 0 1 decap_w0
xfeed_10736 0 1 decap_w0
xfeed_10735 0 1 decap_w0
xfeed_10734 0 1 decap_w0
xfeed_10733 0 1 decap_w0
xfeed_10732 0 1 decap_w0
xfeed_10731 0 1 decap_w0
xfeed_10730 0 1 decap_w0
xfeed_9376 0 1 decap_w0
xfeed_9375 0 1 decap_w0
xfeed_9374 0 1 decap_w0
xfeed_9373 0 1 decap_w0
xfeed_9372 0 1 decap_w0
xfeed_9371 0 1 decap_w0
xfeed_9370 0 1 decap_w0
xfeed_5069 0 1 decap_w0
xfeed_5068 0 1 decap_w0
xfeed_5067 0 1 decap_w0
xfeed_5066 0 1 decap_w0
xfeed_5065 0 1 decap_w0
xfeed_5064 0 1 decap_w0
xfeed_5063 0 1 decap_w0
xfeed_5062 0 1 decap_w0
xfeed_5061 0 1 decap_w0
xfeed_5060 0 1 decap_w0
xfeed_4538 0 1 decap_w0
xfeed_4537 0 1 decap_w0
xfeed_4536 0 1 decap_w0
xfeed_4535 0 1 decap_w0
xfeed_4534 0 1 decap_w0
xfeed_4532 0 1 decap_w0
xfeed_4531 0 1 decap_w0
xfeed_4530 0 1 decap_w0
xsubckt_961_nand2_x0 0 1 1561 1936 1575 nand2_x0
xsubckt_922_mux2_x1 0 1 1894 1600 2034 1579 mux2_x1
xsubckt_784_or21nand_x0 0 1 1687 2058 1742 1740 or21nand_x0
xsubckt_1526_or4_x1 0 1 1067 208 1082 1080 1079 or4_x1
xspare_feed_0 0 1 tie
xspare_feed_1 0 1 tie
xspare_feed_2 0 1 tie
xspare_feed_3 0 1 tie
xspare_feed_4 0 1 tie
xspare_feed_5 0 1 tie
xspare_feed_6 0 1 tie
xspare_feed_7 0 1 tie
xspare_feed_8 0 1 tie
xspare_feed_9 0 1 tie
xfeed_9379 0 1 decap_w0
xfeed_9378 0 1 tie
xfeed_8849 0 1 decap_w0
xfeed_8848 0 1 decap_w0
xfeed_8847 0 1 decap_w0
xfeed_8846 0 1 decap_w0
xfeed_8845 0 1 decap_w0
xfeed_8843 0 1 decap_w0
xfeed_8842 0 1 decap_w0
xfeed_8841 0 1 decap_w0
xfeed_8840 0 1 decap_w0
xsubckt_1168_and3_x1 0 1 1394 1934 608 603 and3_x1
xsubckt_1052_or21nand_x0 0 1 1854 1489 1490 1491 or21nand_x0
xsubckt_1551_nand3_x0 0 1 1043 1103 1050 1048 nand3_x0
xsubckt_1577_and4_x1 0 1 1017 1998 1128 1098 1097 and4_x1
xspare_feed_30 0 1 tie
xspare_feed_31 0 1 tie
xspare_feed_32 0 1 tie
xspare_feed_33 0 1 tie
xspare_feed_34 0 1 tie
xspare_feed_35 0 1 tie
xspare_feed_36 0 1 tie
xspare_feed_37 0 1 tie
xspare_feed_38 0 1 tie
xspare_feed_39 0 1 tie
xfeed_11279 0 1 decap_w0
xfeed_11277 0 1 decap_w0
xfeed_11276 0 1 decap_w0
xfeed_11275 0 1 decap_w0
xfeed_11274 0 1 decap_w0
xfeed_11273 0 1 decap_w0
xfeed_11272 0 1 decap_w0
xfeed_11271 0 1 decap_w0
xfeed_11270 0 1 decap_w0
xfeed_10749 0 1 decap_w0
xfeed_10748 0 1 decap_w0
xfeed_10747 0 1 decap_w0
xfeed_10746 0 1 decap_w0
xfeed_10745 0 1 decap_w0
xfeed_10744 0 1 decap_w0
xfeed_10743 0 1 decap_w0
xfeed_10742 0 1 decap_w0
xfeed_10741 0 1 decap_w0
xfeed_10740 0 1 decap_w0
xfeed_9384 0 1 decap_w0
xfeed_9383 0 1 decap_w0
xfeed_9382 0 1 decap_w0
xfeed_9381 0 1 decap_w0
xfeed_9380 0 1 decap_w0
xfeed_5079 0 1 decap_w0
xfeed_5078 0 1 decap_w0
xfeed_5077 0 1 decap_w0
xfeed_5076 0 1 decap_w0
xfeed_5075 0 1 decap_w0
xfeed_5074 0 1 decap_w0
xfeed_5073 0 1 decap_w0
xfeed_5072 0 1 decap_w0
xfeed_5071 0 1 decap_w0
xfeed_5070 0 1 decap_w0
xfeed_4545 0 1 decap_w0
xfeed_4544 0 1 tie
xfeed_4543 0 1 decap_w0
xfeed_4542 0 1 decap_w0
xfeed_4541 0 1 decap_w0
xsubckt_1242_mux2_x1 0 1 1819 2103 2070 1334 mux2_x1
xsubckt_1002_and3_x1 0 1 1527 652 623 520 and3_x1
xfeed_9389 0 1 decap_w0
xfeed_9388 0 1 decap_w0
xfeed_9387 0 1 tie
xfeed_9386 0 1 decap_w0
xfeed_9385 0 1 decap_w0
xfeed_8859 0 1 decap_w0
xfeed_8858 0 1 decap_w0
xfeed_8857 0 1 decap_w0
xfeed_8856 0 1 decap_w0
xfeed_8855 0 1 decap_w0
xfeed_8854 0 1 decap_w0
xfeed_8853 0 1 decap_w0
xfeed_8852 0 1 decap_w0
xfeed_8851 0 1 decap_w0
xfeed_8850 0 1 decap_w0
xfeed_4549 0 1 decap_w0
xfeed_4548 0 1 decap_w0
xfeed_4547 0 1 decap_w0
xfeed_4546 0 1 decap_w0
xsubckt_1514_and21nor_x0 0 1 1082 736 547 1745 and21nor_x0
xspare_feed_40 0 1 tie
xspare_feed_41 0 1 tie
xspare_feed_42 0 1 tie
xspare_feed_43 0 1 tie
xspare_feed_44 0 1 tie
xspare_feed_45 0 1 tie
xspare_feed_46 0 1 tie
xspare_feed_47 0 1 tie
xspare_feed_48 0 1 tie
xspare_feed_49 0 1 tie
xfeed_11289 0 1 decap_w0
xfeed_11288 0 1 tie
xfeed_11287 0 1 decap_w0
xfeed_11286 0 1 decap_w0
xfeed_11285 0 1 decap_w0
xfeed_11284 0 1 decap_w0
xfeed_11283 0 1 decap_w0
xfeed_11282 0 1 decap_w0
xfeed_11281 0 1 decap_w0
xfeed_11280 0 1 decap_w0
xfeed_10759 0 1 decap_w0
xfeed_10758 0 1 decap_w0
xfeed_10757 0 1 decap_w0
xfeed_10756 0 1 decap_w0
xfeed_10755 0 1 decap_w0
xfeed_10754 0 1 tie
xfeed_10753 0 1 decap_w0
xfeed_10752 0 1 decap_w0
xfeed_10751 0 1 decap_w0
xfeed_10750 0 1 decap_w0
xfeed_9391 0 1 decap_w0
xfeed_9390 0 1 decap_w0
xfeed_5089 0 1 decap_w0
xfeed_5088 0 1 decap_w0
xfeed_5087 0 1 tie
xfeed_5086 0 1 decap_w0
xfeed_5085 0 1 decap_w0
xfeed_5084 0 1 decap_w0
xfeed_5083 0 1 decap_w0
xfeed_5082 0 1 decap_w0
xfeed_5081 0 1 decap_w0
xfeed_5080 0 1 decap_w0
xfeed_4552 0 1 decap_w0
xfeed_4551 0 1 decap_w0
xfeed_4550 0 1 decap_w0
xsubckt_1238_mux2_x1 0 1 1823 2093 2058 1334 mux2_x1
xsubckt_419_nand3_x0 0 1 330 687 680 421 nand3_x0
xsubckt_444_and21nor_x0 0 1 306 663 649 645 and21nor_x0
xsubckt_550_and4_x1 0 1 204 716 1924 1926 599 and4_x1
xsubckt_1547_and2_x1 0 1 1047 1050 1048 and2_x1
xsubckt_1673_mux2_x1 0 1 921 1103 1105 925 mux2_x1
xfeed_9399 0 1 decap_w0
xfeed_9398 0 1 decap_w0
xfeed_9397 0 1 decap_w0
xfeed_9396 0 1 decap_w0
xfeed_9395 0 1 decap_w0
xfeed_9394 0 1 tie
xfeed_9393 0 1 decap_w0
xfeed_9392 0 1 decap_w0
xfeed_8869 0 1 decap_w0
xfeed_8868 0 1 decap_w0
xfeed_8867 0 1 decap_w0
xfeed_8866 0 1 decap_w0
xfeed_8865 0 1 decap_w0
xfeed_8864 0 1 decap_w0
xfeed_8863 0 1 decap_w0
xfeed_8862 0 1 decap_w0
xfeed_8861 0 1 decap_w0
xfeed_8860 0 1 decap_w0
xfeed_4559 0 1 decap_w0
xfeed_4558 0 1 decap_w0
xfeed_4557 0 1 decap_w0
xfeed_4556 0 1 decap_w0
xfeed_4555 0 1 decap_w0
xfeed_4554 0 1 decap_w0
xfeed_4553 0 1 decap_w0
xsubckt_1009_nand4_x0 0 1 1520 643 533 519 1523 nand4_x0
xsubckt_329_nand3_x0 0 1 419 617 557 421 nand3_x0
xspare_feed_50 0 1 tie
xspare_feed_51 0 1 tie
xspare_feed_52 0 1 tie
xspare_feed_53 0 1 tie
xspare_feed_54 0 1 tie
xspare_feed_55 0 1 tie
xspare_feed_56 0 1 tie
xspare_feed_57 0 1 tie
xspare_feed_58 0 1 tie
xspare_feed_59 0 1 tie
xfeed_11299 0 1 decap_w0
xfeed_11298 0 1 tie
xfeed_11297 0 1 decap_w0
xfeed_11296 0 1 decap_w0
xfeed_11295 0 1 decap_w0
xfeed_11294 0 1 decap_w0
xfeed_11293 0 1 tie
xfeed_11292 0 1 decap_w0
xfeed_11291 0 1 decap_w0
xfeed_11290 0 1 decap_w0
xfeed_10769 0 1 decap_w0
xfeed_10768 0 1 decap_w0
xfeed_10767 0 1 decap_w0
xfeed_10766 0 1 tie
xfeed_10765 0 1 decap_w0
xfeed_10764 0 1 decap_w0
xfeed_10763 0 1 decap_w0
xfeed_10762 0 1 decap_w0
xfeed_10761 0 1 tie
xfeed_10760 0 1 decap_w0
xfeed_5098 0 1 decap_w0
xfeed_5097 0 1 decap_w0
xfeed_5096 0 1 decap_w0
xfeed_5095 0 1 decap_w0
xfeed_5094 0 1 decap_w0
xfeed_5093 0 1 decap_w0
xfeed_5092 0 1 decap_w0
xfeed_5091 0 1 decap_w0
xfeed_5090 0 1 decap_w0
xsubckt_1097_nand4_x0 0 1 1450 659 624 529 528 nand4_x0
xsubckt_544_and21nor_x0 0 1 210 408 447 712 and21nor_x0
xfeed_8879 0 1 tie
xfeed_8878 0 1 decap_w0
xfeed_8877 0 1 decap_w0
xfeed_8876 0 1 decap_w0
xfeed_8875 0 1 decap_w0
xfeed_8874 0 1 decap_w0
xfeed_8873 0 1 decap_w0
xfeed_8872 0 1 decap_w0
xfeed_8871 0 1 decap_w0
xfeed_8870 0 1 decap_w0
xfeed_5099 0 1 decap_w0
xfeed_4569 0 1 decap_w0
xfeed_4567 0 1 decap_w0
xfeed_4566 0 1 decap_w0
xfeed_4565 0 1 decap_w0
xfeed_4564 0 1 decap_w0
xfeed_4563 0 1 decap_w0
xfeed_4562 0 1 decap_w0
xfeed_4561 0 1 decap_w0
xfeed_4560 0 1 decap_w0
xspare_feed_60 0 1 tie
xspare_feed_61 0 1 tie
xspare_feed_62 0 1 tie
xspare_feed_63 0 1 tie
xspare_feed_64 0 1 tie
xspare_feed_65 0 1 tie
xspare_feed_66 0 1 tie
xspare_feed_67 0 1 tie
xspare_feed_68 0 1 tie
xspare_feed_69 0 1 tie
xfeed_10779 0 1 decap_w0
xfeed_10778 0 1 decap_w0
xfeed_10777 0 1 decap_w0
xfeed_10776 0 1 decap_w0
xfeed_10775 0 1 decap_w0
xfeed_10774 0 1 decap_w0
xfeed_10773 0 1 decap_w0
xfeed_10772 0 1 decap_w0
xfeed_10771 0 1 tie
xfeed_10770 0 1 decap_w0
xsubckt_576_nand4_x0 0 1 179 709 195 194 189 nand4_x0
xcmpt_abc_11867_new_n333_hfns_0 0 1 775 772 buf_x4
xcmpt_abc_11867_new_n333_hfns_1 0 1 774 772 buf_x4
xcmpt_abc_11867_new_n333_hfns_2 0 1 773 772 buf_x4
xcmpt_abc_11867_new_n333_hfns_3 0 1 772 776 buf_x4
xfeed_8889 0 1 decap_w0
xfeed_8888 0 1 decap_w0
xfeed_8887 0 1 decap_w0
xfeed_8886 0 1 tie
xfeed_8885 0 1 decap_w0
xfeed_8884 0 1 decap_w0
xfeed_8883 0 1 decap_w0
xfeed_8882 0 1 decap_w0
xfeed_8881 0 1 decap_w0
xfeed_8880 0 1 decap_w0
xfeed_4579 0 1 decap_w0
xfeed_4576 0 1 decap_w0
xfeed_4575 0 1 decap_w0
xfeed_4574 0 1 decap_w0
xfeed_4573 0 1 decap_w0
xfeed_4572 0 1 decap_w0
xfeed_4571 0 1 decap_w0
xfeed_4570 0 1 decap_w0
xsubckt_753_nand2_x0 0 1 1714 2000 1746 nand2_x0
xsubckt_476_and3_x1 0 1 274 277 276 275 and3_x1
xsubckt_1535_nor2_x0 0 1 1059 90 1122 nor2_x0
xsubckt_1649_or21nand_x0 0 1 945 1067 957 1072 or21nand_x0
xspare_feed_70 0 1 tie
xspare_feed_71 0 1 tie
xspare_feed_72 0 1 tie
xspare_feed_73 0 1 tie
xspare_feed_74 0 1 tie
xspare_feed_75 0 1 tie
xspare_feed_76 0 1 tie
xspare_feed_77 0 1 tie
xspare_feed_78 0 1 tie
xspare_feed_79 0 1 tie
xfeed_10789 0 1 decap_w0
xfeed_10788 0 1 decap_w0
xfeed_10787 0 1 decap_w0
xfeed_10786 0 1 decap_w0
xfeed_10785 0 1 decap_w0
xfeed_10784 0 1 decap_w0
xfeed_10783 0 1 decap_w0
xfeed_10782 0 1 decap_w0
xfeed_10781 0 1 decap_w0
xfeed_10780 0 1 decap_w0
xfeed_9509 0 1 decap_w0
xfeed_9508 0 1 decap_w0
xfeed_9507 0 1 decap_w0
xfeed_9506 0 1 decap_w0
xfeed_9505 0 1 decap_w0
xfeed_9504 0 1 decap_w0
xfeed_9503 0 1 decap_w0
xfeed_9502 0 1 decap_w0
xfeed_9501 0 1 decap_w0
xfeed_9500 0 1 decap_w0
xsubckt_1012_and21nor_x0 0 1 1865 1533 1519 1518 and21nor_x0
xsubckt_837_or4_x1 0 1 1640 1645 1644 1643 1641 or4_x1
xsubckt_674_nor2_x0 0 1 87 727 212 nor2_x0
xsubckt_1821_dff_x1 0 1 2019 1911 32 dff_x1
xsubckt_1823_dff_x1 0 1 2017 1909 35 dff_x1
xsubckt_1825_dff_x1 0 1 2015 1907 32 dff_x1
xfeed_11400 0 1 decap_w0
xfeed_8899 0 1 decap_w0
xfeed_8898 0 1 decap_w0
xfeed_8896 0 1 tie
xfeed_8895 0 1 decap_w0
xfeed_8894 0 1 decap_w0
xfeed_8893 0 1 decap_w0
xfeed_8892 0 1 decap_w0
xfeed_8890 0 1 decap_w0
xfeed_4589 0 1 decap_w0
xfeed_4588 0 1 decap_w0
xfeed_4587 0 1 decap_w0
xfeed_4586 0 1 decap_w0
xfeed_4585 0 1 decap_w0
xfeed_4584 0 1 decap_w0
xfeed_4583 0 1 decap_w0
xfeed_4582 0 1 decap_w0
xfeed_4581 0 1 decap_w0
xfeed_4580 0 1 decap_w0
xsubckt_1151_or21nand_x0 0 1 1409 1410 175 724 or21nand_x0
xsubckt_855_and2_x1 0 1 1786 2012 1963 and2_x1
xsubckt_844_and21nor_x0 0 1 1634 741 600 1745 and21nor_x0
xsubckt_1827_dff_x1 0 1 1930 29 74 dff_x1
xsubckt_1829_dff_x1 0 1 1928 27 74 dff_x1
xspare_feed_80 0 1 tie
xspare_feed_81 0 1 tie
xspare_feed_82 0 1 tie
xspare_feed_83 0 1 tie
xspare_feed_85 0 1 tie
xspare_feed_86 0 1 tie
xspare_feed_87 0 1 decap_w0
xspare_feed_88 0 1 tie
xspare_feed_89 0 1 tie
xfeed_11409 0 1 decap_w0
xfeed_11408 0 1 decap_w0
xfeed_11407 0 1 decap_w0
xfeed_11406 0 1 decap_w0
xfeed_11405 0 1 tie
xfeed_11404 0 1 decap_w0
xfeed_11403 0 1 decap_w0
xfeed_11402 0 1 decap_w0
xfeed_11401 0 1 decap_w0
xfeed_10799 0 1 decap_w0
xfeed_10798 0 1 decap_w0
xfeed_10797 0 1 tie
xfeed_10796 0 1 decap_w0
xfeed_10795 0 1 decap_w0
xfeed_10794 0 1 decap_w0
xfeed_10793 0 1 decap_w0
xfeed_10792 0 1 tie
xfeed_10791 0 1 decap_w0
xfeed_10790 0 1 decap_w0
xfeed_9517 0 1 decap_w0
xfeed_9516 0 1 decap_w0
xfeed_9515 0 1 decap_w0
xfeed_9514 0 1 tie
xfeed_9513 0 1 decap_w0
xfeed_9512 0 1 decap_w0
xfeed_9511 0 1 decap_w0
xfeed_9510 0 1 decap_w0
xfeed_5209 0 1 decap_w0
xfeed_5208 0 1 decap_w0
xfeed_5207 0 1 decap_w0
xfeed_5206 0 1 decap_w0
xfeed_5205 0 1 decap_w0
xfeed_5204 0 1 decap_w0
xfeed_5203 0 1 decap_w0
xfeed_5202 0 1 decap_w0
xfeed_5201 0 1 decap_w0
xfeed_5200 0 1 decap_w0
xsubckt_1101_and2_x1 0 1 1446 1449 1447 and2_x1
xsubckt_140_or2_x1 0 1 628 653 629 or2_x1
xfeed_9519 0 1 decap_w0
xfeed_9518 0 1 decap_w0
xfeed_4599 0 1 decap_w0
xfeed_4598 0 1 decap_w0
xfeed_4597 0 1 decap_w0
xfeed_4596 0 1 decap_w0
xfeed_4595 0 1 decap_w0
xfeed_4594 0 1 decap_w0
xfeed_4593 0 1 decap_w0
xfeed_4592 0 1 decap_w0
xfeed_4591 0 1 decap_w0
xfeed_4590 0 1 decap_w0
xsubckt_977_mux2_x1 0 1 1868 1551 1960 1576 mux2_x1
xsubckt_240_and2_x1 0 1 511 515 512 and2_x1
xsubckt_1426_nand2_x0 0 1 1167 1917 1168 nand2_x0
xsubckt_1613_and21nor_x0 0 1 981 1102 984 983 and21nor_x0
xspare_feed_90 0 1 decap_w0
xspare_feed_91 0 1 tie
xspare_feed_92 0 1 tie
xspare_feed_93 0 1 decap_w0
xspare_feed_94 0 1 tie
xspare_feed_95 0 1 tie
xspare_feed_96 0 1 decap_w0
xspare_feed_97 0 1 tie
xspare_feed_98 0 1 tie
xspare_feed_99 0 1 decap_w0
xfeed_11419 0 1 decap_w0
xfeed_11418 0 1 decap_w0
xfeed_11417 0 1 tie
xfeed_11416 0 1 decap_w0
xfeed_11415 0 1 decap_w0
xfeed_11414 0 1 decap_w0
xfeed_11413 0 1 decap_w0
xfeed_11412 0 1 decap_w0
xfeed_11411 0 1 decap_w0
xfeed_11410 0 1 decap_w0
xfeed_9524 0 1 decap_w0
xfeed_9523 0 1 decap_w0
xfeed_9522 0 1 decap_w0
xfeed_9521 0 1 decap_w0
xfeed_9520 0 1 decap_w0
xfeed_5219 0 1 decap_w0
xfeed_5217 0 1 tie
xfeed_5216 0 1 decap_w0
xfeed_5215 0 1 decap_w0
xfeed_5214 0 1 decap_w0
xfeed_5213 0 1 decap_w0
xfeed_5212 0 1 decap_w0
xfeed_5211 0 1 decap_w0
xfeed_5210 0 1 tie
xsubckt_1047_or21nand_x0 0 1 1855 1494 1493 1502 or21nand_x0
xsubckt_779_or21nand_x0 0 1 1691 1693 1767 90 or21nand_x0
xsubckt_288_and3_x1 0 1 460 1929 715 599 and3_x1
xsubckt_552_nand3_x0 0 1 202 592 573 203 nand3_x0
xsubckt_1448_or21nand_x0 0 1 1147 1149 1160 1168 or21nand_x0
xsubckt_1752_or21nand_x0 0 1 842 887 886 883 or21nand_x0
xfeed_9529 0 1 decap_w0
xfeed_9528 0 1 decap_w0
xfeed_9527 0 1 tie
xfeed_9526 0 1 decap_w0
xfeed_9525 0 1 decap_w0
xsubckt_1083_and2_x1 0 1 1462 707 1575 and2_x1
xsubckt_1005_and2_x1 0 1 1524 1526 1525 and2_x1
xsubckt_885_mux2_x1 0 1 1910 2018 1600 1619 mux2_x1
xsubckt_759_and2_x1 0 1 1709 2049 1748 and2_x1
xsubckt_60_inv_x0 0 1 722 2004 inv_x0
xfeed_11429 0 1 decap_w0
xfeed_11428 0 1 decap_w0
xfeed_11427 0 1 decap_w0
xfeed_11426 0 1 tie
xfeed_11425 0 1 decap_w0
xfeed_11424 0 1 decap_w0
xfeed_11423 0 1 decap_w0
xfeed_11422 0 1 decap_w0
xfeed_11421 0 1 tie
xfeed_11420 0 1 decap_w0
xfeed_9531 0 1 decap_w0
xfeed_9530 0 1 decap_w0
xfeed_5229 0 1 decap_w0
xfeed_5228 0 1 decap_w0
xfeed_5227 0 1 decap_w0
xfeed_5226 0 1 decap_w0
xfeed_5225 0 1 decap_w0
xfeed_5224 0 1 decap_w0
xfeed_5223 0 1 decap_w0
xfeed_5222 0 1 decap_w0
xfeed_5221 0 1 decap_w0
xfeed_5220 0 1 decap_w0
xsubckt_66_inv_x0 0 1 716 1929 inv_x0
xsubckt_64_inv_x0 0 1 718 2006 inv_x0
xsubckt_62_inv_x0 0 1 720 2005 inv_x0
xsubckt_478_or21nand_x0 0 1 272 273 282 353 or21nand_x0
xsubckt_1389_or2_x1 0 1 1202 693 1323 or2_x1
xsubckt_1583_nand3_x0 0 1 1011 1103 1018 1016 nand3_x0
xfeed_9539 0 1 decap_w0
xfeed_9538 0 1 decap_w0
xfeed_9537 0 1 decap_w0
xfeed_9536 0 1 decap_w0
xfeed_9535 0 1 decap_w0
xfeed_9534 0 1 decap_w0
xfeed_9533 0 1 decap_w0
xfeed_9532 0 1 tie
xsubckt_1108_and21nor_x0 0 1 1440 775 503 430 and21nor_x0
xsubckt_68_inv_x0 0 1 714 1927 inv_x0
xsubckt_527_and4_x1 0 1 225 332 249 228 226 and4_x1
xsubckt_1451_or21nand_x0 0 1 1799 1155 1146 1145 or21nand_x0
xfeed_11439 0 1 decap_w0
xfeed_11438 0 1 decap_w0
xfeed_11437 0 1 decap_w0
xfeed_11436 0 1 decap_w0
xfeed_11435 0 1 decap_w0
xfeed_11434 0 1 decap_w0
xfeed_11433 0 1 decap_w0
xfeed_11432 0 1 decap_w0
xfeed_11431 0 1 decap_w0
xfeed_11430 0 1 decap_w0
xfeed_10909 0 1 decap_w0
xfeed_10908 0 1 decap_w0
xfeed_10907 0 1 decap_w0
xfeed_10906 0 1 decap_w0
xfeed_10905 0 1 decap_w0
xfeed_10904 0 1 decap_w0
xfeed_10903 0 1 decap_w0
xfeed_10902 0 1 decap_w0
xfeed_10901 0 1 decap_w0
xfeed_10900 0 1 decap_w0
xfeed_5238 0 1 decap_w0
xfeed_5237 0 1 decap_w0
xfeed_5236 0 1 decap_w0
xfeed_5235 0 1 decap_w0
xfeed_5234 0 1 decap_w0
xfeed_5233 0 1 decap_w0
xfeed_5232 0 1 tie
xfeed_5231 0 1 decap_w0
xfeed_5230 0 1 decap_w0
xsubckt_1225_nand3_x0 0 1 1339 714 613 609 nand3_x0
xsubckt_455_nand2_x0 0 1 295 524 383 nand2_x0
xsubckt_1609_and21nor_x0 0 1 985 1104 989 987 and21nor_x0
xfeed_9549 0 1 decap_w0
xfeed_9548 0 1 decap_w0
xfeed_9547 0 1 decap_w0
xfeed_9546 0 1 decap_w0
xfeed_9545 0 1 decap_w0
xfeed_9544 0 1 tie
xfeed_9543 0 1 decap_w0
xfeed_9542 0 1 decap_w0
xfeed_9541 0 1 decap_w0
xfeed_9540 0 1 decap_w0
xfeed_5239 0 1 decap_w0
xfeed_4709 0 1 decap_w0
xfeed_4708 0 1 decap_w0
xfeed_4707 0 1 decap_w0
xfeed_4706 0 1 tie
xfeed_4705 0 1 decap_w0
xfeed_4704 0 1 decap_w0
xfeed_4703 0 1 decap_w0
xfeed_4702 0 1 decap_w0
xfeed_4701 0 1 decap_w0
xfeed_4700 0 1 decap_w0
xsubckt_972_nand3_x0 0 1 1553 623 519 1567 nand3_x0
xsubckt_100_mux2_x1 0 1 689 722 721 774 mux2_x1
xsubckt_1558_mux2_x1 0 1 1036 1110 1038 1142 mux2_x1
xfeed_11449 0 1 decap_w0
xfeed_11448 0 1 decap_w0
xfeed_11447 0 1 decap_w0
xfeed_11446 0 1 decap_w0
xfeed_11445 0 1 decap_w0
xfeed_11444 0 1 decap_w0
xfeed_11443 0 1 decap_w0
xfeed_11442 0 1 decap_w0
xfeed_11441 0 1 decap_w0
xfeed_11440 0 1 decap_w0
xfeed_10919 0 1 decap_w0
xfeed_10918 0 1 decap_w0
xfeed_10917 0 1 decap_w0
xfeed_10916 0 1 tie
xfeed_10915 0 1 decap_w0
xfeed_10914 0 1 decap_w0
xfeed_10913 0 1 decap_w0
xfeed_10912 0 1 decap_w0
xfeed_10911 0 1 decap_w0
xfeed_10910 0 1 decap_w0
xfeed_5245 0 1 decap_w0
xfeed_5244 0 1 decap_w0
xfeed_5243 0 1 decap_w0
xfeed_5242 0 1 tie
xfeed_5241 0 1 decap_w0
xfeed_5240 0 1 decap_w0
xsubckt_678_or21nand_x0 0 1 2076 1785 90 206 or21nand_x0
xsubckt_261_nand4_x0 0 1 487 1929 715 714 1928 nand4_x0
xfeed_9559 0 1 decap_w0
xfeed_9558 0 1 decap_w0
xfeed_9557 0 1 decap_w0
xfeed_9556 0 1 decap_w0
xfeed_9555 0 1 decap_w0
xfeed_9554 0 1 decap_w0
xfeed_9553 0 1 decap_w0
xfeed_9552 0 1 decap_w0
xfeed_9551 0 1 decap_w0
xfeed_9550 0 1 decap_w0
xfeed_5249 0 1 tie
xfeed_5248 0 1 decap_w0
xfeed_5247 0 1 decap_w0
xfeed_5246 0 1 decap_w0
xfeed_4719 0 1 decap_w0
xfeed_4718 0 1 decap_w0
xfeed_4717 0 1 decap_w0
xfeed_4716 0 1 decap_w0
xfeed_4715 0 1 decap_w0
xfeed_4714 0 1 decap_w0
xfeed_4713 0 1 decap_w0
xfeed_4712 0 1 tie
xfeed_4711 0 1 decap_w0
xfeed_4710 0 1 decap_w0
xsubckt_1252_and2_x1 0 1 1328 456 438 and2_x1
xsubckt_1396_nand2_x0 0 1 1195 1207 1196 nand2_x0
xfeed_11459 0 1 decap_w0
xfeed_11458 0 1 decap_w0
xfeed_11457 0 1 decap_w0
xfeed_11456 0 1 decap_w0
xfeed_11455 0 1 decap_w0
xfeed_11454 0 1 decap_w0
xfeed_11453 0 1 decap_w0
xfeed_11452 0 1 decap_w0
xfeed_11451 0 1 decap_w0
xfeed_11450 0 1 decap_w0
xfeed_10929 0 1 decap_w0
xfeed_10928 0 1 decap_w0
xfeed_10927 0 1 decap_w0
xfeed_10926 0 1 decap_w0
xfeed_10925 0 1 decap_w0
xfeed_10924 0 1 decap_w0
xfeed_10923 0 1 decap_w0
xfeed_10922 0 1 decap_w0
xfeed_10921 0 1 decap_w0
xfeed_10920 0 1 decap_w0
xfeed_5252 0 1 decap_w0
xfeed_5251 0 1 decap_w0
xfeed_5250 0 1 tie
xsubckt_1248_and2_x1 0 1 1332 314 1756 and2_x1
xsubckt_1186_and4_x1 0 1 1378 574 417 404 196 and4_x1
xsubckt_434_nand3_x0 0 1 316 617 581 557 nand3_x0
xsubckt_542_and21nor_x0 0 1 212 408 447 616 and21nor_x0
xfeed_9569 0 1 decap_w0
xfeed_9568 0 1 decap_w0
xfeed_9567 0 1 decap_w0
xfeed_9566 0 1 decap_w0
xfeed_9565 0 1 decap_w0
xfeed_9564 0 1 decap_w0
xfeed_9563 0 1 decap_w0
xfeed_9562 0 1 decap_w0
xfeed_9561 0 1 decap_w0
xfeed_9560 0 1 decap_w0
xfeed_5259 0 1 decap_w0
xfeed_5258 0 1 decap_w0
xfeed_5257 0 1 decap_w0
xfeed_5256 0 1 decap_w0
xfeed_5255 0 1 decap_w0
xfeed_5254 0 1 decap_w0
xfeed_5253 0 1 decap_w0
xfeed_4729 0 1 decap_w0
xfeed_4728 0 1 decap_w0
xfeed_4727 0 1 decap_w0
xfeed_4726 0 1 decap_w0
xfeed_4725 0 1 decap_w0
xfeed_4724 0 1 tie
xfeed_4723 0 1 decap_w0
xfeed_4722 0 1 decap_w0
xfeed_4721 0 1 decap_w0
xfeed_4720 0 1 decap_w0
xsubckt_1046_or21nand_x0 0 1 1493 1576 520 622 or21nand_x0
xsubckt_875_nand2_x0 0 1 1608 765 1610 nand2_x0
xsubckt_254_nand3_x0 0 1 497 679 571 557 nand3_x0
xsubckt_1731_mux2_x1 0 1 863 867 865 875 mux2_x1
xfeed_11469 0 1 decap_w0
xfeed_11468 0 1 decap_w0
xfeed_11467 0 1 decap_w0
xfeed_11466 0 1 decap_w0
xfeed_11465 0 1 decap_w0
xfeed_11464 0 1 decap_w0
xfeed_11463 0 1 decap_w0
xfeed_11462 0 1 decap_w0
xfeed_11461 0 1 decap_w0
xfeed_11460 0 1 decap_w0
xfeed_10939 0 1 decap_w0
xfeed_10938 0 1 decap_w0
xfeed_10937 0 1 decap_w0
xfeed_10936 0 1 decap_w0
xfeed_10935 0 1 decap_w0
xfeed_10934 0 1 decap_w0
xfeed_10933 0 1 decap_w0
xfeed_10932 0 1 decap_w0
xfeed_10931 0 1 decap_w0
xfeed_10930 0 1 decap_w0
xsubckt_870_mux2_x1 0 1 1612 1613 2002 445 mux2_x1
xsubckt_785_nand2_x0 0 1 1686 1996 1746 nand2_x0
xsubckt_164_nand3_x0 0 1 597 716 1924 599 nand3_x0
xsubckt_387_and2_x1 0 1 362 367 363 and2_x1
xsubckt_449_nexor2_x0 0 1 301 637 633 nexor2_x0
xsubckt_1565_and3_x1 0 1 1029 1037 1033 1031 and3_x1
xfeed_9579 0 1 decap_w0
xfeed_9578 0 1 decap_w0
xfeed_9577 0 1 decap_w0
xfeed_9576 0 1 decap_w0
xfeed_9575 0 1 decap_w0
xfeed_9574 0 1 decap_w0
xfeed_9573 0 1 decap_w0
xfeed_9572 0 1 decap_w0
xfeed_9571 0 1 decap_w0
xfeed_9570 0 1 tie
xfeed_5269 0 1 decap_w0
xfeed_5268 0 1 decap_w0
xfeed_5267 0 1 decap_w0
xfeed_5266 0 1 decap_w0
xfeed_5265 0 1 decap_w0
xfeed_5264 0 1 decap_w0
xfeed_5263 0 1 decap_w0
xfeed_5262 0 1 decap_w0
xfeed_5261 0 1 decap_w0
xfeed_5260 0 1 decap_w0
xfeed_4739 0 1 decap_w0
xfeed_4738 0 1 decap_w0
xfeed_4736 0 1 decap_w0
xfeed_4735 0 1 tie
xfeed_4734 0 1 decap_w0
xfeed_4733 0 1 decap_w0
xfeed_4732 0 1 decap_w0
xfeed_4731 0 1 tie
xsubckt_1042_and3_x1 0 1 1496 623 526 519 and3_x1
xsubckt_1021_nand2_x0 0 1 1512 623 1537 nand2_x0
xsubckt_694_or2_x1 0 1 2075 1776 1770 or2_x1
xsubckt_503_nand4_x0 0 1 248 1925 711 557 405 nand4_x0
xfeed_11479 0 1 decap_w0
xfeed_11478 0 1 decap_w0
xfeed_11477 0 1 decap_w0
xfeed_11476 0 1 decap_w0
xfeed_11475 0 1 decap_w0
xfeed_11474 0 1 decap_w0
xfeed_11473 0 1 decap_w0
xfeed_11472 0 1 tie
xfeed_11471 0 1 decap_w0
xfeed_11470 0 1 decap_w0
xfeed_10949 0 1 decap_w0
xfeed_10948 0 1 decap_w0
xfeed_10947 0 1 decap_w0
xfeed_10946 0 1 decap_w0
xfeed_10945 0 1 decap_w0
xfeed_10944 0 1 decap_w0
xfeed_10943 0 1 decap_w0
xfeed_10942 0 1 decap_w0
xfeed_10941 0 1 decap_w0
xfeed_10940 0 1 decap_w0
xfeed_9589 0 1 decap_w0
xfeed_9588 0 1 decap_w0
xfeed_9587 0 1 tie
xfeed_9586 0 1 decap_w0
xfeed_9585 0 1 decap_w0
xfeed_9584 0 1 decap_w0
xfeed_9583 0 1 decap_w0
xfeed_9581 0 1 decap_w0
xfeed_9580 0 1 decap_w0
xfeed_5279 0 1 decap_w0
xfeed_5278 0 1 decap_w0
xfeed_5277 0 1 tie
xfeed_5276 0 1 tie
xfeed_5275 0 1 decap_w0
xfeed_5274 0 1 decap_w0
xfeed_5273 0 1 decap_w0
xfeed_5272 0 1 decap_w0
xfeed_5271 0 1 decap_w0
xfeed_5270 0 1 decap_w0
xfeed_4749 0 1 decap_w0
xfeed_4748 0 1 decap_w0
xfeed_4747 0 1 decap_w0
xfeed_4746 0 1 decap_w0
xfeed_4745 0 1 tie
xfeed_4744 0 1 decap_w0
xfeed_4743 0 1 decap_w0
xfeed_4742 0 1 decap_w0
xfeed_4741 0 1 decap_w0
xfeed_4740 0 1 decap_w0
xsubckt_1112_mux2_x1 0 1 1845 2003 1994 1438 mux2_x1
xsubckt_652_and2_x1 0 1 107 111 110 and2_x1
xsubckt_177_and3_x1 0 1 581 714 1928 674 and3_x1
xsubckt_480_or21nand_x0 0 1 270 535 311 310 or21nand_x0
xsubckt_586_and4_x1 0 1 169 174 173 171 170 and4_x1
xsubckt_1421_and2_x1 0 1 1172 1178 1173 and2_x1
xsubckt_1548_nand2_x0 0 1 1046 1050 1048 nand2_x0
xsubckt_1550_or21nand_x0 0 1 1044 1105 1051 1049 or21nand_x0
xfeed_11489 0 1 decap_w0
xfeed_11488 0 1 decap_w0
xfeed_11487 0 1 decap_w0
xfeed_11486 0 1 decap_w0
xfeed_11485 0 1 decap_w0
xfeed_11484 0 1 decap_w0
xfeed_11483 0 1 decap_w0
xfeed_11482 0 1 decap_w0
xfeed_11481 0 1 tie
xfeed_11480 0 1 decap_w0
xfeed_10959 0 1 decap_w0
xfeed_10958 0 1 decap_w0
xfeed_10957 0 1 decap_w0
xfeed_10956 0 1 decap_w0
xfeed_10955 0 1 decap_w0
xfeed_10954 0 1 decap_w0
xfeed_10953 0 1 decap_w0
xfeed_10952 0 1 decap_w0
xfeed_10951 0 1 decap_w0
xfeed_10950 0 1 decap_w0
xsubckt_648_and2_x1 0 1 111 166 112 and2_x1
xsubckt_508_and4_x1 0 1 243 254 253 250 244 and4_x1
xsubckt_1747_or21nand_x0 0 1 847 861 859 856 or21nand_x0
xfeed_12100 0 1 decap_w0
xfeed_9599 0 1 decap_w0
xfeed_9598 0 1 decap_w0
xfeed_9597 0 1 decap_w0
xfeed_9596 0 1 decap_w0
xfeed_9595 0 1 decap_w0
xfeed_9594 0 1 decap_w0
xfeed_9593 0 1 decap_w0
xfeed_9592 0 1 decap_w0
xfeed_9591 0 1 decap_w0
xfeed_9590 0 1 decap_w0
xfeed_5289 0 1 tie
xfeed_5288 0 1 decap_w0
xfeed_5287 0 1 decap_w0
xfeed_5286 0 1 decap_w0
xfeed_5285 0 1 decap_w0
xfeed_5284 0 1 decap_w0
xfeed_5283 0 1 decap_w0
xfeed_5282 0 1 tie
xfeed_5281 0 1 decap_w0
xfeed_4759 0 1 decap_w0
xfeed_4758 0 1 decap_w0
xfeed_4757 0 1 decap_w0
xfeed_4756 0 1 decap_w0
xfeed_4755 0 1 decap_w0
xfeed_4754 0 1 decap_w0
xfeed_4753 0 1 decap_w0
xfeed_4751 0 1 decap_w0
xsubckt_1278_nand2_x0 0 1 1303 1308 1304 nand2_x0
xsubckt_1020_mux2_x1 0 1 1862 1548 1933 1576 mux2_x1
xsubckt_1650_or21nand_x0 0 1 944 946 947 1075 or21nand_x0
xsubckt_1708_and21nor_x0 0 1 886 1070 897 1073 and21nor_x0
xfeed_12109 0 1 decap_w0
xfeed_12108 0 1 decap_w0
xfeed_12107 0 1 decap_w0
xfeed_12106 0 1 decap_w0
xfeed_12105 0 1 decap_w0
xfeed_12104 0 1 decap_w0
xfeed_12103 0 1 decap_w0
xfeed_12102 0 1 decap_w0
xfeed_12101 0 1 decap_w0
xfeed_11499 0 1 decap_w0
xfeed_11498 0 1 decap_w0
xfeed_11497 0 1 tie
xfeed_11496 0 1 decap_w0
xfeed_11495 0 1 decap_w0
xfeed_11494 0 1 decap_w0
xfeed_11493 0 1 tie
xfeed_11492 0 1 decap_w0
xfeed_11491 0 1 decap_w0
xfeed_11490 0 1 decap_w0
xfeed_10969 0 1 decap_w0
xfeed_10968 0 1 decap_w0
xfeed_10967 0 1 decap_w0
xfeed_10966 0 1 decap_w0
xfeed_10965 0 1 decap_w0
xfeed_10964 0 1 decap_w0
xfeed_10963 0 1 decap_w0
xfeed_10962 0 1 decap_w0
xfeed_10961 0 1 decap_w0
xfeed_10960 0 1 decap_w0
xsubckt_494_nand3_x0 0 1 257 687 610 495 nand3_x0
xsubckt_1750_or21nand_x0 0 1 844 853 849 848 or21nand_x0
xfeed_5299 0 1 decap_w0
xfeed_5298 0 1 decap_w0
xfeed_5297 0 1 decap_w0
xfeed_5296 0 1 decap_w0
xfeed_5295 0 1 decap_w0
xfeed_5294 0 1 decap_w0
xfeed_5293 0 1 decap_w0
xfeed_5292 0 1 decap_w0
xfeed_5291 0 1 decap_w0
xfeed_5290 0 1 decap_w0
xfeed_4769 0 1 decap_w0
xfeed_4768 0 1 decap_w0
xfeed_4767 0 1 decap_w0
xfeed_4766 0 1 decap_w0
xfeed_4765 0 1 decap_w0
xfeed_4764 0 1 decap_w0
xfeed_4763 0 1 decap_w0
xfeed_4762 0 1 decap_w0
xfeed_4761 0 1 decap_w0
xfeed_4760 0 1 decap_w0
xsubckt_1098_nand2_x0 0 1 1449 631 1450 nand2_x0
xfeed_12119 0 1 decap_w0
xfeed_12118 0 1 decap_w0
xfeed_12117 0 1 decap_w0
xfeed_12116 0 1 decap_w0
xfeed_12115 0 1 decap_w0
xfeed_12114 0 1 decap_w0
xfeed_12113 0 1 decap_w0
xfeed_12112 0 1 decap_w0
xfeed_12111 0 1 decap_w0
xfeed_12110 0 1 decap_w0
xfeed_10979 0 1 decap_w0
xfeed_10978 0 1 decap_w0
xfeed_10977 0 1 decap_w0
xfeed_10976 0 1 decap_w0
xfeed_10975 0 1 decap_w0
xfeed_10974 0 1 decap_w0
xfeed_10973 0 1 decap_w0
xfeed_10972 0 1 decap_w0
xfeed_10971 0 1 decap_w0
xfeed_10970 0 1 decap_w0
xsubckt_909_and2_x1 0 1 1580 172 1620 and2_x1
xsubckt_1830_dff_x1 0 1 1927 26 74 dff_x1
xsubckt_1832_dff_x1 0 1 1925 24 74 dff_x1
xfeed_4779 0 1 decap_w0
xfeed_4778 0 1 tie
xfeed_4777 0 1 decap_w0
xfeed_4776 0 1 decap_w0
xfeed_4775 0 1 decap_w0
xfeed_4774 0 1 decap_w0
xfeed_4773 0 1 tie
xfeed_4772 0 1 decap_w0
xfeed_4771 0 1 decap_w0
xfeed_4770 0 1 decap_w0
xsubckt_1193_and3_x1 0 1 1371 1928 610 604 and3_x1
xsubckt_1834_dff_x1 0 1 2044 1904 35 dff_x1
xsubckt_1836_dff_x1 0 1 2042 1902 32 dff_x1
xfeed_12129 0 1 decap_w0
xfeed_12128 0 1 decap_w0
xfeed_12127 0 1 decap_w0
xfeed_12126 0 1 decap_w0
xfeed_12125 0 1 decap_w0
xfeed_12124 0 1 decap_w0
xfeed_12123 0 1 decap_w0
xfeed_12122 0 1 decap_w0
xfeed_12121 0 1 decap_w0
xfeed_12120 0 1 decap_w0
xfeed_10989 0 1 decap_w0
xfeed_10988 0 1 decap_w0
xfeed_10987 0 1 decap_w0
xfeed_10986 0 1 tie
xfeed_10985 0 1 decap_w0
xfeed_10984 0 1 decap_w0
xfeed_10983 0 1 decap_w0
xfeed_10982 0 1 decap_w0
xfeed_10981 0 1 decap_w0
xfeed_10980 0 1 decap_w0
xsubckt_817_and2_x1 0 1 1658 2050 1740 and2_x1
xsubckt_740_nand2_x0 0 1 2105 1732 1726 nand2_x0
xsubckt_1698_nand2_x0 0 1 896 899 898 nand2_x0
xsubckt_1838_dff_x1 0 1 2040 1900 32 dff_x1
xfeed_9709 0 1 decap_w0
xfeed_9708 0 1 decap_w0
xfeed_9707 0 1 decap_w0
xfeed_9706 0 1 tie
xfeed_9705 0 1 decap_w0
xfeed_9704 0 1 decap_w0
xfeed_9703 0 1 decap_w0
xfeed_9702 0 1 decap_w0
xfeed_9701 0 1 decap_w0
xfeed_9700 0 1 decap_w0
xfeed_4789 0 1 decap_w0
xfeed_4788 0 1 decap_w0
xfeed_4787 0 1 decap_w0
xfeed_4786 0 1 decap_w0
xfeed_4785 0 1 decap_w0
xfeed_4784 0 1 decap_w0
xfeed_4783 0 1 decap_w0
xfeed_4782 0 1 decap_w0
xfeed_4781 0 1 decap_w0
xfeed_4780 0 1 decap_w0
xsubckt_1189_and3_x1 0 1 1375 1378 1377 1376 and3_x1
xfeed_12139 0 1 decap_w0
xfeed_12138 0 1 decap_w0
xfeed_12137 0 1 decap_w0
xfeed_12136 0 1 decap_w0
xfeed_12135 0 1 decap_w0
xfeed_12134 0 1 decap_w0
xfeed_12133 0 1 decap_w0
xfeed_12132 0 1 decap_w0
xfeed_12131 0 1 decap_w0
xfeed_12130 0 1 decap_w0
xfeed_11609 0 1 decap_w0
xfeed_11608 0 1 decap_w0
xfeed_11607 0 1 decap_w0
xfeed_11606 0 1 tie
xfeed_11605 0 1 decap_w0
xfeed_11604 0 1 decap_w0
xfeed_11603 0 1 decap_w0
xfeed_11602 0 1 decap_w0
xfeed_11601 0 1 decap_w0
xfeed_11600 0 1 decap_w0
xfeed_10999 0 1 decap_w0
xfeed_10998 0 1 decap_w0
xfeed_10997 0 1 decap_w0
xfeed_10996 0 1 decap_w0
xfeed_10995 0 1 decap_w0
xfeed_10994 0 1 decap_w0
xfeed_10993 0 1 tie
xfeed_10992 0 1 decap_w0
xfeed_10991 0 1 decap_w0
xfeed_10990 0 1 decap_w0
xsubckt_939_mux2_x1 0 1 1879 1953 520 774 mux2_x1
xsubckt_1345_or21nand_x0 0 1 1807 1253 1246 1243 or21nand_x0
xsubckt_1432_and4_x1 0 1 1162 435 1635 1164 1163 and4_x1
xfeed_9719 0 1 decap_w0
xfeed_9718 0 1 decap_w0
xfeed_9717 0 1 decap_w0
xfeed_9716 0 1 decap_w0
xfeed_9715 0 1 decap_w0
xfeed_9714 0 1 decap_w0
xfeed_9713 0 1 decap_w0
xfeed_9712 0 1 decap_w0
xfeed_9711 0 1 decap_w0
xfeed_9710 0 1 decap_w0
xfeed_5409 0 1 decap_w0
xfeed_5408 0 1 decap_w0
xfeed_5407 0 1 decap_w0
xfeed_5405 0 1 decap_w0
xfeed_5404 0 1 decap_w0
xfeed_5403 0 1 decap_w0
xfeed_5402 0 1 decap_w0
xfeed_5401 0 1 decap_w0
xfeed_5400 0 1 decap_w0
xfeed_4799 0 1 decap_w0
xfeed_4798 0 1 decap_w0
xfeed_4797 0 1 decap_w0
xfeed_4796 0 1 decap_w0
xfeed_4795 0 1 decap_w0
xfeed_4794 0 1 decap_w0
xfeed_4793 0 1 decap_w0
xfeed_4792 0 1 decap_w0
xfeed_4791 0 1 decap_w0
xfeed_4790 0 1 decap_w0
xsubckt_1198_and21nor_x0 0 1 1366 459 606 614 and21nor_x0
xsubckt_1060_nand3_x0 0 1 1482 643 532 1483 nand3_x0
xsubckt_290_nand2_x0 0 1 458 616 460 nand2_x0
xsubckt_112_nand2_x0 0 1 656 1986 1990 nand2_x0
xsubckt_1503_nand2_x0 0 1 1093 1099 1095 nand2_x0
xsubckt_1762_nexor2_x0 0 1 832 935 835 nexor2_x0
xfeed_12149 0 1 decap_w0
xfeed_12148 0 1 decap_w0
xfeed_12147 0 1 decap_w0
xfeed_12146 0 1 decap_w0
xfeed_12145 0 1 decap_w0
xfeed_12144 0 1 decap_w0
xfeed_12143 0 1 decap_w0
xfeed_12142 0 1 decap_w0
xfeed_12141 0 1 decap_w0
xfeed_12140 0 1 decap_w0
xfeed_11619 0 1 decap_w0
xfeed_11618 0 1 decap_w0
xfeed_11617 0 1 decap_w0
xfeed_11616 0 1 decap_w0
xfeed_11615 0 1 decap_w0
xfeed_11614 0 1 decap_w0
xfeed_11613 0 1 tie
xfeed_11612 0 1 decap_w0
xfeed_11611 0 1 decap_w0
xfeed_11610 0 1 decap_w0
xfeed_1106 0 1 decap_w0
xfeed_1105 0 1 decap_w0
xfeed_1104 0 1 decap_w0
xfeed_1103 0 1 decap_w0
xfeed_1102 0 1 decap_w0
xfeed_1101 0 1 decap_w0
xfeed_1100 0 1 decap_w0
xsubckt_236_and21nor_x0 0 1 515 536 535 517 and21nor_x0
xsubckt_73_inv_x0 0 1 709 1932 inv_x0
xsubckt_71_inv_x0 0 1 711 1926 inv_x0
xsubckt_448_nor2_x0 0 1 302 382 303 nor2_x0
xsubckt_1323_nand2_x0 0 1 1809 1271 1263 nand2_x0
xsubckt_1445_or21nand_x0 0 1 1150 1151 1323 689 or21nand_x0
xsubckt_1616_mux2_x1 0 1 978 984 981 992 mux2_x1
xsubckt_1699_and21nor_x0 0 1 895 1104 899 898 and21nor_x0
xsubckt_1753_nexor2_x0 0 1 841 887 881 nexor2_x0
xfeed_9729 0 1 decap_w0
xfeed_9728 0 1 tie
xfeed_9727 0 1 decap_w0
xfeed_9726 0 1 decap_w0
xfeed_9725 0 1 decap_w0
xfeed_9724 0 1 decap_w0
xfeed_9723 0 1 decap_w0
xfeed_9722 0 1 decap_w0
xfeed_9721 0 1 decap_w0
xfeed_9720 0 1 decap_w0
xfeed_5419 0 1 decap_w0
xfeed_5417 0 1 decap_w0
xfeed_5416 0 1 decap_w0
xfeed_5415 0 1 decap_w0
xfeed_5414 0 1 decap_w0
xfeed_5411 0 1 decap_w0
xfeed_5410 0 1 tie
xfeed_1109 0 1 decap_w0
xfeed_1108 0 1 decap_w0
xfeed_1107 0 1 tie
xsubckt_1167_mux2_x1 0 1 1833 1965 1395 1403 mux2_x1
xsubckt_79_inv_x0 0 1 703 2089 inv_x0
xsubckt_77_inv_x0 0 1 705 2090 inv_x0
xsubckt_75_inv_x0 0 1 707 1950 inv_x0
xsubckt_158_and3_x1 0 1 603 1929 715 670 and3_x1
xsubckt_1497_nand3_x0 0 1 1099 1969 682 595 nand3_x0
xfeed_12159 0 1 decap_w0
xfeed_12158 0 1 decap_w0
xfeed_12157 0 1 decap_w0
xfeed_12156 0 1 decap_w0
xfeed_12155 0 1 decap_w0
xfeed_12154 0 1 decap_w0
xfeed_12153 0 1 tie
xfeed_12152 0 1 decap_w0
xfeed_12151 0 1 decap_w0
xfeed_12150 0 1 decap_w0
xfeed_11629 0 1 decap_w0
xfeed_11628 0 1 decap_w0
xfeed_11627 0 1 decap_w0
xfeed_11626 0 1 decap_w0
xfeed_11625 0 1 decap_w0
xfeed_11624 0 1 decap_w0
xfeed_11623 0 1 decap_w0
xfeed_11622 0 1 decap_w0
xfeed_11621 0 1 decap_w0
xfeed_11620 0 1 decap_w0
xfeed_1113 0 1 decap_w0
xfeed_1112 0 1 decap_w0
xfeed_1111 0 1 decap_w0
xfeed_1110 0 1 decap_w0
xsubckt_1143_nand2_x0 0 1 1836 1419 1416 nand2_x0
xsubckt_1310_and2_x1 0 1 1274 1283 1276 and2_x1
xfeed_9739 0 1 decap_w0
xfeed_9738 0 1 decap_w0
xfeed_9737 0 1 decap_w0
xfeed_9736 0 1 decap_w0
xfeed_9735 0 1 decap_w0
xfeed_9734 0 1 decap_w0
xfeed_9733 0 1 decap_w0
xfeed_9732 0 1 decap_w0
xfeed_9731 0 1 decap_w0
xfeed_9730 0 1 decap_w0
xfeed_5429 0 1 decap_w0
xfeed_5428 0 1 decap_w0
xfeed_5427 0 1 decap_w0
xfeed_5426 0 1 decap_w0
xfeed_5425 0 1 tie
xfeed_5424 0 1 decap_w0
xfeed_5423 0 1 decap_w0
xfeed_5422 0 1 decap_w0
xfeed_5421 0 1 decap_w0
xfeed_5420 0 1 tie
xfeed_1119 0 1 decap_w0
xfeed_1118 0 1 decap_w0
xfeed_1117 0 1 decap_w0
xfeed_1116 0 1 decap_w0
xfeed_1115 0 1 decap_w0
xfeed_1114 0 1 decap_w0
xcmpt_abc_11867_new_n543_hfns_0 0 1 533 531 buf_x4
xcmpt_abc_11867_new_n543_hfns_1 0 1 532 531 buf_x4
xcmpt_abc_11867_new_n543_hfns_2 0 1 531 534 buf_x4
xfeed_12169 0 1 decap_w0
xfeed_12168 0 1 decap_w0
xfeed_12167 0 1 decap_w0
xfeed_12166 0 1 decap_w0
xfeed_12165 0 1 decap_w0
xfeed_12164 0 1 decap_w0
xfeed_12163 0 1 decap_w0
xfeed_12162 0 1 decap_w0
xfeed_12161 0 1 decap_w0
xfeed_12160 0 1 decap_w0
xfeed_11639 0 1 decap_w0
xfeed_11638 0 1 decap_w0
xfeed_11637 0 1 decap_w0
xfeed_11636 0 1 tie
xfeed_11635 0 1 decap_w0
xfeed_11634 0 1 decap_w0
xfeed_11633 0 1 decap_w0
xfeed_11632 0 1 decap_w0
xfeed_11631 0 1 decap_w0
xfeed_11630 0 1 decap_w0
xfeed_1120 0 1 decap_w0
xsubckt_1306_and2_x1 0 1 1278 435 1279 and2_x1
xfeed_9749 0 1 decap_w0
xfeed_9748 0 1 decap_w0
xfeed_9747 0 1 decap_w0
xfeed_9746 0 1 decap_w0
xfeed_9745 0 1 tie
xfeed_9744 0 1 decap_w0
xfeed_9743 0 1 decap_w0
xfeed_9742 0 1 decap_w0
xfeed_9741 0 1 decap_w0
xfeed_9740 0 1 decap_w0
xfeed_5439 0 1 decap_w0
xfeed_5438 0 1 decap_w0
xfeed_5437 0 1 decap_w0
xfeed_5436 0 1 decap_w0
xfeed_5435 0 1 decap_w0
xfeed_5434 0 1 decap_w0
xfeed_5433 0 1 decap_w0
xfeed_5432 0 1 decap_w0
xfeed_5430 0 1 tie
xfeed_4909 0 1 decap_w0
xfeed_4908 0 1 decap_w0
xfeed_4907 0 1 decap_w0
xfeed_4906 0 1 decap_w0
xfeed_4905 0 1 decap_w0
xfeed_4904 0 1 decap_w0
xfeed_4903 0 1 tie
xfeed_4902 0 1 decap_w0
xfeed_4901 0 1 decap_w0
xfeed_4900 0 1 decap_w0
xfeed_1129 0 1 decap_w0
xfeed_1128 0 1 decap_w0
xfeed_1127 0 1 decap_w0
xfeed_1126 0 1 decap_w0
xfeed_1125 0 1 decap_w0
xfeed_1124 0 1 tie
xfeed_1123 0 1 decap_w0
xfeed_1122 0 1 decap_w0
xfeed_1121 0 1 decap_w0
xsubckt_1266_and3_x1 0 1 1314 2065 666 657 and3_x1
xsubckt_1786_nexor2_x0 0 1 808 1036 1030 nexor2_x0
xsubckt_1795_nexor2_x0 0 1 799 816 813 nexor2_x0
xfeed_12179 0 1 decap_w0
xfeed_12178 0 1 decap_w0
xfeed_12177 0 1 decap_w0
xfeed_12176 0 1 decap_w0
xfeed_12175 0 1 decap_w0
xfeed_12174 0 1 decap_w0
xfeed_12173 0 1 decap_w0
xfeed_12172 0 1 decap_w0
xfeed_12171 0 1 decap_w0
xfeed_12170 0 1 decap_w0
xfeed_11649 0 1 decap_w0
xfeed_11648 0 1 decap_w0
xfeed_11647 0 1 decap_w0
xfeed_11646 0 1 decap_w0
xfeed_11645 0 1 decap_w0
xfeed_11644 0 1 decap_w0
xfeed_11643 0 1 decap_w0
xfeed_11642 0 1 decap_w0
xfeed_11641 0 1 decap_w0
xfeed_11640 0 1 decap_w0
xsubckt_1214_and2_x1 0 1 1350 592 587 and2_x1
xsubckt_840_and21nor_x0 0 1 1638 690 1755 1754 and21nor_x0
xsubckt_172_nor2_x0 0 1 586 2055 1921 nor2_x0
xsubckt_1623_and3_x1 0 1 971 977 974 973 and3_x1
xsubckt_1739_nand3_x0 0 1 855 1069 873 871 nand3_x0
xfeed_9759 0 1 decap_w0
xfeed_9758 0 1 decap_w0
xfeed_9757 0 1 decap_w0
xfeed_9756 0 1 decap_w0
xfeed_9755 0 1 decap_w0
xfeed_9754 0 1 decap_w0
xfeed_9753 0 1 decap_w0
xfeed_9752 0 1 tie
xfeed_9751 0 1 decap_w0
xfeed_9750 0 1 decap_w0
xfeed_5449 0 1 decap_w0
xfeed_5448 0 1 decap_w0
xfeed_5447 0 1 decap_w0
xfeed_5446 0 1 tie
xfeed_5445 0 1 decap_w0
xfeed_5444 0 1 decap_w0
xfeed_5443 0 1 decap_w0
xfeed_5442 0 1 decap_w0
xfeed_5441 0 1 decap_w0
xfeed_5440 0 1 decap_w0
xfeed_4919 0 1 decap_w0
xfeed_4918 0 1 decap_w0
xfeed_4917 0 1 decap_w0
xfeed_4916 0 1 decap_w0
xfeed_4915 0 1 tie
xfeed_4914 0 1 decap_w0
xfeed_4913 0 1 decap_w0
xfeed_4912 0 1 decap_w0
xfeed_4911 0 1 decap_w0
xfeed_4910 0 1 decap_w0
xfeed_1139 0 1 decap_w0
xfeed_1138 0 1 decap_w0
xfeed_1137 0 1 decap_w0
xfeed_1136 0 1 tie
xfeed_1135 0 1 decap_w0
xfeed_1134 0 1 decap_w0
xfeed_1133 0 1 decap_w0
xfeed_1132 0 1 decap_w0
xfeed_1131 0 1 decap_w0
xfeed_1130 0 1 decap_w0
xsubckt_969_nand2_x0 0 1 1556 1956 1575 nand2_x0
xsubckt_924_mux2_x1 0 1 1892 1593 2032 1579 mux2_x1
xsubckt_353_and2_x1 0 1 395 680 405 and2_x1
xsubckt_1768_nexor2_x0 0 1 826 839 836 nexor2_x0
xfeed_12189 0 1 decap_w0
xfeed_12188 0 1 decap_w0
xfeed_12187 0 1 decap_w0
xfeed_12186 0 1 decap_w0
xfeed_12185 0 1 decap_w0
xfeed_12184 0 1 decap_w0
xfeed_12183 0 1 decap_w0
xfeed_12182 0 1 decap_w0
xfeed_12181 0 1 decap_w0
xfeed_12180 0 1 decap_w0
xfeed_11659 0 1 tie
xfeed_11658 0 1 decap_w0
xfeed_11657 0 1 decap_w0
xfeed_11656 0 1 decap_w0
xfeed_11655 0 1 decap_w0
xfeed_11654 0 1 decap_w0
xfeed_11653 0 1 decap_w0
xfeed_11652 0 1 decap_w0
xfeed_11651 0 1 decap_w0
xfeed_11650 0 1 decap_w0
xsubckt_401_mux2_x1 0 1 348 1965 1966 1952 mux2_x1
xfeed_9769 0 1 decap_w0
xfeed_9768 0 1 decap_w0
xfeed_9767 0 1 decap_w0
xfeed_9766 0 1 tie
xfeed_9765 0 1 decap_w0
xfeed_9764 0 1 decap_w0
xfeed_9763 0 1 decap_w0
xfeed_9762 0 1 decap_w0
xfeed_9761 0 1 decap_w0
xfeed_9760 0 1 decap_w0
xfeed_5459 0 1 decap_w0
xfeed_5458 0 1 decap_w0
xfeed_5457 0 1 decap_w0
xfeed_5456 0 1 decap_w0
xfeed_5455 0 1 decap_w0
xfeed_5454 0 1 tie
xfeed_5453 0 1 decap_w0
xfeed_5452 0 1 decap_w0
xfeed_5451 0 1 decap_w0
xfeed_5450 0 1 decap_w0
xfeed_4929 0 1 decap_w0
xfeed_4928 0 1 decap_w0
xfeed_4927 0 1 tie
xfeed_4926 0 1 decap_w0
xfeed_4925 0 1 decap_w0
xfeed_4924 0 1 decap_w0
xfeed_4923 0 1 decap_w0
xfeed_4922 0 1 tie
xfeed_4921 0 1 decap_w0
xfeed_4920 0 1 decap_w0
xfeed_1149 0 1 decap_w0
xfeed_1148 0 1 decap_w0
xfeed_1147 0 1 tie
xfeed_1146 0 1 decap_w0
xfeed_1145 0 1 decap_w0
xfeed_1144 0 1 decap_w0
xfeed_1143 0 1 decap_w0
xfeed_1142 0 1 decap_w0
xfeed_1141 0 1 decap_w0
xfeed_1140 0 1 tie
xsubckt_1244_mux2_x1 0 1 1817 2101 2068 1334 mux2_x1
xsubckt_952_nand2_x0 0 1 1568 1937 1575 nand2_x0
xsubckt_775_or21nand_x0 0 1 1695 2059 1742 1740 or21nand_x0
xsubckt_758_and3_x1 0 1 1710 1972 1749 1739 and3_x1
xsubckt_699_nand2_x0 0 1 1765 168 1766 nand2_x0
xsubckt_1293_nand2_x0 0 1 1290 775 1973 nand2_x0
xfeed_12199 0 1 decap_w0
xfeed_12198 0 1 decap_w0
xfeed_12197 0 1 decap_w0
xfeed_12196 0 1 tie
xfeed_12195 0 1 decap_w0
xfeed_12194 0 1 decap_w0
xfeed_12193 0 1 decap_w0
xfeed_12192 0 1 decap_w0
xfeed_12191 0 1 decap_w0
xfeed_12190 0 1 decap_w0
xfeed_11669 0 1 decap_w0
xfeed_11668 0 1 decap_w0
xfeed_11667 0 1 decap_w0
xfeed_11666 0 1 decap_w0
xfeed_11665 0 1 decap_w0
xfeed_11664 0 1 decap_w0
xfeed_11663 0 1 decap_w0
xfeed_11662 0 1 decap_w0
xfeed_11661 0 1 decap_w0
xfeed_11660 0 1 decap_w0
xsubckt_1798_and21nor_x0 0 1 796 830 799 797 and21nor_x0
xfeed_9779 0 1 decap_w0
xfeed_9778 0 1 decap_w0
xfeed_9777 0 1 decap_w0
xfeed_9775 0 1 decap_w0
xfeed_9774 0 1 decap_w0
xfeed_9773 0 1 decap_w0
xfeed_9772 0 1 decap_w0
xfeed_9771 0 1 decap_w0
xfeed_9770 0 1 decap_w0
xfeed_5469 0 1 tie
xfeed_5468 0 1 decap_w0
xfeed_5467 0 1 decap_w0
xfeed_5466 0 1 decap_w0
xfeed_5465 0 1 decap_w0
xfeed_5464 0 1 tie
xfeed_5463 0 1 decap_w0
xfeed_5462 0 1 decap_w0
xfeed_5461 0 1 decap_w0
xfeed_5460 0 1 decap_w0
xfeed_4939 0 1 decap_w0
xfeed_4938 0 1 decap_w0
xfeed_4936 0 1 decap_w0
xfeed_4935 0 1 decap_w0
xfeed_4934 0 1 tie
xfeed_4933 0 1 decap_w0
xfeed_4932 0 1 decap_w0
xfeed_4931 0 1 decap_w0
xfeed_4930 0 1 decap_w0
xfeed_1159 0 1 decap_w0
xfeed_1158 0 1 decap_w0
xfeed_1157 0 1 decap_w0
xfeed_1156 0 1 tie
xfeed_1155 0 1 decap_w0
xfeed_1154 0 1 decap_w0
xfeed_1153 0 1 decap_w0
xfeed_1152 0 1 decap_w0
xfeed_1151 0 1 decap_w0
xfeed_1150 0 1 decap_w0
xsubckt_1397_and21nor_x0 0 1 1194 774 1206 1197 and21nor_x0
xfeed_11679 0 1 decap_w0
xfeed_11678 0 1 decap_w0
xfeed_11677 0 1 decap_w0
xfeed_11676 0 1 decap_w0
xfeed_11675 0 1 decap_w0
xfeed_11674 0 1 decap_w0
xfeed_11673 0 1 decap_w0
xfeed_11672 0 1 decap_w0
xfeed_11671 0 1 decap_w0
xfeed_11670 0 1 decap_w0
xsubckt_1148_mux2_x1 0 1 1411 1412 2000 484 mux2_x1
xsubckt_836_and21nor_x0 0 1 1641 742 600 1745 and21nor_x0
xsubckt_682_nand2_x0 0 1 1781 1784 1783 nand2_x0
xsubckt_504_nand2_x0 0 1 247 686 506 nand2_x0
xsubckt_574_and3_x1 0 1 181 195 194 182 and3_x1
xfeed_9789 0 1 decap_w0
xfeed_9788 0 1 decap_w0
xfeed_9787 0 1 decap_w0
xfeed_9786 0 1 decap_w0
xfeed_9785 0 1 decap_w0
xfeed_9784 0 1 decap_w0
xfeed_9783 0 1 tie
xfeed_9782 0 1 decap_w0
xfeed_9781 0 1 decap_w0
xfeed_9780 0 1 decap_w0
xfeed_5479 0 1 decap_w0
xfeed_5478 0 1 tie
xfeed_5477 0 1 decap_w0
xfeed_5476 0 1 decap_w0
xfeed_5475 0 1 decap_w0
xfeed_5474 0 1 decap_w0
xfeed_5473 0 1 decap_w0
xfeed_5472 0 1 decap_w0
xfeed_5471 0 1 decap_w0
xfeed_5470 0 1 decap_w0
xfeed_4949 0 1 decap_w0
xfeed_4948 0 1 decap_w0
xfeed_4947 0 1 decap_w0
xfeed_4946 0 1 decap_w0
xfeed_4945 0 1 decap_w0
xfeed_4944 0 1 decap_w0
xfeed_4943 0 1 decap_w0
xfeed_4942 0 1 decap_w0
xfeed_4941 0 1 decap_w0
xfeed_4940 0 1 decap_w0
xfeed_1169 0 1 decap_w0
xfeed_1168 0 1 decap_w0
xfeed_1167 0 1 decap_w0
xfeed_1166 0 1 tie
xfeed_1165 0 1 decap_w0
xfeed_1164 0 1 decap_w0
xfeed_1163 0 1 decap_w0
xfeed_1162 0 1 decap_w0
xfeed_1161 0 1 decap_w0
xfeed_1160 0 1 decap_w0
xsubckt_1004_nand3_x0 0 1 1525 627 532 1563 nand3_x0
xsubckt_310_nand4_x0 0 1 438 1927 713 681 589 nand4_x0
xfeed_11689 0 1 decap_w0
xfeed_11688 0 1 decap_w0
xfeed_11687 0 1 decap_w0
xfeed_11686 0 1 decap_w0
xfeed_11685 0 1 decap_w0
xfeed_11684 0 1 decap_w0
xfeed_11683 0 1 decap_w0
xfeed_11682 0 1 decap_w0
xfeed_11681 0 1 decap_w0
xfeed_11680 0 1 decap_w0
xsubckt_1056_mux2_x1 0 1 1853 1486 1948 1576 mux2_x1
xsubckt_979_and4_x1 0 1 1548 637 633 622 520 and4_x1
xsubckt_596_and2_x1 0 1 159 162 161 and2_x1
xsubckt_1491_mux2_x1 0 1 1105 1107 739 1143 mux2_x1
xsubckt_1541_nor2_x0 0 1 1053 1059 1054 nor2_x0
xfeed_9799 0 1 decap_w0
xfeed_9798 0 1 decap_w0
xfeed_9797 0 1 decap_w0
xfeed_9796 0 1 decap_w0
xfeed_9795 0 1 decap_w0
xfeed_9794 0 1 decap_w0
xfeed_9793 0 1 decap_w0
xfeed_9792 0 1 decap_w0
xfeed_9791 0 1 decap_w0
xfeed_9790 0 1 decap_w0
xfeed_5489 0 1 decap_w0
xfeed_5488 0 1 decap_w0
xfeed_5487 0 1 decap_w0
xfeed_5486 0 1 decap_w0
xfeed_5485 0 1 decap_w0
xfeed_5484 0 1 decap_w0
xfeed_5483 0 1 decap_w0
xfeed_5482 0 1 decap_w0
xfeed_5481 0 1 decap_w0
xfeed_5480 0 1 decap_w0
xfeed_4959 0 1 decap_w0
xfeed_4958 0 1 decap_w0
xfeed_4957 0 1 decap_w0
xfeed_4956 0 1 decap_w0
xfeed_4955 0 1 decap_w0
xfeed_4954 0 1 decap_w0
xfeed_4953 0 1 tie
xfeed_4952 0 1 decap_w0
xfeed_4951 0 1 decap_w0
xfeed_4950 0 1 decap_w0
xfeed_1179 0 1 decap_w0
xfeed_1178 0 1 decap_w0
xfeed_1177 0 1 decap_w0
xfeed_1175 0 1 decap_w0
xfeed_1174 0 1 decap_w0
xfeed_1173 0 1 tie
xfeed_1172 0 1 decap_w0
xfeed_1171 0 1 decap_w0
xfeed_1170 0 1 decap_w0
xsubckt_430_and2_x1 0 1 319 332 320 and2_x1
xsubckt_518_and2_x1 0 1 233 271 234 and2_x1
xsubckt_1355_nand2_x0 0 1 1233 1245 1234 nand2_x0
xsubckt_1365_and2_x1 0 1 1224 1228 1225 and2_x1
xfeed_12309 0 1 tie
xfeed_12308 0 1 decap_w0
xfeed_12307 0 1 decap_w0
xfeed_12306 0 1 decap_w0
xfeed_12305 0 1 decap_w0
xfeed_12304 0 1 decap_w0
xfeed_12303 0 1 decap_w0
xfeed_12302 0 1 decap_w0
xfeed_12301 0 1 decap_w0
xfeed_12300 0 1 tie
xfeed_11699 0 1 decap_w0
xfeed_11698 0 1 decap_w0
xfeed_11697 0 1 decap_w0
xfeed_11696 0 1 decap_w0
xfeed_11695 0 1 decap_w0
xfeed_11694 0 1 decap_w0
xfeed_11693 0 1 decap_w0
xfeed_11692 0 1 decap_w0
xfeed_11691 0 1 decap_w0
xfeed_11690 0 1 decap_w0
xsubckt_1251_nand4_x0 0 1 1329 716 1924 711 670 nand4_x0
xsubckt_1139_or21nand_x0 0 1 1419 1995 1424 1422 or21nand_x0
xsubckt_117_mux2_x1 0 1 651 1991 2000 1986 mux2_x1
xsubckt_1299_and4_x1 0 1 1284 1311 1303 1293 1285 and4_x1
xsubckt_1304_and21nor_x0 0 1 1280 751 478 1317 and21nor_x0
xsubckt_1659_nexor2_x0 0 1 935 948 941 nexor2_x0
xfeed_6109 0 1 decap_w0
xfeed_6108 0 1 decap_w0
xfeed_6107 0 1 decap_w0
xfeed_6106 0 1 decap_w0
xfeed_6105 0 1 decap_w0
xfeed_6104 0 1 decap_w0
xfeed_6103 0 1 decap_w0
xfeed_6102 0 1 decap_w0
xfeed_6101 0 1 decap_w0
xfeed_6100 0 1 tie
xfeed_5499 0 1 decap_w0
xfeed_5498 0 1 decap_w0
xfeed_5497 0 1 decap_w0
xfeed_5496 0 1 decap_w0
xfeed_5495 0 1 decap_w0
xfeed_5494 0 1 decap_w0
xfeed_5492 0 1 decap_w0
xfeed_5491 0 1 decap_w0
xfeed_5490 0 1 decap_w0
xfeed_4969 0 1 decap_w0
xfeed_4968 0 1 decap_w0
xfeed_4967 0 1 decap_w0
xfeed_4966 0 1 decap_w0
xfeed_4965 0 1 decap_w0
xfeed_4964 0 1 decap_w0
xfeed_4963 0 1 decap_w0
xfeed_4962 0 1 decap_w0
xfeed_4961 0 1 tie
xfeed_4960 0 1 decap_w0
xfeed_1189 0 1 decap_w0
xfeed_1188 0 1 tie
xfeed_1187 0 1 decap_w0
xfeed_1186 0 1 decap_w0
xfeed_1185 0 1 decap_w0
xfeed_1184 0 1 decap_w0
xfeed_1183 0 1 decap_w0
xfeed_1182 0 1 decap_w0
xfeed_1181 0 1 decap_w0
xfeed_1180 0 1 decap_w0
xsubckt_1085_nand2_x0 0 1 1460 313 1496 nand2_x0
xsubckt_853_or4_x1 0 1 1626 1631 1630 1629 1627 or4_x1
xsubckt_676_nor2_x0 0 1 85 87 86 nor2_x0
xsubckt_200_or2_x1 0 1 554 1917 18 or2_x1
xsubckt_426_and2_x1 0 1 323 326 324 and2_x1
xsubckt_481_nand3_x0 0 1 269 610 581 558 nand3_x0
xsubckt_1604_and3_x1 0 1 990 1972 680 594 and3_x1
xsubckt_1841_dff_x1 0 1 2037 1897 35 dff_x1
xsubckt_1843_dff_x1 0 1 2035 1895 35 dff_x1
xfeed_12319 0 1 decap_w0
xfeed_12318 0 1 decap_w0
xfeed_12317 0 1 decap_w0
xfeed_12316 0 1 decap_w0
xfeed_12315 0 1 decap_w0
xfeed_12314 0 1 decap_w0
xfeed_12313 0 1 decap_w0
xfeed_12312 0 1 decap_w0
xfeed_12311 0 1 decap_w0
xfeed_12310 0 1 decap_w0
xsubckt_386_and3_x1 0 1 363 366 365 364 and3_x1
xsubckt_1845_dff_x1 0 1 2033 1893 35 dff_x1
xsubckt_1847_dff_x1 0 1 2031 1891 32 dff_x1
xsubckt_1849_dff_x1 0 1 2029 1889 32 dff_x1
xfeed_6119 0 1 decap_w0
xfeed_6118 0 1 decap_w0
xfeed_6117 0 1 tie
xfeed_6116 0 1 decap_w0
xfeed_6115 0 1 decap_w0
xfeed_6114 0 1 decap_w0
xfeed_6113 0 1 decap_w0
xfeed_6112 0 1 decap_w0
xfeed_6111 0 1 decap_w0
xfeed_6110 0 1 decap_w0
xfeed_4979 0 1 decap_w0
xfeed_4978 0 1 decap_w0
xfeed_4977 0 1 decap_w0
xfeed_4976 0 1 decap_w0
xfeed_4975 0 1 decap_w0
xfeed_4974 0 1 decap_w0
xfeed_4973 0 1 tie
xfeed_4972 0 1 decap_w0
xfeed_4971 0 1 decap_w0
xfeed_4970 0 1 decap_w0
xfeed_1199 0 1 decap_w0
xfeed_1198 0 1 decap_w0
xfeed_1197 0 1 tie
xfeed_1196 0 1 decap_w0
xfeed_1195 0 1 decap_w0
xfeed_1194 0 1 decap_w0
xfeed_1193 0 1 decap_w0
xfeed_1192 0 1 decap_w0
xfeed_1191 0 1 decap_w0
xfeed_1190 0 1 decap_w0
xsubckt_1626_and2_x1 0 1 968 1656 969 and2_x1
xfeed_12329 0 1 tie
xfeed_12328 0 1 decap_w0
xfeed_12327 0 1 decap_w0
xfeed_12326 0 1 decap_w0
xfeed_12325 0 1 decap_w0
xfeed_12324 0 1 decap_w0
xfeed_12323 0 1 decap_w0
xfeed_12322 0 1 decap_w0
xfeed_12321 0 1 decap_w0
xfeed_12320 0 1 decap_w0
xsubckt_1154_nand3_x0 0 1 1406 484 1437 1408 nand3_x0
xsubckt_1103_and21nor_x0 0 1 1444 1575 1451 1445 and21nor_x0
xsubckt_474_nand2_x0 0 1 276 558 552 nand2_x0
xsubckt_1504_and21nor_x0 0 1 1092 1104 1099 1095 and21nor_x0
xfeed_9909 0 1 decap_w0
xfeed_9908 0 1 decap_w0
xfeed_9907 0 1 decap_w0
xfeed_9906 0 1 decap_w0
xfeed_9905 0 1 decap_w0
xfeed_9904 0 1 decap_w0
xfeed_9903 0 1 decap_w0
xfeed_9902 0 1 decap_w0
xfeed_9901 0 1 decap_w0
xfeed_9900 0 1 decap_w0
xfeed_6129 0 1 decap_w0
xfeed_6128 0 1 decap_w0
xfeed_6127 0 1 decap_w0
xfeed_6125 0 1 decap_w0
xfeed_6124 0 1 decap_w0
xfeed_6123 0 1 decap_w0
xfeed_6122 0 1 decap_w0
xfeed_6121 0 1 decap_w0
xfeed_6120 0 1 decap_w0
xfeed_4989 0 1 decap_w0
xfeed_4988 0 1 decap_w0
xfeed_4987 0 1 decap_w0
xfeed_4986 0 1 decap_w0
xfeed_4985 0 1 tie
xfeed_4984 0 1 decap_w0
xfeed_4983 0 1 decap_w0
xfeed_4982 0 1 decap_w0
xfeed_4981 0 1 decap_w0
xfeed_4980 0 1 decap_w0
xsubckt_1064_nand3_x0 0 1 1478 1484 1481 1479 nand3_x0
xsubckt_1447_or2_x1 0 1 1148 1154 1150 or2_x1
xsubckt_1507_nand2_x0 0 1 1089 1091 1090 nand2_x0
xfeed_12339 0 1 decap_w0
xfeed_12338 0 1 decap_w0
xfeed_12337 0 1 decap_w0
xfeed_12336 0 1 decap_w0
xfeed_12335 0 1 decap_w0
xfeed_12334 0 1 decap_w0
xfeed_12333 0 1 decap_w0
xfeed_12332 0 1 decap_w0
xfeed_12331 0 1 decap_w0
xfeed_12330 0 1 decap_w0
xfeed_11809 0 1 decap_w0
xfeed_11808 0 1 decap_w0
xfeed_11807 0 1 decap_w0
xfeed_11806 0 1 decap_w0
xfeed_11805 0 1 decap_w0
xfeed_11804 0 1 decap_w0
xfeed_11803 0 1 decap_w0
xfeed_11802 0 1 decap_w0
xfeed_11801 0 1 decap_w0
xfeed_11800 0 1 decap_w0
xsubckt_1133_mux2_x1 0 1 1837 1425 1966 1431 mux2_x1
xsubckt_987_nand4_x0 0 1 1540 1550 1549 1547 1542 nand4_x0
xsubckt_887_mux2_x1 0 1 1909 2017 1599 1619 mux2_x1
xsubckt_80_inv_x0 0 1 702 2009 inv_x0
xsubckt_116_nand2_x0 0 1 652 659 654 nand2_x0
xsubckt_150_and2_x1 0 1 618 712 1926 and2_x1
xsubckt_533_and4_x1 0 1 220 442 441 415 413 and4_x1
xsubckt_1417_nand2_x0 0 1 1176 2048 479 nand2_x0
xfeed_9919 0 1 tie
xfeed_9918 0 1 decap_w0
xfeed_9917 0 1 decap_w0
xfeed_9916 0 1 decap_w0
xfeed_9915 0 1 decap_w0
xfeed_9914 0 1 decap_w0
xfeed_9913 0 1 decap_w0
xfeed_9912 0 1 decap_w0
xfeed_9911 0 1 decap_w0
xfeed_9910 0 1 decap_w0
xfeed_6139 0 1 decap_w0
xfeed_6138 0 1 decap_w0
xfeed_6137 0 1 decap_w0
xfeed_6136 0 1 decap_w0
xfeed_6135 0 1 decap_w0
xfeed_6134 0 1 decap_w0
xfeed_6133 0 1 decap_w0
xfeed_6132 0 1 decap_w0
xfeed_6131 0 1 decap_w0
xfeed_6130 0 1 decap_w0
xfeed_5609 0 1 decap_w0
xfeed_5608 0 1 decap_w0
xfeed_5606 0 1 decap_w0
xfeed_5605 0 1 decap_w0
xfeed_5603 0 1 decap_w0
xfeed_5602 0 1 decap_w0
xfeed_5601 0 1 decap_w0
xfeed_5600 0 1 decap_w0
xfeed_4999 0 1 decap_w0
xfeed_4998 0 1 decap_w0
xfeed_4997 0 1 decap_w0
xfeed_4996 0 1 decap_w0
xfeed_4995 0 1 decap_w0
xfeed_4994 0 1 decap_w0
xfeed_4993 0 1 decap_w0
xfeed_4991 0 1 decap_w0
xfeed_4990 0 1 decap_w0
xsubckt_673_or21nand_x0 0 1 88 1966 436 167 or21nand_x0
xsubckt_82_inv_x0 0 1 700 2008 inv_x0
xsubckt_84_inv_x0 0 1 698 2007 inv_x0
xfeed_12349 0 1 decap_w0
xfeed_12348 0 1 decap_w0
xfeed_12347 0 1 decap_w0
xfeed_12346 0 1 tie
xfeed_12345 0 1 decap_w0
xfeed_12344 0 1 decap_w0
xfeed_12343 0 1 decap_w0
xfeed_12342 0 1 decap_w0
xfeed_12341 0 1 decap_w0
xfeed_12340 0 1 decap_w0
xfeed_11819 0 1 decap_w0
xfeed_11818 0 1 decap_w0
xfeed_11817 0 1 decap_w0
xfeed_11816 0 1 decap_w0
xfeed_11815 0 1 decap_w0
xfeed_11814 0 1 tie
xfeed_11813 0 1 decap_w0
xfeed_11812 0 1 decap_w0
xfeed_11811 0 1 decap_w0
xfeed_11810 0 1 decap_w0
xsubckt_1041_mux2_x1 0 1 1857 1497 1949 1576 mux2_x1
xsubckt_731_nor3_x0 0 1 1733 1738 1737 1734 nor3_x0
xsubckt_634_and21nor_x0 0 1 124 752 449 410 and21nor_x0
xsubckt_1400_nand2_x0 0 1 1192 774 1978 nand2_x0
xcmpt_MOS6502_state_bit0_hfns_0 0 1 1924 1922 buf_x4
xcmpt_MOS6502_state_bit0_hfns_1 0 1 1923 1922 buf_x4
xcmpt_MOS6502_state_bit0_hfns_2 0 1 1922 1930 buf_x4
xdiode_209 0 1 1916 diode_w1
xdiode_208 0 1 1916 diode_w1
xdiode_207 0 1 661 diode_w1
xdiode_206 0 1 661 diode_w1
xdiode_205 0 1 661 diode_w1
xdiode_204 0 1 660 diode_w1
xdiode_203 0 1 660 diode_w1
xdiode_202 0 1 660 diode_w1
xdiode_201 0 1 775 diode_w1
xdiode_200 0 1 775 diode_w1
xfeed_9929 0 1 decap_w0
xfeed_9928 0 1 decap_w0
xfeed_9927 0 1 decap_w0
xfeed_9926 0 1 decap_w0
xfeed_9925 0 1 decap_w0
xfeed_9924 0 1 decap_w0
xfeed_9923 0 1 decap_w0
xfeed_9922 0 1 decap_w0
xfeed_9921 0 1 decap_w0
xfeed_9920 0 1 decap_w0
xfeed_6149 0 1 decap_w0
xfeed_6148 0 1 decap_w0
xfeed_6147 0 1 decap_w0
xfeed_6146 0 1 decap_w0
xfeed_6145 0 1 tie
xfeed_6144 0 1 decap_w0
xfeed_6143 0 1 decap_w0
xfeed_6142 0 1 decap_w0
xfeed_6141 0 1 decap_w0
xfeed_6140 0 1 decap_w0
xfeed_5619 0 1 decap_w0
xfeed_5618 0 1 decap_w0
xfeed_5616 0 1 decap_w0
xfeed_5615 0 1 decap_w0
xfeed_5614 0 1 decap_w0
xfeed_5613 0 1 decap_w0
xfeed_5612 0 1 decap_w0
xfeed_5611 0 1 decap_w0
xfeed_5610 0 1 decap_w0
xfeed_1309 0 1 decap_w0
xfeed_1308 0 1 decap_w0
xfeed_1307 0 1 decap_w0
xfeed_1306 0 1 decap_w0
xfeed_1305 0 1 decap_w0
xfeed_1304 0 1 decap_w0
xfeed_1303 0 1 decap_w0
xfeed_1302 0 1 decap_w0
xfeed_1301 0 1 decap_w0
xfeed_1300 0 1 decap_w0
xsubckt_702_nand4_x0 0 1 1762 1927 1925 711 674 nand4_x0
xsubckt_1804_and21nor_x0 0 1 791 850 847 853 and21nor_x0
xfeed_12359 0 1 decap_w0
xfeed_12358 0 1 decap_w0
xfeed_12357 0 1 decap_w0
xfeed_12356 0 1 decap_w0
xfeed_12355 0 1 decap_w0
xfeed_12354 0 1 decap_w0
xfeed_12353 0 1 decap_w0
xfeed_12352 0 1 decap_w0
xfeed_12351 0 1 decap_w0
xfeed_12350 0 1 tie
xfeed_11829 0 1 decap_w0
xfeed_11828 0 1 decap_w0
xfeed_11827 0 1 decap_w0
xfeed_11826 0 1 decap_w0
xfeed_11825 0 1 decap_w0
xfeed_11824 0 1 decap_w0
xfeed_11823 0 1 decap_w0
xfeed_11822 0 1 decap_w0
xfeed_11821 0 1 decap_w0
xfeed_11820 0 1 decap_w0
xsubckt_1220_nand2_x0 0 1 1344 284 1345 nand2_x0
xsubckt_1130_nand2_x0 0 1 1427 1940 2047 nand2_x0
xsubckt_1037_mux2_x1 0 1 1858 1506 1963 1510 mux2_x1
xsubckt_437_and4_x1 0 1 313 659 641 640 634 and4_x1
xsubckt_1639_or21nand_x0 0 1 955 1105 962 960 or21nand_x0
xdiode_219 0 1 1928 diode_w1
xdiode_218 0 1 1928 diode_w1
xdiode_217 0 1 1928 diode_w1
xdiode_216 0 1 1925 diode_w1
xdiode_215 0 1 1925 diode_w1
xdiode_214 0 1 1925 diode_w1
xdiode_213 0 1 1925 diode_w1
xdiode_212 0 1 1926 diode_w1
xdiode_211 0 1 1916 diode_w1
xdiode_210 0 1 1916 diode_w1
xfeed_9939 0 1 decap_w0
xfeed_9938 0 1 decap_w0
xfeed_9937 0 1 decap_w0
xfeed_9936 0 1 decap_w0
xfeed_9935 0 1 decap_w0
xfeed_9934 0 1 tie
xfeed_9933 0 1 decap_w0
xfeed_9932 0 1 decap_w0
xfeed_9931 0 1 decap_w0
xfeed_9930 0 1 decap_w0
xfeed_6159 0 1 decap_w0
xfeed_6158 0 1 decap_w0
xfeed_6157 0 1 tie
xfeed_6156 0 1 decap_w0
xfeed_6155 0 1 decap_w0
xfeed_6154 0 1 decap_w0
xfeed_6153 0 1 decap_w0
xfeed_6152 0 1 decap_w0
xfeed_6151 0 1 decap_w0
xfeed_6150 0 1 decap_w0
xfeed_5629 0 1 tie
xfeed_5628 0 1 decap_w0
xfeed_5627 0 1 decap_w0
xfeed_5626 0 1 decap_w0
xfeed_5625 0 1 decap_w0
xfeed_5624 0 1 decap_w0
xfeed_5623 0 1 decap_w0
xfeed_5622 0 1 tie
xfeed_5621 0 1 decap_w0
xfeed_5620 0 1 decap_w0
xfeed_1319 0 1 decap_w0
xfeed_1318 0 1 decap_w0
xfeed_1317 0 1 decap_w0
xfeed_1316 0 1 decap_w0
xfeed_1315 0 1 decap_w0
xfeed_1314 0 1 decap_w0
xfeed_1313 0 1 decap_w0
xfeed_1312 0 1 decap_w0
xfeed_1311 0 1 decap_w0
xfeed_1310 0 1 tie
xsubckt_1040_nand2_x0 0 1 1497 1499 1498 nand2_x0
xsubckt_361_inv_x0 0 1 29 388 inv_x0
xsubckt_1542_or21nand_x0 0 1 1052 1055 1122 90 or21nand_x0
xfeed_12369 0 1 decap_w0
xfeed_12368 0 1 decap_w0
xfeed_12367 0 1 decap_w0
xfeed_12366 0 1 decap_w0
xfeed_12365 0 1 decap_w0
xfeed_12364 0 1 decap_w0
xfeed_12363 0 1 decap_w0
xfeed_12362 0 1 decap_w0
xfeed_12361 0 1 decap_w0
xfeed_12360 0 1 decap_w0
xfeed_11839 0 1 decap_w0
xfeed_11838 0 1 decap_w0
xfeed_11837 0 1 decap_w0
xfeed_11836 0 1 decap_w0
xfeed_11835 0 1 decap_w0
xfeed_11834 0 1 decap_w0
xfeed_11833 0 1 decap_w0
xfeed_11832 0 1 decap_w0
xfeed_11831 0 1 decap_w0
xfeed_11830 0 1 decap_w0
xsubckt_1338_or21nand_x0 0 1 1249 1250 1322 759 or21nand_x0
xdiode_229 0 1 589 diode_w1
xdiode_228 0 1 589 diode_w1
xdiode_227 0 1 663 diode_w1
xdiode_226 0 1 663 diode_w1
xdiode_225 0 1 663 diode_w1
xdiode_224 0 1 1927 diode_w1
xdiode_223 0 1 1927 diode_w1
xdiode_222 0 1 1927 diode_w1
xdiode_221 0 1 1928 diode_w1
xdiode_220 0 1 1928 diode_w1
xfeed_9949 0 1 tie
xfeed_9948 0 1 decap_w0
xfeed_9947 0 1 decap_w0
xfeed_9946 0 1 decap_w0
xfeed_9945 0 1 decap_w0
xfeed_9944 0 1 decap_w0
xfeed_9943 0 1 decap_w0
xfeed_9942 0 1 decap_w0
xfeed_9941 0 1 tie
xfeed_9940 0 1 decap_w0
xfeed_6169 0 1 decap_w0
xfeed_6168 0 1 decap_w0
xfeed_6167 0 1 decap_w0
xfeed_6166 0 1 decap_w0
xfeed_6165 0 1 decap_w0
xfeed_6164 0 1 decap_w0
xfeed_6163 0 1 decap_w0
xfeed_6162 0 1 decap_w0
xfeed_6161 0 1 decap_w0
xfeed_6160 0 1 decap_w0
xfeed_5639 0 1 decap_w0
xfeed_5638 0 1 decap_w0
xfeed_5637 0 1 decap_w0
xfeed_5636 0 1 decap_w0
xfeed_5635 0 1 decap_w0
xfeed_5633 0 1 decap_w0
xfeed_5632 0 1 decap_w0
xfeed_5631 0 1 decap_w0
xfeed_5630 0 1 decap_w0
xfeed_1329 0 1 decap_w0
xfeed_1328 0 1 decap_w0
xfeed_1327 0 1 decap_w0
xfeed_1326 0 1 decap_w0
xfeed_1325 0 1 decap_w0
xfeed_1324 0 1 tie
xfeed_1323 0 1 decap_w0
xfeed_1322 0 1 decap_w0
xfeed_1321 0 1 decap_w0
xfeed_1320 0 1 tie
xsubckt_973_or21nand_x0 0 1 1869 1556 1553 1573 or21nand_x0
xsubckt_959_nand4_x0 0 1 1562 643 532 1576 1563 nand4_x0
xsubckt_873_nand3_x0 0 1 1610 1962 1964 2054 nand3_x0
xsubckt_266_nand2_x0 0 1 482 609 489 nand2_x0
xsubckt_367_and3_x1 0 1 382 652 526 383 and3_x1
xfeed_12379 0 1 decap_w0
xfeed_12378 0 1 decap_w0
xfeed_12377 0 1 decap_w0
xfeed_12376 0 1 decap_w0
xfeed_12375 0 1 decap_w0
xfeed_12374 0 1 decap_w0
xfeed_12373 0 1 decap_w0
xfeed_12372 0 1 decap_w0
xfeed_12371 0 1 decap_w0
xfeed_12370 0 1 decap_w0
xfeed_11849 0 1 decap_w0
xfeed_11848 0 1 decap_w0
xfeed_11847 0 1 decap_w0
xfeed_11846 0 1 decap_w0
xfeed_11845 0 1 decap_w0
xfeed_11844 0 1 decap_w0
xfeed_11843 0 1 decap_w0
xfeed_11842 0 1 tie
xfeed_11841 0 1 decap_w0
xfeed_11840 0 1 decap_w0
xsubckt_693_nand3_x0 0 1 1770 1775 1774 1771 nand3_x0
xsubckt_315_and2_x1 0 1 433 437 434 and2_x1
xsubckt_1387_nand2_x0 0 1 1204 775 1979 nand2_x0
xsubckt_1545_and4_x1 0 1 1049 1997 1128 1098 1097 and4_x1
xsubckt_1730_nand2_x0 0 1 864 1101 866 nand2_x0
xsubckt_1733_mux2_x1 0 1 861 901 863 1142 mux2_x1
xdiode_239 0 1 657 diode_w1
xdiode_238 0 1 657 diode_w1
xdiode_237 0 1 175 diode_w1
xdiode_236 0 1 175 diode_w1
xdiode_235 0 1 1749 diode_w1
xdiode_234 0 1 1749 diode_w1
xdiode_233 0 1 1749 diode_w1
xdiode_232 0 1 1749 diode_w1
xdiode_231 0 1 1749 diode_w1
xdiode_230 0 1 1749 diode_w1
xfeed_9959 0 1 decap_w0
xfeed_9958 0 1 decap_w0
xfeed_9957 0 1 decap_w0
xfeed_9956 0 1 decap_w0
xfeed_9955 0 1 decap_w0
xfeed_9954 0 1 decap_w0
xfeed_9953 0 1 decap_w0
xfeed_9952 0 1 decap_w0
xfeed_9951 0 1 decap_w0
xfeed_9950 0 1 decap_w0
xfeed_6179 0 1 decap_w0
xfeed_6178 0 1 decap_w0
xfeed_6177 0 1 decap_w0
xfeed_6176 0 1 tie
xfeed_6175 0 1 decap_w0
xfeed_6174 0 1 decap_w0
xfeed_6173 0 1 decap_w0
xfeed_6172 0 1 decap_w0
xfeed_6171 0 1 decap_w0
xfeed_6170 0 1 decap_w0
xfeed_5649 0 1 decap_w0
xfeed_5648 0 1 decap_w0
xfeed_5647 0 1 decap_w0
xfeed_5646 0 1 decap_w0
xfeed_5645 0 1 decap_w0
xfeed_5644 0 1 decap_w0
xfeed_5643 0 1 decap_w0
xfeed_5642 0 1 tie
xfeed_5641 0 1 decap_w0
xfeed_5640 0 1 decap_w0
xfeed_1339 0 1 decap_w0
xfeed_1338 0 1 decap_w0
xfeed_1337 0 1 decap_w0
xfeed_1336 0 1 decap_w0
xfeed_1335 0 1 decap_w0
xfeed_1334 0 1 decap_w0
xfeed_1333 0 1 decap_w0
xfeed_1332 0 1 decap_w0
xfeed_1331 0 1 tie
xfeed_1330 0 1 decap_w0
xsubckt_1202_and21nor_x0 0 1 1362 614 602 459 and21nor_x0
xsubckt_672_or21nand_x0 0 1 89 2047 601 163 or21nand_x0
xsubckt_275_and3_x1 0 1 473 1916 771 475 and3_x1
xsubckt_425_nand3_x0 0 1 324 610 557 460 nand3_x0
xfeed_12389 0 1 decap_w0
xfeed_12388 0 1 decap_w0
xfeed_12387 0 1 decap_w0
xfeed_12386 0 1 decap_w0
xfeed_12385 0 1 decap_w0
xfeed_12384 0 1 decap_w0
xfeed_12383 0 1 decap_w0
xfeed_12382 0 1 decap_w0
xfeed_12381 0 1 decap_w0
xfeed_12380 0 1 decap_w0
xfeed_11859 0 1 decap_w0
xfeed_11858 0 1 decap_w0
xfeed_11857 0 1 decap_w0
xfeed_11856 0 1 decap_w0
xfeed_11855 0 1 decap_w0
xfeed_11854 0 1 decap_w0
xfeed_11853 0 1 tie
xfeed_11852 0 1 decap_w0
xfeed_11851 0 1 decap_w0
xfeed_11850 0 1 decap_w0
xsubckt_1015_nand4_x0 0 1 1516 643 622 526 313 nand4_x0
xsubckt_942_nand4_x0 0 1 1575 1917 680 673 669 nand4_x0
xsubckt_335_nand3_x0 0 1 413 686 608 418 nand3_x0
xsubckt_1460_nand2_x0 0 1 1136 1955 548 nand2_x0
xsubckt_1538_or21nand_x0 0 1 1056 1635 1116 690 or21nand_x0
xdiode_249 0 1 1739 diode_w1
xdiode_248 0 1 1739 diode_w1
xdiode_247 0 1 1739 diode_w1
xdiode_246 0 1 447 diode_w1
xdiode_245 0 1 447 diode_w1
xdiode_244 0 1 447 diode_w1
xdiode_243 0 1 771 diode_w1
xdiode_242 0 1 771 diode_w1
xdiode_241 0 1 657 diode_w1
xdiode_240 0 1 657 diode_w1
xfeed_9969 0 1 decap_w0
xfeed_9968 0 1 decap_w0
xfeed_9967 0 1 decap_w0
xfeed_9966 0 1 decap_w0
xfeed_9965 0 1 decap_w0
xfeed_9964 0 1 decap_w0
xfeed_9963 0 1 decap_w0
xfeed_9962 0 1 decap_w0
xfeed_9961 0 1 decap_w0
xfeed_9960 0 1 decap_w0
xfeed_6188 0 1 decap_w0
xfeed_6187 0 1 decap_w0
xfeed_6185 0 1 decap_w0
xfeed_6184 0 1 decap_w0
xfeed_6183 0 1 decap_w0
xfeed_6182 0 1 decap_w0
xfeed_6181 0 1 decap_w0
xfeed_6180 0 1 tie
xfeed_5659 0 1 decap_w0
xfeed_5658 0 1 decap_w0
xfeed_5657 0 1 tie
xfeed_5656 0 1 decap_w0
xfeed_5655 0 1 decap_w0
xfeed_5654 0 1 decap_w0
xfeed_5653 0 1 decap_w0
xfeed_5652 0 1 decap_w0
xfeed_5651 0 1 decap_w0
xfeed_5650 0 1 decap_w0
xfeed_1349 0 1 decap_w0
xfeed_1348 0 1 decap_w0
xfeed_1347 0 1 decap_w0
xfeed_1346 0 1 decap_w0
xfeed_1345 0 1 decap_w0
xfeed_1344 0 1 decap_w0
xfeed_1343 0 1 tie
xfeed_1342 0 1 decap_w0
xfeed_1341 0 1 decap_w0
xfeed_1340 0 1 decap_w0
xsubckt_1137_or21nand_x0 0 1 1421 287 1625 1436 or21nand_x0
xsubckt_1066_and2_x1 0 1 1477 708 1575 and2_x1
xsubckt_776_nand2_x0 0 1 1694 1997 1746 nand2_x0
xsubckt_219_and2_x1 0 1 535 687 666 and2_x1
xfeed_13009 0 1 decap_w0
xfeed_13008 0 1 decap_w0
xfeed_13007 0 1 decap_w0
xfeed_13006 0 1 decap_w0
xfeed_13005 0 1 decap_w0
xfeed_13004 0 1 decap_w0
xfeed_13003 0 1 decap_w0
xfeed_13002 0 1 decap_w0
xfeed_13001 0 1 decap_w0
xfeed_13000 0 1 decap_w0
xfeed_12399 0 1 decap_w0
xfeed_12398 0 1 decap_w0
xfeed_12397 0 1 decap_w0
xfeed_12396 0 1 decap_w0
xfeed_12395 0 1 decap_w0
xfeed_12394 0 1 decap_w0
xfeed_12393 0 1 decap_w0
xfeed_12392 0 1 decap_w0
xfeed_12391 0 1 decap_w0
xfeed_12390 0 1 decap_w0
xfeed_11869 0 1 decap_w0
xfeed_11868 0 1 decap_w0
xfeed_11867 0 1 decap_w0
xfeed_11866 0 1 tie
xfeed_11865 0 1 decap_w0
xfeed_11864 0 1 decap_w0
xfeed_11863 0 1 decap_w0
xfeed_11862 0 1 decap_w0
xfeed_11861 0 1 tie
xfeed_11860 0 1 decap_w0
xsubckt_1114_mux2_x1 0 1 1843 2001 1992 1438 mux2_x1
xsubckt_686_nand2_x0 0 1 1777 1780 1779 nand2_x0
xsubckt_654_and2_x1 0 1 105 107 106 and2_x1
xsubckt_429_and21nor_x0 0 1 320 321 331 535 and21nor_x0
xsubckt_540_and3_x1 0 1 213 425 270 269 and3_x1
xsubckt_1294_and21nor_x0 0 1 1289 752 478 1317 and21nor_x0
xsubckt_1423_and2_x1 0 1 1170 1181 1172 and2_x1
xdiode_259 0 1 1745 diode_w1
xdiode_258 0 1 1745 diode_w1
xdiode_257 0 1 1745 diode_w1
xdiode_256 0 1 1740 diode_w1
xdiode_255 0 1 1740 diode_w1
xdiode_254 0 1 1740 diode_w1
xdiode_253 0 1 1740 diode_w1
xdiode_252 0 1 1739 diode_w1
xdiode_251 0 1 1739 diode_w1
xdiode_250 0 1 1739 diode_w1
xfeed_9979 0 1 decap_w0
xfeed_9978 0 1 decap_w0
xfeed_9977 0 1 decap_w0
xfeed_9976 0 1 decap_w0
xfeed_9975 0 1 decap_w0
xfeed_9974 0 1 decap_w0
xfeed_9973 0 1 decap_w0
xfeed_9972 0 1 decap_w0
xfeed_9971 0 1 decap_w0
xfeed_9970 0 1 decap_w0
xfeed_6199 0 1 decap_w0
xfeed_6197 0 1 tie
xfeed_6196 0 1 decap_w0
xfeed_6195 0 1 decap_w0
xfeed_6194 0 1 decap_w0
xfeed_6193 0 1 decap_w0
xfeed_6192 0 1 decap_w0
xfeed_6191 0 1 decap_w0
xfeed_6190 0 1 tie
xfeed_5669 0 1 decap_w0
xfeed_5668 0 1 decap_w0
xfeed_5667 0 1 tie
xfeed_5666 0 1 decap_w0
xfeed_5665 0 1 decap_w0
xfeed_5664 0 1 decap_w0
xfeed_5663 0 1 decap_w0
xfeed_5662 0 1 decap_w0
xfeed_5661 0 1 decap_w0
xfeed_5660 0 1 decap_w0
xfeed_1359 0 1 decap_w0
xfeed_1358 0 1 decap_w0
xfeed_1357 0 1 decap_w0
xfeed_1356 0 1 decap_w0
xfeed_1355 0 1 decap_w0
xfeed_1354 0 1 decap_w0
xfeed_1353 0 1 tie
xfeed_1352 0 1 decap_w0
xfeed_1351 0 1 decap_w0
xfeed_1350 0 1 decap_w0
xsubckt_1124_nor3_x0 0 1 1433 1940 1963 1956 nor3_x0
xsubckt_1008_nand3_x0 0 1 1521 643 533 1523 nand3_x0
xsubckt_971_and3_x1 0 1 1554 623 519 1567 and3_x1
xsubckt_562_and2_x1 0 1 193 456 403 and2_x1
xfeed_13019 0 1 decap_w0
xfeed_13018 0 1 decap_w0
xfeed_13017 0 1 decap_w0
xfeed_13016 0 1 decap_w0
xfeed_13015 0 1 decap_w0
xfeed_13014 0 1 decap_w0
xfeed_13013 0 1 decap_w0
xfeed_13012 0 1 decap_w0
xfeed_13011 0 1 decap_w0
xfeed_13010 0 1 tie
xfeed_11877 0 1 decap_w0
xfeed_11876 0 1 decap_w0
xfeed_11875 0 1 decap_w0
xfeed_11874 0 1 decap_w0
xfeed_11873 0 1 decap_w0
xfeed_11872 0 1 tie
xfeed_11871 0 1 decap_w0
xfeed_11870 0 1 decap_w0
xsubckt_1740_and3_x1 0 1 854 860 857 855 and3_x1
xdiode_267 0 1 711 diode_w1
xdiode_266 0 1 711 diode_w1
xdiode_265 0 1 1745 diode_w1
xdiode_264 0 1 1745 diode_w1
xdiode_263 0 1 1745 diode_w1
xdiode_262 0 1 1745 diode_w1
xdiode_261 0 1 1745 diode_w1
xdiode_260 0 1 1745 diode_w1
xfeed_11879 0 1 decap_w0
xfeed_11878 0 1 decap_w0
xfeed_9989 0 1 decap_w0
xfeed_9988 0 1 decap_w0
xfeed_9987 0 1 decap_w0
xfeed_9986 0 1 decap_w0
xfeed_9985 0 1 decap_w0
xfeed_9984 0 1 decap_w0
xfeed_9983 0 1 decap_w0
xfeed_9982 0 1 decap_w0
xfeed_9981 0 1 decap_w0
xfeed_9980 0 1 decap_w0
xfeed_5679 0 1 decap_w0
xfeed_5678 0 1 decap_w0
xfeed_5677 0 1 tie
xfeed_5676 0 1 decap_w0
xfeed_5675 0 1 decap_w0
xfeed_5674 0 1 decap_w0
xfeed_5673 0 1 decap_w0
xfeed_5672 0 1 decap_w0
xfeed_5671 0 1 decap_w0
xfeed_5670 0 1 decap_w0
xfeed_1369 0 1 decap_w0
xfeed_1368 0 1 tie
xfeed_1367 0 1 decap_w0
xfeed_1366 0 1 decap_w0
xfeed_1365 0 1 decap_w0
xfeed_1364 0 1 decap_w0
xfeed_1363 0 1 decap_w0
xfeed_1362 0 1 decap_w0
xfeed_1361 0 1 decap_w0
xfeed_1360 0 1 decap_w0
xsubckt_877_nexor2_x0 0 1 1606 1614 1607 nexor2_x0
xsubckt_558_and2_x1 0 1 197 551 543 and2_x1
xdiode_269 0 1 600 diode_w1
xdiode_268 0 1 711 diode_w1
xfeed_13029 0 1 decap_w0
xfeed_13028 0 1 decap_w0
xfeed_13027 0 1 decap_w0
xfeed_13026 0 1 decap_w0
xfeed_13025 0 1 decap_w0
xfeed_13024 0 1 decap_w0
xfeed_13023 0 1 decap_w0
xfeed_13022 0 1 decap_w0
xfeed_13021 0 1 decap_w0
xfeed_13020 0 1 decap_w0
xfeed_11884 0 1 decap_w0
xfeed_11883 0 1 decap_w0
xfeed_11882 0 1 decap_w0
xfeed_11881 0 1 decap_w0
xfeed_11880 0 1 decap_w0
xsubckt_1213_and3_x1 0 1 1351 205 1756 1354 and3_x1
xsubckt_1093_and21nor_x0 0 1 1454 386 1563 524 and21nor_x0
xsubckt_311_nand2_x0 0 1 437 557 439 nand2_x0
xsubckt_1327_and2_x1 0 1 1259 435 1260 and2_x1
xsubckt_1359_nand2_x0 0 1 1230 775 1967 nand2_x0
xsubckt_1612_nand2_x0 0 1 982 984 983 nand2_x0
xdiode_274 0 1 600 diode_w1
xdiode_273 0 1 600 diode_w1
xdiode_272 0 1 600 diode_w1
xdiode_271 0 1 600 diode_w1
xdiode_270 0 1 600 diode_w1
xfeed_11889 0 1 decap_w0
xfeed_11888 0 1 decap_w0
xfeed_11887 0 1 decap_w0
xfeed_11886 0 1 decap_w0
xfeed_11885 0 1 decap_w0
xfeed_9999 0 1 decap_w0
xfeed_9998 0 1 decap_w0
xfeed_9997 0 1 decap_w0
xfeed_9996 0 1 decap_w0
xfeed_9995 0 1 decap_w0
xfeed_9994 0 1 decap_w0
xfeed_9993 0 1 decap_w0
xfeed_9992 0 1 decap_w0
xfeed_9991 0 1 decap_w0
xfeed_9990 0 1 decap_w0
xfeed_5689 0 1 decap_w0
xfeed_5688 0 1 decap_w0
xfeed_5687 0 1 decap_w0
xfeed_5686 0 1 decap_w0
xfeed_5685 0 1 decap_w0
xfeed_5684 0 1 tie
xfeed_5683 0 1 decap_w0
xfeed_5682 0 1 decap_w0
xfeed_5681 0 1 decap_w0
xfeed_5680 0 1 decap_w0
xfeed_1379 0 1 decap_w0
xfeed_1378 0 1 decap_w0
xfeed_1377 0 1 decap_w0
xfeed_1376 0 1 decap_w0
xfeed_1375 0 1 tie
xfeed_1374 0 1 decap_w0
xfeed_1373 0 1 decap_w0
xfeed_1372 0 1 decap_w0
xfeed_1371 0 1 decap_w0
xfeed_1370 0 1 decap_w0
xsubckt_307_nand3_x0 0 1 441 687 609 447 nand3_x0
xsubckt_131_nand2_x0 0 1 637 660 639 nand2_x0
xsubckt_352_and3_x1 0 1 396 401 398 397 and3_x1
xsubckt_1850_dff_x1 0 1 2028 1888 35 dff_x1
xdiode_279 0 1 1964 diode_w1
xdiode_278 0 1 1964 diode_w1
xdiode_277 0 1 1964 diode_w1
xdiode_276 0 1 600 diode_w1
xdiode_275 0 1 600 diode_w1
xfeed_13039 0 1 decap_w0
xfeed_13038 0 1 decap_w0
xfeed_13037 0 1 decap_w0
xfeed_13036 0 1 decap_w0
xfeed_13035 0 1 decap_w0
xfeed_13034 0 1 decap_w0
xfeed_13033 0 1 decap_w0
xfeed_13032 0 1 decap_w0
xfeed_13031 0 1 decap_w0
xfeed_13030 0 1 decap_w0
xfeed_12509 0 1 decap_w0
xfeed_12508 0 1 decap_w0
xfeed_12507 0 1 decap_w0
xfeed_12506 0 1 decap_w0
xfeed_12505 0 1 decap_w0
xfeed_12504 0 1 decap_w0
xfeed_12503 0 1 decap_w0
xfeed_12502 0 1 decap_w0
xfeed_12501 0 1 decap_w0
xfeed_12500 0 1 decap_w0
xfeed_11891 0 1 decap_w0
xfeed_11890 0 1 decap_w0
xsubckt_748_nand2_x0 0 1 2098 1725 1719 nand2_x0
xsubckt_193_nor2_x0 0 1 565 570 567 nor2_x0
xsubckt_1852_dff_x1 0 1 2026 1886 32 dff_x1
xsubckt_1854_dff_x1 0 1 2024 1884 32 dff_x1
xsubckt_1856_dff_x1 0 1 2022 1882 32 dff_x1
xdiode_281 0 1 1334 diode_w1
xdiode_280 0 1 1964 diode_w1
xfeed_11899 0 1 decap_w0
xfeed_11898 0 1 decap_w0
xfeed_11897 0 1 decap_w0
xfeed_11896 0 1 decap_w0
xfeed_11895 0 1 decap_w0
xfeed_11894 0 1 decap_w0
xfeed_11893 0 1 decap_w0
xfeed_11892 0 1 decap_w0
xfeed_6309 0 1 decap_w0
xfeed_6308 0 1 decap_w0
xfeed_6307 0 1 decap_w0
xfeed_6306 0 1 decap_w0
xfeed_6305 0 1 decap_w0
xfeed_6304 0 1 decap_w0
xfeed_6303 0 1 decap_w0
xfeed_6302 0 1 tie
xfeed_6301 0 1 decap_w0
xfeed_6300 0 1 decap_w0
xfeed_5699 0 1 decap_w0
xfeed_5698 0 1 decap_w0
xfeed_5697 0 1 decap_w0
xfeed_5696 0 1 tie
xfeed_5695 0 1 decap_w0
xfeed_5694 0 1 decap_w0
xfeed_5693 0 1 decap_w0
xfeed_5692 0 1 decap_w0
xfeed_5691 0 1 decap_w0
xfeed_5690 0 1 decap_w0
xfeed_1389 0 1 decap_w0
xfeed_1388 0 1 decap_w0
xfeed_1387 0 1 decap_w0
xfeed_1386 0 1 decap_w0
xfeed_1385 0 1 decap_w0
xfeed_1384 0 1 decap_w0
xfeed_1383 0 1 decap_w0
xfeed_1382 0 1 tie
xfeed_1381 0 1 decap_w0
xfeed_1380 0 1 decap_w0
xsubckt_705_and3_x1 0 1 1759 211 1763 1760 and3_x1
xsubckt_658_nand2_x0 0 1 102 2032 175 nand2_x0
xsubckt_234_and4_x1 0 1 517 533 530 524 518 and4_x1
xsubckt_348_and3_x1 0 1 400 712 1926 405 and3_x1
xsubckt_1858_dff_x1 0 1 1984 1919 54 dff_x1
xdiode_288 0 1 599 diode_w1
xdiode_287 0 1 599 diode_w1
xdiode_286 0 1 599 diode_w1
xdiode_285 0 1 599 diode_w1
xdiode_284 0 1 1334 diode_w1
xdiode_283 0 1 1334 diode_w1
xdiode_282 0 1 1334 diode_w1
xfeed_13049 0 1 decap_w0
xfeed_13048 0 1 decap_w0
xfeed_13047 0 1 decap_w0
xfeed_13046 0 1 decap_w0
xfeed_13045 0 1 decap_w0
xfeed_13044 0 1 decap_w0
xfeed_13043 0 1 decap_w0
xfeed_13042 0 1 decap_w0
xfeed_13041 0 1 decap_w0
xfeed_13040 0 1 decap_w0
xfeed_12519 0 1 decap_w0
xfeed_12518 0 1 decap_w0
xfeed_12517 0 1 decap_w0
xfeed_12516 0 1 decap_w0
xfeed_12515 0 1 decap_w0
xfeed_12514 0 1 tie
xfeed_12513 0 1 decap_w0
xfeed_12512 0 1 decap_w0
xfeed_12511 0 1 decap_w0
xfeed_12510 0 1 decap_w0
xsubckt_968_or21nand_x0 0 1 1870 1558 1557 1573 or21nand_x0
xsubckt_771_or21nand_x0 0 1 1698 1700 1767 100 or21nand_x0
xsubckt_256_and3_x1 0 1 495 714 1928 589 and3_x1
xsubckt_173_or2_x1 0 1 585 2055 1921 or2_x1
xsubckt_464_nand4_x0 0 1 286 715 1925 711 599 nand4_x0
xfeed_6319 0 1 decap_w0
xfeed_6318 0 1 decap_w0
xfeed_6317 0 1 decap_w0
xfeed_6316 0 1 decap_w0
xfeed_6315 0 1 decap_w0
xfeed_6314 0 1 decap_w0
xfeed_6313 0 1 decap_w0
xfeed_6312 0 1 decap_w0
xfeed_6311 0 1 tie
xfeed_6310 0 1 decap_w0
xfeed_2009 0 1 decap_w0
xfeed_2008 0 1 decap_w0
xfeed_2007 0 1 decap_w0
xfeed_2006 0 1 decap_w0
xfeed_2005 0 1 decap_w0
xfeed_2004 0 1 decap_w0
xfeed_2003 0 1 decap_w0
xfeed_2002 0 1 decap_w0
xfeed_2001 0 1 decap_w0
xfeed_2000 0 1 decap_w0
xfeed_1399 0 1 tie
xfeed_1398 0 1 decap_w0
xfeed_1397 0 1 decap_w0
xfeed_1396 0 1 decap_w0
xfeed_1395 0 1 decap_w0
xfeed_1394 0 1 decap_w0
xfeed_1393 0 1 decap_w0
xfeed_1392 0 1 tie
xfeed_1391 0 1 decap_w0
xfeed_1390 0 1 decap_w0
xsubckt_727_and2_x1 0 1 1737 2053 1748 and2_x1
xsubckt_641_nand2_x0 0 1 118 2033 175 nand2_x0
xsubckt_374_nand4_x0 0 1 375 532 530 518 384 nand4_x0
xsubckt_1411_nand3_x0 0 1 1181 1207 1196 1184 nand3_x0
xsubckt_1540_or21nand_x0 0 1 1054 1057 1118 760 or21nand_x0
xfeed_13059 0 1 decap_w0
xfeed_13058 0 1 decap_w0
xfeed_13057 0 1 decap_w0
xfeed_13056 0 1 tie
xfeed_13055 0 1 decap_w0
xfeed_13054 0 1 decap_w0
xfeed_13053 0 1 decap_w0
xfeed_13052 0 1 decap_w0
xfeed_13051 0 1 tie
xfeed_13050 0 1 decap_w0
xfeed_12529 0 1 decap_w0
xfeed_12528 0 1 decap_w0
xfeed_12527 0 1 decap_w0
xfeed_12526 0 1 tie
xfeed_12525 0 1 decap_w0
xfeed_12524 0 1 decap_w0
xfeed_12523 0 1 decap_w0
xfeed_12522 0 1 decap_w0
xfeed_12521 0 1 decap_w0
xfeed_12520 0 1 decap_w0
xsubckt_1099_and3_x1 0 1 1448 623 621 519 and3_x1
xsubckt_278_and2_x1 0 1 470 480 471 and2_x1
xsubckt_190_and2_x1 0 1 568 1925 1926 and2_x1
xsubckt_1737_or21nand_x0 0 1 857 859 861 1075 or21nand_x0
xfeed_6329 0 1 decap_w0
xfeed_6328 0 1 decap_w0
xfeed_6327 0 1 decap_w0
xfeed_6326 0 1 decap_w0
xfeed_6325 0 1 decap_w0
xfeed_6324 0 1 decap_w0
xfeed_6323 0 1 decap_w0
xfeed_6322 0 1 decap_w0
xfeed_6321 0 1 decap_w0
xfeed_6320 0 1 tie
xfeed_2019 0 1 tie
xfeed_2018 0 1 decap_w0
xfeed_2017 0 1 decap_w0
xfeed_2016 0 1 decap_w0
xfeed_2015 0 1 decap_w0
xfeed_2014 0 1 decap_w0
xfeed_2013 0 1 decap_w0
xfeed_2012 0 1 decap_w0
xfeed_2011 0 1 decap_w0
xfeed_2010 0 1 decap_w0
xsubckt_832_and21nor_x0 0 1 1645 691 1755 1754 and21nor_x0
xsubckt_91_inv_x0 0 1 2001 694 inv_x0
xsubckt_93_inv_x0 0 1 2000 693 inv_x0
xsubckt_461_nand2_x0 0 1 289 314 290 nand2_x0
xsubckt_1342_and4_x1 0 1 1245 1273 1266 1257 1247 and4_x1
xsubckt_1482_and2_x1 0 1 1114 1628 1115 and2_x1
xsubckt_1618_mux2_x1 0 1 976 1021 978 1142 mux2_x1
xfeed_13069 0 1 decap_w0
xfeed_13068 0 1 decap_w0
xfeed_13067 0 1 decap_w0
xfeed_13066 0 1 decap_w0
xfeed_13065 0 1 decap_w0
xfeed_13064 0 1 decap_w0
xfeed_13063 0 1 tie
xfeed_13062 0 1 decap_w0
xfeed_13061 0 1 decap_w0
xfeed_13060 0 1 decap_w0
xfeed_12539 0 1 decap_w0
xfeed_12538 0 1 decap_w0
xfeed_12537 0 1 decap_w0
xfeed_12536 0 1 decap_w0
xfeed_12535 0 1 decap_w0
xfeed_12534 0 1 decap_w0
xfeed_12533 0 1 tie
xfeed_12532 0 1 decap_w0
xfeed_12531 0 1 decap_w0
xfeed_12530 0 1 decap_w0
xsubckt_95_inv_x0 0 1 1999 692 inv_x0
xsubckt_97_inv_x0 0 1 1998 691 inv_x0
xsubckt_99_inv_x0 0 1 1997 690 inv_x0
xsubckt_103_nand2_x0 0 1 684 1916 771 nand2_x0
xsubckt_1601_and21nor_x0 0 1 993 994 1117 2049 and21nor_x0
xsubckt_1672_nand2_x0 0 1 922 1105 924 nand2_x0
xfeed_6339 0 1 decap_w0
xfeed_6338 0 1 decap_w0
xfeed_6337 0 1 decap_w0
xfeed_6336 0 1 decap_w0
xfeed_6335 0 1 decap_w0
xfeed_6334 0 1 decap_w0
xfeed_6333 0 1 decap_w0
xfeed_6332 0 1 decap_w0
xfeed_6331 0 1 decap_w0
xfeed_6330 0 1 decap_w0
xfeed_5809 0 1 decap_w0
xfeed_5808 0 1 decap_w0
xfeed_5807 0 1 decap_w0
xfeed_5806 0 1 tie
xfeed_5805 0 1 decap_w0
xfeed_5804 0 1 decap_w0
xfeed_5803 0 1 decap_w0
xfeed_5802 0 1 decap_w0
xfeed_5801 0 1 decap_w0
xfeed_5800 0 1 decap_w0
xfeed_2029 0 1 decap_w0
xfeed_2028 0 1 decap_w0
xfeed_2027 0 1 decap_w0
xfeed_2026 0 1 decap_w0
xfeed_2025 0 1 decap_w0
xfeed_2024 0 1 decap_w0
xfeed_2023 0 1 decap_w0
xfeed_2022 0 1 decap_w0
xfeed_2021 0 1 decap_w0
xfeed_2020 0 1 decap_w0
xsubckt_898_nand2_x0 0 1 1589 760 1591 nand2_x0
xsubckt_767_or21nand_x0 0 1 1702 2060 1742 1740 or21nand_x0
xsubckt_543_and2_x1 0 1 211 449 410 and2_x1
xsubckt_1300_nand4_x0 0 1 1283 1311 1303 1293 1285 nand4_x0
xsubckt_1314_nand2_x0 0 1 1271 775 1971 nand2_x0
xfeed_13079 0 1 decap_w0
xfeed_13078 0 1 decap_w0
xfeed_13077 0 1 decap_w0
xfeed_13076 0 1 decap_w0
xfeed_13075 0 1 decap_w0
xfeed_13074 0 1 decap_w0
xfeed_13073 0 1 decap_w0
xfeed_13072 0 1 decap_w0
xfeed_13071 0 1 decap_w0
xfeed_13070 0 1 decap_w0
xfeed_12549 0 1 decap_w0
xfeed_12548 0 1 decap_w0
xfeed_12547 0 1 decap_w0
xfeed_12546 0 1 decap_w0
xfeed_12545 0 1 decap_w0
xfeed_12544 0 1 decap_w0
xfeed_12543 0 1 decap_w0
xfeed_12542 0 1 decap_w0
xfeed_12541 0 1 decap_w0
xfeed_12540 0 1 decap_w0
xsubckt_366_or21nand_x0 0 1 383 660 624 521 or21nand_x0
xsubckt_539_and2_x1 0 1 214 515 374 and2_x1
xfeed_6349 0 1 decap_w0
xfeed_6348 0 1 decap_w0
xfeed_6347 0 1 decap_w0
xfeed_6346 0 1 decap_w0
xfeed_6345 0 1 decap_w0
xfeed_6344 0 1 decap_w0
xfeed_6342 0 1 decap_w0
xfeed_6341 0 1 decap_w0
xfeed_6340 0 1 decap_w0
xfeed_5819 0 1 decap_w0
xfeed_5818 0 1 tie
xfeed_5817 0 1 decap_w0
xfeed_5816 0 1 decap_w0
xfeed_5815 0 1 decap_w0
xfeed_5814 0 1 decap_w0
xfeed_5813 0 1 decap_w0
xfeed_5812 0 1 decap_w0
xfeed_5811 0 1 tie
xfeed_5810 0 1 decap_w0
xfeed_2039 0 1 decap_w0
xfeed_2038 0 1 decap_w0
xfeed_2037 0 1 decap_w0
xfeed_2036 0 1 tie
xfeed_2035 0 1 decap_w0
xfeed_2034 0 1 decap_w0
xfeed_2033 0 1 decap_w0
xfeed_2032 0 1 decap_w0
xfeed_2031 0 1 decap_w0
xfeed_2030 0 1 decap_w0
xfeed_1509 0 1 decap_w0
xfeed_1508 0 1 decap_w0
xfeed_1507 0 1 decap_w0
xfeed_1506 0 1 decap_w0
xfeed_1505 0 1 decap_w0
xfeed_1504 0 1 decap_w0
xfeed_1503 0 1 decap_w0
xfeed_1502 0 1 decap_w0
xfeed_1501 0 1 decap_w0
xfeed_1500 0 1 decap_w0
xsubckt_974_and2_x1 0 1 1552 645 533 and2_x1
xsubckt_860_and3_x1 0 1 1621 200 1762 1622 and3_x1
xsubckt_1741_nand3_x0 0 1 853 860 857 855 nand3_x0
xfeed_13089 0 1 decap_w0
xfeed_13088 0 1 decap_w0
xfeed_13087 0 1 decap_w0
xfeed_13086 0 1 decap_w0
xfeed_13085 0 1 decap_w0
xfeed_13084 0 1 decap_w0
xfeed_13083 0 1 decap_w0
xfeed_13082 0 1 tie
xfeed_13081 0 1 decap_w0
xfeed_13080 0 1 decap_w0
xfeed_12559 0 1 decap_w0
xfeed_12558 0 1 decap_w0
xfeed_12557 0 1 decap_w0
xfeed_12556 0 1 decap_w0
xfeed_12555 0 1 decap_w0
xfeed_12554 0 1 decap_w0
xfeed_12553 0 1 decap_w0
xfeed_12552 0 1 decap_w0
xfeed_12551 0 1 decap_w0
xfeed_12550 0 1 decap_w0
xsubckt_1268_and3_x1 0 1 1312 1324 1315 1313 and3_x1
xsubckt_967_nand3_x0 0 1 1557 622 520 1567 nand3_x0
xsubckt_828_and21nor_x0 0 1 1648 743 600 1745 and21nor_x0
xsubckt_1693_and21nor_x0 0 1 901 902 1121 152 and21nor_x0
xfeed_6359 0 1 decap_w0
xfeed_6358 0 1 decap_w0
xfeed_6357 0 1 decap_w0
xfeed_6356 0 1 decap_w0
xfeed_6355 0 1 decap_w0
xfeed_6354 0 1 decap_w0
xfeed_6353 0 1 decap_w0
xfeed_6352 0 1 decap_w0
xfeed_6351 0 1 decap_w0
xfeed_6350 0 1 decap_w0
xfeed_5829 0 1 decap_w0
xfeed_5828 0 1 decap_w0
xfeed_5827 0 1 decap_w0
xfeed_5826 0 1 decap_w0
xfeed_5825 0 1 tie
xfeed_5824 0 1 decap_w0
xfeed_5823 0 1 decap_w0
xfeed_5822 0 1 decap_w0
xfeed_5821 0 1 decap_w0
xfeed_5820 0 1 decap_w0
xfeed_2049 0 1 decap_w0
xfeed_2048 0 1 tie
xfeed_2047 0 1 decap_w0
xfeed_2046 0 1 decap_w0
xfeed_2045 0 1 decap_w0
xfeed_2044 0 1 decap_w0
xfeed_2043 0 1 decap_w0
xfeed_2042 0 1 decap_w0
xfeed_2041 0 1 decap_w0
xfeed_2040 0 1 decap_w0
xfeed_1519 0 1 decap_w0
xfeed_1518 0 1 decap_w0
xfeed_1517 0 1 decap_w0
xfeed_1516 0 1 decap_w0
xfeed_1515 0 1 decap_w0
xfeed_1514 0 1 decap_w0
xfeed_1513 0 1 decap_w0
xfeed_1512 0 1 decap_w0
xfeed_1511 0 1 decap_w0
xfeed_1510 0 1 decap_w0
xsubckt_1102_and3_x1 0 1 1445 1455 1453 1446 and3_x1
xsubckt_930_mux2_x1 0 1 1887 2027 1605 1578 mux2_x1
xsubckt_1471_nand3_x0 0 1 1125 1142 1137 1126 nand3_x0
xfeed_13099 0 1 decap_w0
xfeed_13098 0 1 decap_w0
xfeed_13097 0 1 decap_w0
xfeed_13096 0 1 decap_w0
xfeed_13095 0 1 decap_w0
xfeed_13094 0 1 decap_w0
xfeed_13093 0 1 decap_w0
xfeed_13092 0 1 decap_w0
xfeed_13091 0 1 decap_w0
xfeed_13090 0 1 decap_w0
xfeed_12569 0 1 decap_w0
xfeed_12568 0 1 decap_w0
xfeed_12567 0 1 decap_w0
xfeed_12566 0 1 decap_w0
xfeed_12565 0 1 tie
xfeed_12564 0 1 decap_w0
xfeed_12563 0 1 decap_w0
xfeed_12562 0 1 decap_w0
xfeed_12561 0 1 decap_w0
xfeed_12560 0 1 decap_w0
xsubckt_1088_and21nor_x0 0 1 1849 1462 1458 1576 and21nor_x0
xsubckt_926_mux2_x1 0 1 1890 1581 2030 1579 mux2_x1
xsubckt_241_and3_x1 0 1 510 560 540 511 and3_x1
xsubckt_1736_or21nand_x0 0 1 858 1067 869 1072 or21nand_x0
xfeed_6369 0 1 decap_w0
xfeed_6368 0 1 decap_w0
xfeed_6366 0 1 decap_w0
xfeed_6365 0 1 tie
xfeed_6364 0 1 decap_w0
xfeed_6363 0 1 decap_w0
xfeed_6362 0 1 decap_w0
xfeed_6361 0 1 decap_w0
xfeed_6360 0 1 decap_w0
xfeed_5839 0 1 decap_w0
xfeed_5838 0 1 decap_w0
xfeed_5837 0 1 decap_w0
xfeed_5836 0 1 decap_w0
xfeed_5835 0 1 decap_w0
xfeed_5834 0 1 decap_w0
xfeed_5833 0 1 decap_w0
xfeed_5832 0 1 decap_w0
xfeed_5831 0 1 decap_w0
xfeed_5830 0 1 decap_w0
xfeed_2059 0 1 decap_w0
xfeed_2058 0 1 decap_w0
xfeed_2057 0 1 decap_w0
xfeed_2056 0 1 tie
xfeed_2055 0 1 decap_w0
xfeed_2054 0 1 decap_w0
xfeed_2053 0 1 decap_w0
xfeed_2052 0 1 decap_w0
xfeed_2051 0 1 decap_w0
xfeed_2050 0 1 decap_w0
xfeed_1529 0 1 decap_w0
xfeed_1528 0 1 decap_w0
xfeed_1527 0 1 decap_w0
xfeed_1526 0 1 decap_w0
xfeed_1525 0 1 decap_w0
xfeed_1524 0 1 decap_w0
xfeed_1523 0 1 decap_w0
xfeed_1522 0 1 decap_w0
xfeed_1521 0 1 decap_w0
xfeed_1520 0 1 decap_w0
xsubckt_950_nand3_x0 0 1 1569 653 525 383 nand3_x0
xsubckt_666_or21nand_x0 0 1 2077 95 100 206 or21nand_x0
xsubckt_253_nand2_x0 0 1 498 679 571 nand2_x0
xsubckt_403_mux2_x1 0 1 346 348 347 1953 mux2_x1
xfeed_12577 0 1 decap_w0
xfeed_12576 0 1 decap_w0
xfeed_12575 0 1 decap_w0
xfeed_12574 0 1 decap_w0
xfeed_12573 0 1 decap_w0
xfeed_12572 0 1 decap_w0
xfeed_12571 0 1 decap_w0
xfeed_12570 0 1 decap_w0
xsubckt_1246_mux2_x1 0 1 1815 2099 2066 1334 mux2_x1
xsubckt_263_and2_x1 0 1 485 609 495 and2_x1
xsubckt_339_nand3_x0 0 1 409 682 558 421 nand3_x0
xsubckt_1529_and3_x1 0 1 1064 1099 1095 1070 and3_x1
xsubckt_1554_nand2_x0 0 1 1040 1101 1042 nand2_x0
xfeed_12579 0 1 decap_w0
xfeed_12578 0 1 decap_w0
xfeed_6379 0 1 decap_w0
xfeed_6378 0 1 decap_w0
xfeed_6377 0 1 decap_w0
xfeed_6376 0 1 decap_w0
xfeed_6375 0 1 decap_w0
xfeed_6374 0 1 decap_w0
xfeed_6373 0 1 decap_w0
xfeed_6372 0 1 decap_w0
xfeed_6371 0 1 decap_w0
xfeed_6370 0 1 tie
xfeed_5849 0 1 decap_w0
xfeed_5848 0 1 decap_w0
xfeed_5847 0 1 decap_w0
xfeed_5846 0 1 decap_w0
xfeed_5845 0 1 decap_w0
xfeed_5844 0 1 decap_w0
xfeed_5843 0 1 decap_w0
xfeed_5842 0 1 decap_w0
xfeed_5841 0 1 decap_w0
xfeed_5840 0 1 decap_w0
xfeed_2069 0 1 decap_w0
xfeed_2068 0 1 decap_w0
xfeed_2067 0 1 decap_w0
xfeed_2066 0 1 decap_w0
xfeed_2065 0 1 decap_w0
xfeed_2064 0 1 decap_w0
xfeed_2063 0 1 decap_w0
xfeed_2062 0 1 decap_w0
xfeed_2061 0 1 decap_w0
xfeed_2060 0 1 decap_w0
xfeed_1539 0 1 decap_w0
xfeed_1538 0 1 decap_w0
xfeed_1537 0 1 decap_w0
xfeed_1536 0 1 decap_w0
xfeed_1535 0 1 decap_w0
xfeed_1534 0 1 decap_w0
xfeed_1533 0 1 tie
xfeed_1532 0 1 decap_w0
xfeed_1531 0 1 decap_w0
xfeed_1530 0 1 decap_w0
xsubckt_680_nand3_x0 0 1 1783 2014 184 177 nand3_x0
xsubckt_249_nand3_x0 0 1 502 687 617 603 nand3_x0
xsubckt_159_nand3_x0 0 1 602 1929 715 670 nand3_x0
xsubckt_1374_nand2_x0 0 1 1216 1980 1316 nand2_x0
xfeed_12584 0 1 decap_w0
xfeed_12583 0 1 decap_w0
xfeed_12582 0 1 decap_w0
xfeed_12581 0 1 decap_w0
xfeed_12580 0 1 decap_w0
xsubckt_943_nand2_x0 0 1 1574 1940 1575 nand2_x0
xsubckt_1677_mux2_x1 0 1 917 922 920 929 mux2_x1
xfeed_12589 0 1 decap_w0
xfeed_12588 0 1 decap_w0
xfeed_12587 0 1 decap_w0
xfeed_12586 0 1 tie
xfeed_12585 0 1 decap_w0
xfeed_6389 0 1 decap_w0
xfeed_6388 0 1 decap_w0
xfeed_6387 0 1 decap_w0
xfeed_6386 0 1 decap_w0
xfeed_6385 0 1 decap_w0
xfeed_6384 0 1 decap_w0
xfeed_6383 0 1 decap_w0
xfeed_6382 0 1 decap_w0
xfeed_6381 0 1 decap_w0
xfeed_6380 0 1 decap_w0
xfeed_5858 0 1 decap_w0
xfeed_5857 0 1 decap_w0
xfeed_5856 0 1 decap_w0
xfeed_5855 0 1 tie
xfeed_5854 0 1 decap_w0
xfeed_5853 0 1 decap_w0
xfeed_5852 0 1 decap_w0
xfeed_5851 0 1 decap_w0
xfeed_5850 0 1 decap_w0
xfeed_2079 0 1 decap_w0
xfeed_2078 0 1 decap_w0
xfeed_2077 0 1 decap_w0
xfeed_2076 0 1 decap_w0
xfeed_2075 0 1 decap_w0
xfeed_2074 0 1 decap_w0
xfeed_2073 0 1 tie
xfeed_2072 0 1 decap_w0
xfeed_2071 0 1 decap_w0
xfeed_2070 0 1 decap_w0
xfeed_1549 0 1 decap_w0
xfeed_1548 0 1 decap_w0
xfeed_1547 0 1 decap_w0
xfeed_1546 0 1 decap_w0
xfeed_1545 0 1 decap_w0
xfeed_1544 0 1 decap_w0
xfeed_1543 0 1 decap_w0
xfeed_1542 0 1 decap_w0
xfeed_1541 0 1 decap_w0
xfeed_1540 0 1 tie
xsubckt_502_and3_x1 0 1 249 254 253 250 and3_x1
xcmpt_RDY_hfns_0 0 1 1917 1915 buf_x4
xcmpt_RDY_hfns_1 0 1 1916 1915 buf_x4
xcmpt_RDY_hfns_2 0 1 1915 1918 buf_x4
xdiode_19 0 1 679 diode_w1
xdiode_18 0 1 679 diode_w1
xdiode_17 0 1 679 diode_w1
xdiode_16 0 1 679 diode_w1
xdiode_15 0 1 679 diode_w1
xdiode_14 0 1 678 diode_w1
xdiode_13 0 1 678 diode_w1
xdiode_12 0 1 678 diode_w1
xdiode_11 0 1 678 diode_w1
xdiode_10 0 1 610 diode_w1
xfeed_13209 0 1 decap_w0
xfeed_13208 0 1 decap_w0
xfeed_13207 0 1 decap_w0
xfeed_13206 0 1 decap_w0
xfeed_13205 0 1 decap_w0
xfeed_13204 0 1 decap_w0
xfeed_13203 0 1 decap_w0
xfeed_13202 0 1 decap_w0
xfeed_13201 0 1 decap_w0
xfeed_13200 0 1 decap_w0
xfeed_12591 0 1 decap_w0
xfeed_12590 0 1 decap_w0
xsubckt_410_and3_x1 0 1 339 679 558 490 and3_x1
xsubckt_524_and2_x1 0 1 228 278 229 and2_x1
xsubckt_1443_nand3_x0 0 1 1152 2066 666 657 nand3_x0
xfeed_12599 0 1 decap_w0
xfeed_12598 0 1 decap_w0
xfeed_12597 0 1 decap_w0
xfeed_12596 0 1 decap_w0
xfeed_12595 0 1 decap_w0
xfeed_12594 0 1 decap_w0
xfeed_12593 0 1 decap_w0
xfeed_12592 0 1 decap_w0
xfeed_7009 0 1 decap_w0
xfeed_7008 0 1 decap_w0
xfeed_7007 0 1 decap_w0
xfeed_7006 0 1 decap_w0
xfeed_7005 0 1 decap_w0
xfeed_7004 0 1 tie
xfeed_7003 0 1 decap_w0
xfeed_7002 0 1 decap_w0
xfeed_7001 0 1 decap_w0
xfeed_7000 0 1 tie
xfeed_6399 0 1 decap_w0
xfeed_6398 0 1 decap_w0
xfeed_6397 0 1 decap_w0
xfeed_6396 0 1 decap_w0
xfeed_6395 0 1 decap_w0
xfeed_6394 0 1 tie
xfeed_6393 0 1 decap_w0
xfeed_6392 0 1 decap_w0
xfeed_6391 0 1 decap_w0
xfeed_6390 0 1 decap_w0
xfeed_5869 0 1 decap_w0
xfeed_5868 0 1 decap_w0
xfeed_5867 0 1 decap_w0
xfeed_5866 0 1 decap_w0
xfeed_5865 0 1 decap_w0
xfeed_5864 0 1 decap_w0
xfeed_5863 0 1 decap_w0
xfeed_5862 0 1 decap_w0
xfeed_5861 0 1 decap_w0
xfeed_2089 0 1 decap_w0
xfeed_2088 0 1 decap_w0
xfeed_2087 0 1 decap_w0
xfeed_2086 0 1 decap_w0
xfeed_2085 0 1 decap_w0
xfeed_2084 0 1 decap_w0
xfeed_2083 0 1 decap_w0
xfeed_2082 0 1 tie
xfeed_2081 0 1 decap_w0
xfeed_2080 0 1 decap_w0
xfeed_1559 0 1 decap_w0
xfeed_1558 0 1 decap_w0
xfeed_1557 0 1 decap_w0
xfeed_1556 0 1 decap_w0
xfeed_1555 0 1 decap_w0
xfeed_1554 0 1 decap_w0
xfeed_1553 0 1 tie
xfeed_1552 0 1 decap_w0
xfeed_1551 0 1 decap_w0
xfeed_1550 0 1 decap_w0
xsubckt_138_nand4_x0 0 1 630 660 639 636 635 nand4_x0
xsubckt_1488_and21nor_x0 0 1 1108 665 598 681 and21nor_x0
xsubckt_1493_mux2_x1 0 1 1103 1107 738 1143 mux2_x1
xdiode_29 0 1 682 diode_w1
xdiode_28 0 1 681 diode_w1
xdiode_27 0 1 681 diode_w1
xdiode_26 0 1 681 diode_w1
xdiode_25 0 1 680 diode_w1
xdiode_24 0 1 680 diode_w1
xdiode_23 0 1 680 diode_w1
xdiode_22 0 1 679 diode_w1
xdiode_21 0 1 679 diode_w1
xdiode_20 0 1 679 diode_w1
xfeed_13219 0 1 decap_w0
xfeed_13218 0 1 decap_w0
xfeed_13217 0 1 tie
xfeed_13216 0 1 decap_w0
xfeed_13215 0 1 decap_w0
xfeed_13214 0 1 decap_w0
xfeed_13213 0 1 decap_w0
xfeed_13212 0 1 decap_w0
xfeed_13211 0 1 decap_w0
xfeed_13210 0 1 decap_w0
xsubckt_1259_nand4_x0 0 1 1321 605 493 476 1756 nand4_x0
xsubckt_1227_and4_x1 0 1 1337 203 1353 1341 1338 and4_x1
xsubckt_406_and3_x1 0 1 343 687 678 595 and3_x1
xsubckt_1901_dff_x1 0 1 1986 1846 67 dff_x1
xfeed_7019 0 1 decap_w0
xfeed_7018 0 1 decap_w0
xfeed_7017 0 1 tie
xfeed_7016 0 1 decap_w0
xfeed_7015 0 1 decap_w0
xfeed_7014 0 1 decap_w0
xfeed_7013 0 1 decap_w0
xfeed_7012 0 1 decap_w0
xfeed_7011 0 1 decap_w0
xfeed_7010 0 1 decap_w0
xfeed_5876 0 1 decap_w0
xfeed_5875 0 1 decap_w0
xfeed_5874 0 1 tie
xfeed_5873 0 1 decap_w0
xfeed_5872 0 1 decap_w0
xfeed_5871 0 1 decap_w0
xfeed_5870 0 1 decap_w0
xfeed_2099 0 1 decap_w0
xfeed_2098 0 1 decap_w0
xfeed_2097 0 1 decap_w0
xfeed_2096 0 1 decap_w0
xfeed_2095 0 1 decap_w0
xfeed_2094 0 1 decap_w0
xfeed_2093 0 1 decap_w0
xfeed_2092 0 1 decap_w0
xfeed_2091 0 1 decap_w0
xfeed_2090 0 1 decap_w0
xfeed_1569 0 1 decap_w0
xfeed_1568 0 1 decap_w0
xfeed_1567 0 1 decap_w0
xfeed_1566 0 1 tie
xfeed_1565 0 1 decap_w0
xfeed_1564 0 1 decap_w0
xfeed_1563 0 1 decap_w0
xfeed_1562 0 1 decap_w0
xfeed_1561 0 1 decap_w0
xfeed_1560 0 1 decap_w0
xsubckt_211_nand4_x0 0 1 543 712 1926 674 670 nand4_x0
xsubckt_489_nand3_x0 0 1 27 315 271 262 nand3_x0
xsubckt_1724_and2_x1 0 1 870 873 871 and2_x1
xsubckt_1903_dff_x1 0 1 1993 1844 67 dff_x1
xsubckt_1905_dff_x1 0 1 1991 1842 67 dff_x1
xsubckt_1907_dff_x1 0 1 1989 1840 67 dff_x1
xspare_feed_100 0 1 tie
xspare_feed_101 0 1 tie
xspare_feed_102 0 1 decap_w0
xspare_feed_103 0 1 tie
xspare_feed_104 0 1 tie
xspare_feed_105 0 1 decap_w0
xspare_feed_106 0 1 tie
xspare_feed_107 0 1 tie
xspare_feed_108 0 1 decap_w0
xspare_feed_109 0 1 tie
xdiode_39 0 1 1575 diode_w1
xdiode_38 0 1 435 diode_w1
xdiode_37 0 1 435 diode_w1
xdiode_36 0 1 435 diode_w1
xdiode_35 0 1 435 diode_w1
xdiode_34 0 1 682 diode_w1
xdiode_33 0 1 682 diode_w1
xdiode_32 0 1 682 diode_w1
xdiode_31 0 1 682 diode_w1
xdiode_30 0 1 682 diode_w1
xfeed_13229 0 1 decap_w0
xfeed_13228 0 1 decap_w0
xfeed_13227 0 1 decap_w0
xfeed_13226 0 1 decap_w0
xfeed_13225 0 1 decap_w0
xfeed_13224 0 1 tie
xfeed_13223 0 1 decap_w0
xfeed_13222 0 1 decap_w0
xfeed_13221 0 1 decap_w0
xfeed_13220 0 1 decap_w0
xfeed_5879 0 1 tie
xfeed_5878 0 1 decap_w0
xfeed_5877 0 1 decap_w0
xsubckt_911_mux2_x1 0 1 1904 1612 2044 1580 mux2_x1
xsubckt_399_nand3_x0 0 1 350 617 558 489 nand3_x0
xsubckt_1346_nand2_x0 0 1 1242 774 1968 nand2_x0
xsubckt_1436_nand2_x0 0 1 1158 1169 1159 nand2_x0
xsubckt_1861_dff_x1 0 1 1952 1878 67 dff_x1
xsubckt_1863_dff_x1 0 1 1941 1876 67 dff_x1
xsubckt_1909_dff_x1 0 1 1987 1838 67 dff_x1
xfeed_7029 0 1 decap_w0
xfeed_7028 0 1 decap_w0
xfeed_7027 0 1 decap_w0
xfeed_7026 0 1 decap_w0
xfeed_7025 0 1 decap_w0
xfeed_7024 0 1 tie
xfeed_7023 0 1 decap_w0
xfeed_7022 0 1 decap_w0
xfeed_7021 0 1 decap_w0
xfeed_7020 0 1 decap_w0
xfeed_5883 0 1 tie
xfeed_5882 0 1 decap_w0
xfeed_5881 0 1 decap_w0
xfeed_5880 0 1 decap_w0
xfeed_1579 0 1 decap_w0
xfeed_1578 0 1 decap_w0
xfeed_1577 0 1 decap_w0
xfeed_1576 0 1 decap_w0
xfeed_1575 0 1 decap_w0
xfeed_1574 0 1 decap_w0
xfeed_1573 0 1 decap_w0
xfeed_1572 0 1 decap_w0
xfeed_1571 0 1 decap_w0
xfeed_1570 0 1 decap_w0
xsubckt_1865_dff_x1 0 1 1937 1874 64 dff_x1
xsubckt_1867_dff_x1 0 1 1936 1872 67 dff_x1
xsubckt_1869_dff_x1 0 1 1935 1870 67 dff_x1
xspare_feed_110 0 1 tie
xspare_feed_111 0 1 decap_w0
xspare_feed_112 0 1 tie
xspare_feed_113 0 1 tie
xdiode_49 0 1 595 diode_w1
xdiode_48 0 1 595 diode_w1
xdiode_47 0 1 595 diode_w1
xdiode_46 0 1 595 diode_w1
xdiode_45 0 1 595 diode_w1
xdiode_44 0 1 595 diode_w1
xdiode_43 0 1 1576 diode_w1
xdiode_42 0 1 1576 diode_w1
xdiode_41 0 1 1575 diode_w1
xdiode_40 0 1 1575 diode_w1
xfeed_13239 0 1 decap_w0
xfeed_13238 0 1 decap_w0
xfeed_13237 0 1 decap_w0
xfeed_13236 0 1 decap_w0
xfeed_13235 0 1 decap_w0
xfeed_13234 0 1 decap_w0
xfeed_13233 0 1 decap_w0
xfeed_13232 0 1 decap_w0
xfeed_13231 0 1 decap_w0
xfeed_13230 0 1 decap_w0
xfeed_12709 0 1 decap_w0
xfeed_12708 0 1 decap_w0
xfeed_12707 0 1 tie
xfeed_12706 0 1 decap_w0
xfeed_12705 0 1 decap_w0
xfeed_12704 0 1 decap_w0
xfeed_12703 0 1 decap_w0
xfeed_12702 0 1 tie
xfeed_12701 0 1 decap_w0
xfeed_12700 0 1 decap_w0
xfeed_5889 0 1 tie
xfeed_5888 0 1 decap_w0
xfeed_5887 0 1 decap_w0
xfeed_5886 0 1 decap_w0
xfeed_5885 0 1 decap_w0
xfeed_5884 0 1 decap_w0
xsubckt_1231_mux2_x1 0 1 1830 2106 2065 1334 mux2_x1
xsubckt_907_mux2_x1 0 1 1581 1582 1996 445 mux2_x1
xsubckt_336_and2_x1 0 1 412 415 413 and2_x1
xsubckt_382_nand3_x0 0 1 367 652 535 369 nand3_x0
xsubckt_1591_and21nor_x0 0 1 1003 1070 1015 1073 and21nor_x0
xfeed_7039 0 1 decap_w0
xfeed_7038 0 1 tie
xfeed_7037 0 1 decap_w0
xfeed_7036 0 1 decap_w0
xfeed_7035 0 1 decap_w0
xfeed_7034 0 1 decap_w0
xfeed_7033 0 1 decap_w0
xfeed_7032 0 1 decap_w0
xfeed_7031 0 1 tie
xfeed_7030 0 1 decap_w0
xfeed_6509 0 1 decap_w0
xfeed_6508 0 1 decap_w0
xfeed_6507 0 1 decap_w0
xfeed_6506 0 1 decap_w0
xfeed_6505 0 1 decap_w0
xfeed_6504 0 1 decap_w0
xfeed_6503 0 1 decap_w0
xfeed_6502 0 1 decap_w0
xfeed_6501 0 1 decap_w0
xfeed_6500 0 1 decap_w0
xfeed_5890 0 1 decap_w0
xfeed_1589 0 1 decap_w0
xfeed_1588 0 1 decap_w0
xfeed_1587 0 1 decap_w0
xfeed_1586 0 1 decap_w0
xfeed_1585 0 1 tie
xfeed_1584 0 1 decap_w0
xfeed_1583 0 1 decap_w0
xfeed_1582 0 1 decap_w0
xfeed_1581 0 1 decap_w0
xfeed_1580 0 1 decap_w0
xsubckt_893_mux2_x1 0 1 1593 1594 1998 445 mux2_x1
xsubckt_244_and2_x1 0 1 507 509 508 and2_x1
xsubckt_218_and3_x1 0 1 536 610 595 558 and3_x1
xsubckt_182_and4_x1 0 1 576 716 1924 681 599 and4_x1
xsubckt_1474_and4_x1 0 1 1122 1768 1360 1124 1123 and4_x1
xdiode_59 0 1 1996 diode_w1
xdiode_58 0 1 1996 diode_w1
xdiode_57 0 1 1996 diode_w1
xdiode_56 0 1 1996 diode_w1
xdiode_55 0 1 1996 diode_w1
xdiode_54 0 1 1996 diode_w1
xdiode_53 0 1 670 diode_w1
xdiode_52 0 1 670 diode_w1
xdiode_51 0 1 670 diode_w1
xdiode_50 0 1 670 diode_w1
xfeed_13249 0 1 tie
xfeed_13248 0 1 decap_w0
xfeed_13247 0 1 decap_w0
xfeed_13246 0 1 decap_w0
xfeed_13245 0 1 decap_w0
xfeed_13244 0 1 decap_w0
xfeed_13243 0 1 decap_w0
xfeed_13242 0 1 decap_w0
xfeed_13241 0 1 decap_w0
xfeed_13240 0 1 decap_w0
xfeed_12717 0 1 decap_w0
xfeed_12716 0 1 decap_w0
xfeed_12715 0 1 decap_w0
xfeed_12714 0 1 decap_w0
xfeed_12713 0 1 decap_w0
xfeed_12712 0 1 decap_w0
xfeed_12711 0 1 decap_w0
xfeed_12710 0 1 decap_w0
xfeed_5899 0 1 decap_w0
xfeed_5898 0 1 decap_w0
xfeed_5897 0 1 decap_w0
xfeed_5896 0 1 tie
xfeed_5895 0 1 decap_w0
xfeed_5894 0 1 decap_w0
xfeed_5893 0 1 decap_w0
xfeed_5892 0 1 decap_w0
xfeed_5891 0 1 decap_w0
xsubckt_1691_and21nor_x0 0 1 903 904 1117 2052 and21nor_x0
xfeed_12719 0 1 decap_w0
xfeed_12718 0 1 decap_w0
xfeed_7049 0 1 decap_w0
xfeed_7048 0 1 decap_w0
xfeed_7047 0 1 decap_w0
xfeed_7046 0 1 decap_w0
xfeed_7045 0 1 tie
xfeed_7044 0 1 decap_w0
xfeed_7043 0 1 decap_w0
xfeed_7042 0 1 decap_w0
xfeed_7041 0 1 decap_w0
xfeed_7040 0 1 decap_w0
xfeed_6519 0 1 tie
xfeed_6518 0 1 decap_w0
xfeed_6517 0 1 decap_w0
xfeed_6516 0 1 decap_w0
xfeed_6515 0 1 decap_w0
xfeed_6514 0 1 decap_w0
xfeed_6513 0 1 decap_w0
xfeed_6512 0 1 decap_w0
xfeed_6511 0 1 decap_w0
xfeed_6510 0 1 decap_w0
xfeed_2209 0 1 decap_w0
xfeed_2208 0 1 decap_w0
xfeed_2207 0 1 tie
xfeed_2206 0 1 decap_w0
xfeed_2205 0 1 decap_w0
xfeed_2204 0 1 decap_w0
xfeed_2203 0 1 decap_w0
xfeed_2202 0 1 decap_w0
xfeed_2201 0 1 decap_w0
xfeed_2200 0 1 decap_w0
xfeed_1597 0 1 decap_w0
xfeed_1596 0 1 decap_w0
xfeed_1595 0 1 decap_w0
xfeed_1594 0 1 decap_w0
xfeed_1593 0 1 decap_w0
xfeed_1592 0 1 tie
xfeed_1591 0 1 decap_w0
xfeed_1590 0 1 decap_w0
xsubckt_970_and4_x1 0 1 1555 660 624 523 522 and4_x1
xsubckt_965_or21nand_x0 0 1 1871 1560 1559 1573 or21nand_x0
xsubckt_152_and2_x1 0 1 613 716 1924 and2_x1
xsubckt_535_and4_x1 0 1 218 277 276 258 257 and4_x1
xsubckt_1496_and3_x1 0 1 1100 1969 682 595 and3_x1
xdiode_69 0 1 1998 diode_w1
xdiode_68 0 1 1998 diode_w1
xdiode_67 0 1 1998 diode_w1
xdiode_66 0 1 1998 diode_w1
xdiode_65 0 1 1998 diode_w1
xdiode_64 0 1 1997 diode_w1
xdiode_63 0 1 1997 diode_w1
xdiode_62 0 1 1997 diode_w1
xdiode_61 0 1 1997 diode_w1
xdiode_60 0 1 1997 diode_w1
xfeed_13259 0 1 decap_w0
xfeed_13258 0 1 decap_w0
xfeed_13257 0 1 decap_w0
xfeed_13256 0 1 decap_w0
xfeed_13255 0 1 decap_w0
xfeed_13254 0 1 decap_w0
xfeed_13253 0 1 decap_w0
xfeed_13252 0 1 decap_w0
xfeed_13251 0 1 decap_w0
xfeed_13250 0 1 decap_w0
xfeed_12724 0 1 decap_w0
xfeed_12723 0 1 decap_w0
xfeed_12722 0 1 decap_w0
xfeed_12721 0 1 decap_w0
xfeed_12720 0 1 decap_w0
xfeed_1599 0 1 tie
xfeed_1598 0 1 decap_w0
xsubckt_1055_nand3_x0 0 1 1486 629 334 1487 nand3_x0
xfeed_12729 0 1 decap_w0
xfeed_12728 0 1 decap_w0
xfeed_12727 0 1 decap_w0
xfeed_12726 0 1 decap_w0
xfeed_12725 0 1 decap_w0
xfeed_7059 0 1 decap_w0
xfeed_7058 0 1 decap_w0
xfeed_7057 0 1 decap_w0
xfeed_7056 0 1 decap_w0
xfeed_7055 0 1 decap_w0
xfeed_7054 0 1 tie
xfeed_7053 0 1 decap_w0
xfeed_7052 0 1 decap_w0
xfeed_7051 0 1 decap_w0
xfeed_7050 0 1 tie
xfeed_6529 0 1 decap_w0
xfeed_6528 0 1 decap_w0
xfeed_6527 0 1 decap_w0
xfeed_6526 0 1 decap_w0
xfeed_6525 0 1 decap_w0
xfeed_6524 0 1 decap_w0
xfeed_6523 0 1 tie
xfeed_6522 0 1 decap_w0
xfeed_6521 0 1 decap_w0
xfeed_6520 0 1 decap_w0
xfeed_2219 0 1 decap_w0
xfeed_2218 0 1 decap_w0
xfeed_2217 0 1 decap_w0
xfeed_2216 0 1 decap_w0
xfeed_2215 0 1 decap_w0
xfeed_2214 0 1 tie
xfeed_2213 0 1 decap_w0
xfeed_2212 0 1 decap_w0
xfeed_2211 0 1 decap_w0
xfeed_2210 0 1 decap_w0
xsubckt_1378_and4_x1 0 1 1212 435 1663 1214 1213 and4_x1
xsubckt_1408_nand2_x0 0 1 1184 1191 1186 nand2_x0
xsubckt_1586_nand2_x0 0 1 1008 1101 1010 nand2_x0
xdiode_79 0 1 2002 diode_w1
xdiode_78 0 1 2002 diode_w1
xdiode_77 0 1 2001 diode_w1
xdiode_76 0 1 2001 diode_w1
xdiode_75 0 1 2000 diode_w1
xdiode_74 0 1 2000 diode_w1
xdiode_73 0 1 2000 diode_w1
xdiode_72 0 1 1999 diode_w1
xdiode_71 0 1 1999 diode_w1
xdiode_70 0 1 1999 diode_w1
xfeed_13269 0 1 decap_w0
xfeed_13268 0 1 decap_w0
xfeed_13267 0 1 decap_w0
xfeed_13266 0 1 decap_w0
xfeed_13265 0 1 decap_w0
xfeed_13264 0 1 decap_w0
xfeed_13263 0 1 decap_w0
xfeed_13262 0 1 decap_w0
xfeed_13261 0 1 decap_w0
xfeed_13260 0 1 decap_w0
xfeed_12731 0 1 decap_w0
xfeed_12730 0 1 decap_w0
xsubckt_1228_nand2_x0 0 1 1336 1346 1337 nand2_x0
xsubckt_505_and2_x1 0 1 246 248 247 and2_x1
xsubckt_1333_or21nand_x0 0 1 1808 1262 1256 1254 or21nand_x0
xsubckt_1352_and2_x1 0 1 1236 1240 1237 and2_x1
xfeed_12739 0 1 tie
xfeed_12738 0 1 decap_w0
xfeed_12737 0 1 decap_w0
xfeed_12736 0 1 decap_w0
xfeed_12735 0 1 tie
xfeed_12734 0 1 decap_w0
xfeed_12733 0 1 decap_w0
xfeed_12732 0 1 decap_w0
xfeed_7068 0 1 decap_w0
xfeed_7066 0 1 decap_w0
xfeed_7065 0 1 decap_w0
xfeed_7064 0 1 decap_w0
xfeed_7063 0 1 decap_w0
xfeed_7062 0 1 decap_w0
xfeed_7061 0 1 decap_w0
xfeed_7060 0 1 decap_w0
xfeed_6539 0 1 decap_w0
xfeed_6538 0 1 decap_w0
xfeed_6537 0 1 tie
xfeed_6536 0 1 decap_w0
xfeed_6535 0 1 decap_w0
xfeed_6534 0 1 decap_w0
xfeed_6533 0 1 decap_w0
xfeed_6532 0 1 decap_w0
xfeed_6531 0 1 decap_w0
xfeed_6530 0 1 tie
xfeed_2229 0 1 decap_w0
xfeed_2228 0 1 decap_w0
xfeed_2227 0 1 decap_w0
xfeed_2226 0 1 decap_w0
xfeed_2225 0 1 decap_w0
xfeed_2224 0 1 decap_w0
xfeed_2223 0 1 decap_w0
xfeed_2222 0 1 decap_w0
xfeed_2221 0 1 decap_w0
xfeed_2220 0 1 decap_w0
xsubckt_1260_and2_x1 0 1 1320 663 478 and2_x1
xsubckt_936_and2_x1 0 1 1577 1919 725 and2_x1
xsubckt_874_and4_x1 0 1 1609 1962 1964 2054 2051 and4_x1
xsubckt_439_and4_x1 0 1 311 650 644 637 633 and4_x1
xsubckt_579_and2_x1 0 1 176 181 178 and2_x1
xsubckt_1433_or21nand_x0 0 1 1161 1162 1323 690 or21nand_x0
xdiode_89 0 1 666 diode_w1
xdiode_88 0 1 666 diode_w1
xdiode_87 0 1 674 diode_w1
xdiode_86 0 1 674 diode_w1
xdiode_85 0 1 674 diode_w1
xdiode_84 0 1 674 diode_w1
xdiode_83 0 1 674 diode_w1
xdiode_82 0 1 2003 diode_w1
xdiode_81 0 1 2003 diode_w1
xdiode_80 0 1 2003 diode_w1
xfeed_13277 0 1 decap_w0
xfeed_13276 0 1 decap_w0
xfeed_13275 0 1 decap_w0
xfeed_13274 0 1 decap_w0
xfeed_13273 0 1 decap_w0
xfeed_13272 0 1 decap_w0
xfeed_13271 0 1 decap_w0
xfeed_13270 0 1 decap_w0
xsubckt_1034_nand4_x0 0 1 1501 645 637 633 622 nand4_x0
xsubckt_363_or21nand_x0 0 1 386 661 654 624 or21nand_x0
xsubckt_487_and2_x1 0 1 263 265 264 and2_x1
xsubckt_1655_nand3_x0 0 1 939 948 944 942 nand3_x0
xfeed_200 0 1 decap_w0
xfeed_201 0 1 decap_w0
xfeed_202 0 1 decap_w0
xfeed_203 0 1 decap_w0
xfeed_204 0 1 decap_w0
xfeed_205 0 1 decap_w0
xfeed_206 0 1 decap_w0
xfeed_207 0 1 decap_w0
xfeed_208 0 1 decap_w0
xfeed_209 0 1 decap_w0
xfeed_13279 0 1 decap_w0
xfeed_13278 0 1 decap_w0
xfeed_12749 0 1 decap_w0
xfeed_12748 0 1 decap_w0
xfeed_12747 0 1 decap_w0
xfeed_12746 0 1 tie
xfeed_12745 0 1 decap_w0
xfeed_12744 0 1 decap_w0
xfeed_12743 0 1 decap_w0
xfeed_12742 0 1 decap_w0
xfeed_12741 0 1 decap_w0
xfeed_12740 0 1 decap_w0
xfeed_7079 0 1 decap_w0
xfeed_7078 0 1 decap_w0
xfeed_7077 0 1 decap_w0
xfeed_7076 0 1 decap_w0
xfeed_7075 0 1 decap_w0
xfeed_7074 0 1 decap_w0
xfeed_7072 0 1 decap_w0
xfeed_7071 0 1 decap_w0
xfeed_7070 0 1 decap_w0
xfeed_6549 0 1 decap_w0
xfeed_6548 0 1 decap_w0
xfeed_6547 0 1 decap_w0
xfeed_6546 0 1 decap_w0
xfeed_6545 0 1 decap_w0
xfeed_6544 0 1 decap_w0
xfeed_6543 0 1 decap_w0
xfeed_6542 0 1 decap_w0
xfeed_6541 0 1 decap_w0
xfeed_6540 0 1 decap_w0
xfeed_2239 0 1 decap_w0
xfeed_2238 0 1 decap_w0
xfeed_2237 0 1 decap_w0
xfeed_2236 0 1 decap_w0
xfeed_2235 0 1 decap_w0
xfeed_2234 0 1 decap_w0
xfeed_2233 0 1 decap_w0
xfeed_2232 0 1 decap_w0
xfeed_2231 0 1 decap_w0
xfeed_2230 0 1 decap_w0
xfeed_1709 0 1 decap_w0
xfeed_1708 0 1 decap_w0
xfeed_1707 0 1 decap_w0
xfeed_1706 0 1 decap_w0
xfeed_1705 0 1 decap_w0
xfeed_1704 0 1 decap_w0
xfeed_1703 0 1 decap_w0
xfeed_1702 0 1 decap_w0
xfeed_1701 0 1 decap_w0
xfeed_1700 0 1 decap_w0
xsubckt_818_and3_x1 0 1 1657 2070 680 489 and3_x1
xsubckt_409_and2_x1 0 1 340 342 341 and2_x1
xsubckt_1787_and21nor_x0 0 1 807 1029 811 809 and21nor_x0
xdiode_99 0 1 2049 diode_w1
xdiode_98 0 1 2049 diode_w1
xdiode_97 0 1 2049 diode_w1
xdiode_96 0 1 2048 diode_w1
xdiode_95 0 1 2048 diode_w1
xdiode_94 0 1 2048 diode_w1
xdiode_93 0 1 2048 diode_w1
xdiode_92 0 1 666 diode_w1
xdiode_91 0 1 666 diode_w1
xdiode_90 0 1 666 diode_w1
xfeed_13284 0 1 decap_w0
xfeed_13283 0 1 decap_w0
xfeed_13282 0 1 decap_w0
xfeed_13281 0 1 decap_w0
xfeed_13280 0 1 decap_w0
xsubckt_1031_nand2_x0 0 1 1860 1508 1504 nand2_x0
xsubckt_814_or2_x1 0 1 2104 1667 1661 or2_x1
xsubckt_255_and4_x1 0 1 496 504 502 500 497 and4_x1
xsubckt_369_and3_x1 0 1 380 532 530 382 and3_x1
xsubckt_1295_nand3_x0 0 1 1288 2062 666 657 nand3_x0
xfeed_210 0 1 decap_w0
xfeed_211 0 1 decap_w0
xfeed_212 0 1 decap_w0
xfeed_213 0 1 decap_w0
xfeed_214 0 1 decap_w0
xfeed_215 0 1 decap_w0
xfeed_216 0 1 decap_w0
xfeed_217 0 1 decap_w0
xfeed_218 0 1 decap_w0
xfeed_219 0 1 decap_w0
xfeed_13289 0 1 decap_w0
xfeed_13288 0 1 decap_w0
xfeed_13287 0 1 decap_w0
xfeed_13286 0 1 decap_w0
xfeed_13285 0 1 decap_w0
xfeed_12759 0 1 decap_w0
xfeed_12758 0 1 decap_w0
xfeed_12757 0 1 decap_w0
xfeed_12756 0 1 decap_w0
xfeed_12755 0 1 decap_w0
xfeed_12754 0 1 decap_w0
xfeed_12753 0 1 decap_w0
xfeed_12752 0 1 decap_w0
xfeed_12751 0 1 tie
xfeed_12750 0 1 decap_w0
xfeed_7089 0 1 tie
xfeed_7088 0 1 decap_w0
xfeed_7087 0 1 decap_w0
xfeed_7086 0 1 decap_w0
xfeed_7085 0 1 decap_w0
xfeed_7084 0 1 decap_w0
xfeed_7083 0 1 decap_w0
xfeed_7082 0 1 tie
xfeed_7081 0 1 decap_w0
xfeed_7080 0 1 decap_w0
xfeed_6559 0 1 tie
xfeed_6558 0 1 decap_w0
xfeed_6557 0 1 decap_w0
xfeed_6556 0 1 decap_w0
xfeed_6555 0 1 decap_w0
xfeed_6554 0 1 decap_w0
xfeed_6553 0 1 decap_w0
xfeed_6552 0 1 decap_w0
xfeed_6551 0 1 decap_w0
xfeed_6550 0 1 decap_w0
xfeed_2249 0 1 decap_w0
xfeed_2248 0 1 decap_w0
xfeed_2247 0 1 decap_w0
xfeed_2246 0 1 decap_w0
xfeed_2245 0 1 decap_w0
xfeed_2244 0 1 decap_w0
xfeed_2243 0 1 decap_w0
xfeed_2242 0 1 decap_w0
xfeed_2241 0 1 decap_w0
xfeed_2240 0 1 decap_w0
xfeed_1719 0 1 decap_w0
xfeed_1718 0 1 decap_w0
xfeed_1717 0 1 decap_w0
xfeed_1716 0 1 decap_w0
xfeed_1715 0 1 decap_w0
xfeed_1714 0 1 decap_w0
xfeed_1713 0 1 decap_w0
xfeed_1712 0 1 decap_w0
xfeed_1711 0 1 decap_w0
xfeed_1710 0 1 decap_w0
xsubckt_1164_and2_x1 0 1 1397 1399 1398 and2_x1
xsubckt_1024_and4_x1 0 1 1510 1916 1927 679 674 and4_x1
xsubckt_954_nand3_x0 0 1 1566 660 654 527 nand3_x0
xsubckt_772_or2_x1 0 1 2095 1699 1698 or2_x1
xsubckt_770_or2_x1 0 1 1699 1704 1703 or2_x1
xsubckt_726_and3_x1 0 1 1738 1982 1749 1739 and3_x1
xfeed_13291 0 1 decap_w0
xfeed_13290 0 1 decap_w0
xsubckt_778_or2_x1 0 1 1692 1697 1696 or2_x1
xsubckt_243_nand4_x0 0 1 508 652 649 645 535 nand4_x0
xsubckt_383_or2_x1 0 1 366 554 501 or2_x1
xsubckt_1319_or2_x1 0 1 1266 1270 1267 or2_x1
xsubckt_1660_or2_x1 0 1 934 694 1116 or2_x1
xsubckt_1790_and21nor_x0 0 1 804 1060 806 805 and21nor_x0
xfeed_220 0 1 decap_w0
xfeed_221 0 1 decap_w0
xfeed_223 0 1 decap_w0
xfeed_224 0 1 decap_w0
xfeed_225 0 1 decap_w0
xfeed_226 0 1 decap_w0
xfeed_227 0 1 tie
xfeed_228 0 1 decap_w0
xfeed_229 0 1 decap_w0
xfeed_13299 0 1 decap_w0
xfeed_13298 0 1 decap_w0
xfeed_13297 0 1 decap_w0
xfeed_13296 0 1 decap_w0
xfeed_13295 0 1 decap_w0
xfeed_13294 0 1 tie
xfeed_13293 0 1 decap_w0
xfeed_13292 0 1 decap_w0
xfeed_12769 0 1 decap_w0
xfeed_12768 0 1 decap_w0
xfeed_12767 0 1 decap_w0
xfeed_12766 0 1 decap_w0
xfeed_12765 0 1 decap_w0
xfeed_12764 0 1 decap_w0
xfeed_12763 0 1 decap_w0
xfeed_12762 0 1 decap_w0
xfeed_12761 0 1 decap_w0
xfeed_12760 0 1 decap_w0
xfeed_7099 0 1 decap_w0
xfeed_7098 0 1 decap_w0
xfeed_7097 0 1 decap_w0
xfeed_7096 0 1 decap_w0
xfeed_7095 0 1 decap_w0
xfeed_7094 0 1 decap_w0
xfeed_7093 0 1 decap_w0
xfeed_7092 0 1 decap_w0
xfeed_7091 0 1 decap_w0
xfeed_7090 0 1 decap_w0
xfeed_6569 0 1 decap_w0
xfeed_6568 0 1 decap_w0
xfeed_6567 0 1 decap_w0
xfeed_6566 0 1 tie
xfeed_6565 0 1 decap_w0
xfeed_6564 0 1 decap_w0
xfeed_6563 0 1 decap_w0
xfeed_6562 0 1 decap_w0
xfeed_6561 0 1 decap_w0
xfeed_6560 0 1 decap_w0
xfeed_2259 0 1 decap_w0
xfeed_2258 0 1 decap_w0
xfeed_2257 0 1 decap_w0
xfeed_2256 0 1 decap_w0
xfeed_2255 0 1 decap_w0
xfeed_2254 0 1 decap_w0
xfeed_2253 0 1 decap_w0
xfeed_2252 0 1 decap_w0
xfeed_2251 0 1 decap_w0
xfeed_2250 0 1 tie
xfeed_1729 0 1 decap_w0
xfeed_1728 0 1 decap_w0
xfeed_1727 0 1 decap_w0
xfeed_1726 0 1 tie
xfeed_1725 0 1 decap_w0
xfeed_1724 0 1 decap_w0
xfeed_1723 0 1 decap_w0
xfeed_1722 0 1 decap_w0
xfeed_1721 0 1 decap_w0
xfeed_1720 0 1 decap_w0
xsubckt_225_and2_x1 0 1 526 661 527 and2_x1
xsubckt_506_nand3_x0 0 1 245 679 557 405 nand3_x0
xsubckt_520_and4_x1 0 1 232 378 355 349 259 and4_x1
xsubckt_1185_and21nor_x0 0 1 1379 666 617 581 and21nor_x0
xsubckt_416_nand3_x0 0 1 333 653 535 369 nand3_x0
xfeed_230 0 1 decap_w0
xfeed_231 0 1 decap_w0
xfeed_232 0 1 decap_w0
xfeed_233 0 1 decap_w0
xfeed_234 0 1 decap_w0
xfeed_235 0 1 decap_w0
xfeed_236 0 1 decap_w0
xfeed_237 0 1 decap_w0
xfeed_238 0 1 decap_w0
xfeed_239 0 1 tie
xfeed_12779 0 1 decap_w0
xfeed_12778 0 1 decap_w0
xfeed_12777 0 1 decap_w0
xfeed_12776 0 1 decap_w0
xfeed_12775 0 1 decap_w0
xfeed_12774 0 1 decap_w0
xfeed_12773 0 1 decap_w0
xfeed_12772 0 1 decap_w0
xfeed_12771 0 1 decap_w0
xfeed_12770 0 1 decap_w0
xfeed_6576 0 1 decap_w0
xfeed_6575 0 1 decap_w0
xfeed_6574 0 1 decap_w0
xfeed_6573 0 1 decap_w0
xfeed_6572 0 1 decap_w0
xfeed_6571 0 1 decap_w0
xfeed_6570 0 1 decap_w0
xfeed_2269 0 1 decap_w0
xfeed_2268 0 1 decap_w0
xfeed_2267 0 1 decap_w0
xfeed_2266 0 1 decap_w0
xfeed_2265 0 1 tie
xfeed_2264 0 1 decap_w0
xfeed_2263 0 1 decap_w0
xfeed_2262 0 1 decap_w0
xfeed_2261 0 1 decap_w0
xfeed_2260 0 1 decap_w0
xfeed_1737 0 1 decap_w0
xfeed_1736 0 1 tie
xfeed_1735 0 1 decap_w0
xfeed_1734 0 1 decap_w0
xfeed_1733 0 1 decap_w0
xfeed_1732 0 1 decap_w0
xfeed_1731 0 1 decap_w0
xfeed_1730 0 1 decap_w0
xsubckt_1116_mux2_x1 0 1 1841 1999 1990 1438 mux2_x1
xsubckt_516_and4_x1 0 1 235 373 361 255 236 and4_x1
xfeed_6579 0 1 decap_w0
xfeed_6578 0 1 decap_w0
xfeed_6577 0 1 decap_w0
xfeed_1739 0 1 decap_w0
xfeed_1738 0 1 decap_w0
xsubckt_1271_nand2_x0 0 1 1814 1333 1310 nand2_x0
xfeed_0 0 1 decap_w0
xfeed_240 0 1 decap_w0
xfeed_241 0 1 decap_w0
xfeed_242 0 1 decap_w0
xfeed_243 0 1 decap_w0
xfeed_244 0 1 decap_w0
xfeed_245 0 1 decap_w0
xfeed_246 0 1 tie
xfeed_247 0 1 decap_w0
xfeed_248 0 1 decap_w0
xfeed_249 0 1 decap_w0
xfeed_12789 0 1 decap_w0
xfeed_12788 0 1 decap_w0
xfeed_12787 0 1 decap_w0
xfeed_12786 0 1 decap_w0
xfeed_12785 0 1 decap_w0
xfeed_12784 0 1 decap_w0
xfeed_12783 0 1 decap_w0
xfeed_12782 0 1 decap_w0
xfeed_12781 0 1 decap_w0
xfeed_12780 0 1 decap_w0
xfeed_6583 0 1 decap_w0
xfeed_6582 0 1 decap_w0
xfeed_6581 0 1 decap_w0
xfeed_6580 0 1 decap_w0
xfeed_2279 0 1 decap_w0
xfeed_2278 0 1 decap_w0
xfeed_2277 0 1 decap_w0
xfeed_2276 0 1 decap_w0
xfeed_2275 0 1 decap_w0
xfeed_2274 0 1 decap_w0
xfeed_2273 0 1 decap_w0
xfeed_2272 0 1 decap_w0
xfeed_2271 0 1 decap_w0
xfeed_2270 0 1 decap_w0
xfeed_1744 0 1 decap_w0
xfeed_1743 0 1 decap_w0
xfeed_1742 0 1 decap_w0
xfeed_1741 0 1 decap_w0
xfeed_1740 0 1 decap_w0
xsubckt_1629_or21nand_x0 0 1 965 968 1118 764 or21nand_x0
xfeed_1 0 1 decap_w0
xfeed_2 0 1 decap_w0
xfeed_3 0 1 decap_w0
xfeed_4 0 1 decap_w0
xfeed_5 0 1 decap_w0
xfeed_6 0 1 decap_w0
xfeed_7 0 1 tie
xfeed_8 0 1 decap_w0
xfeed_9 0 1 decap_w0
xfeed_13409 0 1 decap_w0
xfeed_13408 0 1 decap_w0
xfeed_13407 0 1 decap_w0
xfeed_13406 0 1 decap_w0
xfeed_13405 0 1 decap_w0
xfeed_13404 0 1 decap_w0
xfeed_13403 0 1 decap_w0
xfeed_13402 0 1 decap_w0
xfeed_13401 0 1 tie
xfeed_13400 0 1 decap_w0
xfeed_6589 0 1 tie
xfeed_6588 0 1 decap_w0
xfeed_6587 0 1 decap_w0
xfeed_6586 0 1 decap_w0
xfeed_6585 0 1 decap_w0
xfeed_6584 0 1 decap_w0
xfeed_1749 0 1 decap_w0
xfeed_1748 0 1 decap_w0
xfeed_1747 0 1 decap_w0
xfeed_1746 0 1 decap_w0
xfeed_1745 0 1 decap_w0
xsubckt_1177_nand3_x0 0 1 1385 2013 1393 1386 nand3_x0
xsubckt_1131_or21nand_x0 0 1 1426 1427 1428 1434 or21nand_x0
xsubckt_881_and3_x1 0 1 1603 1962 767 766 and3_x1
xsubckt_323_and21nor_x0 0 1 425 429 427 535 and21nor_x0
xsubckt_472_and2_x1 0 1 278 280 279 and2_x1
xsubckt_1532_or21nand_x0 0 1 1798 1144 1062 774 or21nand_x0
xfeed_250 0 1 decap_w0
xfeed_251 0 1 decap_w0
xfeed_252 0 1 decap_w0
xfeed_253 0 1 decap_w0
xfeed_254 0 1 decap_w0
xfeed_256 0 1 tie
xfeed_257 0 1 decap_w0
xfeed_258 0 1 decap_w0
xfeed_259 0 1 decap_w0
xfeed_12799 0 1 decap_w0
xfeed_12798 0 1 decap_w0
xfeed_12797 0 1 decap_w0
xfeed_12796 0 1 decap_w0
xfeed_12795 0 1 decap_w0
xfeed_12794 0 1 decap_w0
xfeed_12793 0 1 decap_w0
xfeed_12792 0 1 decap_w0
xfeed_12791 0 1 decap_w0
xfeed_12790 0 1 decap_w0
xfeed_7209 0 1 decap_w0
xfeed_7208 0 1 decap_w0
xfeed_7207 0 1 tie
xfeed_7206 0 1 decap_w0
xfeed_7205 0 1 decap_w0
xfeed_7204 0 1 decap_w0
xfeed_7203 0 1 decap_w0
xfeed_7202 0 1 decap_w0
xfeed_7201 0 1 decap_w0
xfeed_7200 0 1 decap_w0
xfeed_6590 0 1 decap_w0
xfeed_2289 0 1 decap_w0
xfeed_2288 0 1 decap_w0
xfeed_2287 0 1 decap_w0
xfeed_2286 0 1 decap_w0
xfeed_2285 0 1 decap_w0
xfeed_2284 0 1 decap_w0
xfeed_2283 0 1 decap_w0
xfeed_2282 0 1 decap_w0
xfeed_2281 0 1 decap_w0
xfeed_2280 0 1 decap_w0
xfeed_1751 0 1 decap_w0
xfeed_1750 0 1 decap_w0
xsubckt_824_and21nor_x0 0 1 1652 692 1755 1754 and21nor_x0
xsubckt_229_nand2_x0 0 1 522 785 1997 nand2_x0
xsubckt_393_nand4_x0 0 1 356 533 524 518 360 nand4_x0
xsubckt_1328_or21nand_x0 0 1 1258 1259 1322 760 or21nand_x0
xsubckt_1738_and3_x1 0 1 856 1069 873 871 and3_x1
xsubckt_1910_dff_x1 0 1 1966 1837 61 dff_x1
xsubckt_1912_dff_x1 0 1 2012 1835 61 dff_x1
xsubckt_1914_dff_x1 0 1 1965 1833 61 dff_x1
xfeed_13417 0 1 decap_w0
xfeed_13416 0 1 decap_w0
xfeed_13415 0 1 decap_w0
xfeed_13414 0 1 decap_w0
xfeed_13413 0 1 decap_w0
xfeed_13412 0 1 decap_w0
xfeed_13411 0 1 decap_w0
xfeed_13410 0 1 decap_w0
xfeed_6599 0 1 tie
xfeed_6598 0 1 decap_w0
xfeed_6597 0 1 decap_w0
xfeed_6596 0 1 decap_w0
xfeed_6595 0 1 decap_w0
xfeed_6594 0 1 decap_w0
xfeed_6593 0 1 decap_w0
xfeed_6592 0 1 decap_w0
xfeed_6591 0 1 decap_w0
xfeed_1759 0 1 decap_w0
xfeed_1758 0 1 decap_w0
xfeed_1757 0 1 decap_w0
xfeed_1756 0 1 decap_w0
xfeed_1755 0 1 tie
xfeed_1754 0 1 decap_w0
xfeed_1753 0 1 decap_w0
xfeed_1752 0 1 decap_w0
xsubckt_656_nand3_x0 0 1 104 2024 184 176 nand3_x0
xsubckt_1781_nexor2_x0 0 1 813 1004 998 nexor2_x0
xsubckt_1870_dff_x1 0 1 1956 1869 67 dff_x1
xsubckt_1916_dff_x1 0 1 1962 1786 61 dff_x1
xsubckt_1918_dff_x1 0 1 2065 1830 51 dff_x1
xfeed_260 0 1 decap_w0
xfeed_261 0 1 tie
xfeed_262 0 1 decap_w0
xfeed_263 0 1 decap_w0
xfeed_264 0 1 decap_w0
xfeed_265 0 1 decap_w0
xfeed_266 0 1 decap_w0
xfeed_267 0 1 decap_w0
xfeed_268 0 1 decap_w0
xfeed_269 0 1 decap_w0
xfeed_13419 0 1 decap_w0
xfeed_13418 0 1 decap_w0
xfeed_7219 0 1 decap_w0
xfeed_7218 0 1 tie
xfeed_7217 0 1 decap_w0
xfeed_7215 0 1 decap_w0
xfeed_7214 0 1 decap_w0
xfeed_7213 0 1 decap_w0
xfeed_7211 0 1 tie
xfeed_7210 0 1 decap_w0
xfeed_2297 0 1 decap_w0
xfeed_2296 0 1 decap_w0
xfeed_2295 0 1 decap_w0
xfeed_2294 0 1 decap_w0
xfeed_2293 0 1 decap_w0
xfeed_2292 0 1 decap_w0
xfeed_2291 0 1 tie
xfeed_2290 0 1 decap_w0
xsubckt_825_and2_x1 0 1 1651 2049 1740 and2_x1
xsubckt_302_and2_x1 0 1 446 616 447 and2_x1
xsubckt_212_nand2_x0 0 1 542 687 544 nand2_x0
xsubckt_1603_nand2_x0 0 1 991 995 993 nand2_x0
xsubckt_1808_mux2_x1 0 1 1794 2051 827 773 mux2_x1
xsubckt_1872_dff_x1 0 1 1945 1867 77 dff_x1
xsubckt_1874_dff_x1 0 1 1943 1865 77 dff_x1
xsubckt_1876_dff_x1 0 1 1938 1863 77 dff_x1
xfeed_13424 0 1 decap_w0
xfeed_13423 0 1 decap_w0
xfeed_13422 0 1 decap_w0
xfeed_13421 0 1 decap_w0
xfeed_13420 0 1 decap_w0
xfeed_2299 0 1 decap_w0
xfeed_2298 0 1 decap_w0
xfeed_1769 0 1 tie
xfeed_1768 0 1 decap_w0
xfeed_1767 0 1 decap_w0
xfeed_1766 0 1 decap_w0
xfeed_1765 0 1 decap_w0
xfeed_1764 0 1 decap_w0
xfeed_1763 0 1 decap_w0
xfeed_1762 0 1 tie
xfeed_1761 0 1 decap_w0
xfeed_1760 0 1 decap_w0
xsubckt_1123_or2_x1 0 1 1434 1940 1956 or2_x1
xsubckt_671_and4_x1 0 1 90 94 93 92 91 and4_x1
xsubckt_662_or21nand_x0 0 1 98 1971 450 411 or21nand_x0
xsubckt_376_and2_x1 0 1 373 378 374 and2_x1
xsubckt_1513_nand2_x0 0 1 1083 1125 1085 nand2_x0
xsubckt_1585_and21nor_x0 0 1 1009 1102 1012 1011 and21nor_x0
xsubckt_1878_dff_x1 0 1 1955 1861 67 dff_x1
xfeed_270 0 1 decap_w0
xfeed_271 0 1 decap_w0
xfeed_272 0 1 decap_w0
xfeed_273 0 1 decap_w0
xfeed_274 0 1 decap_w0
xfeed_275 0 1 decap_w0
xfeed_276 0 1 decap_w0
xfeed_277 0 1 decap_w0
xfeed_278 0 1 decap_w0
xfeed_279 0 1 decap_w0
xfeed_13429 0 1 decap_w0
xfeed_13428 0 1 decap_w0
xfeed_13427 0 1 decap_w0
xfeed_13426 0 1 tie
xfeed_13425 0 1 decap_w0
xfeed_7229 0 1 decap_w0
xfeed_7228 0 1 decap_w0
xfeed_7227 0 1 decap_w0
xfeed_7226 0 1 decap_w0
xfeed_7225 0 1 tie
xfeed_7224 0 1 decap_w0
xfeed_7222 0 1 decap_w0
xfeed_7221 0 1 decap_w0
xfeed_7220 0 1 decap_w0
xsubckt_1184_and21nor_x0 0 1 1380 544 581 608 and21nor_x0
xsubckt_1502_and2_x1 0 1 1094 1099 1095 and2_x1
xsubckt_1509_nand3_x0 0 1 1087 1119 1112 1092 nand3_x0
xsubckt_1528_or21nand_x0 0 1 1065 1067 1072 1093 or21nand_x0
xfeed_13431 0 1 decap_w0
xfeed_13430 0 1 decap_w0
xfeed_1779 0 1 decap_w0
xfeed_1778 0 1 decap_w0
xfeed_1777 0 1 decap_w0
xfeed_1776 0 1 decap_w0
xfeed_1775 0 1 decap_w0
xfeed_1774 0 1 decap_w0
xfeed_1773 0 1 decap_w0
xfeed_1772 0 1 decap_w0
xfeed_1771 0 1 decap_w0
xfeed_1770 0 1 decap_w0
xsubckt_1203_nor3_x0 0 1 1361 1369 1367 1362 nor3_x0
xsubckt_1153_nand2_x0 0 1 1407 484 1408 nand2_x0
xsubckt_1027_and3_x1 0 1 1507 638 632 1510 and3_x1
xsubckt_170_and3_x1 0 1 588 680 599 589 and3_x1
xfeed_280 0 1 decap_w0
xfeed_281 0 1 decap_w0
xfeed_282 0 1 decap_w0
xfeed_283 0 1 decap_w0
xfeed_284 0 1 decap_w0
xfeed_285 0 1 decap_w0
xfeed_286 0 1 decap_w0
xfeed_287 0 1 decap_w0
xfeed_288 0 1 tie
xfeed_289 0 1 decap_w0
xfeed_13439 0 1 decap_w0
xfeed_13438 0 1 decap_w0
xfeed_13437 0 1 decap_w0
xfeed_13436 0 1 decap_w0
xfeed_13435 0 1 decap_w0
xfeed_13434 0 1 decap_w0
xfeed_13433 0 1 decap_w0
xfeed_13432 0 1 decap_w0
xfeed_12909 0 1 decap_w0
xfeed_12908 0 1 decap_w0
xfeed_12907 0 1 decap_w0
xfeed_12906 0 1 decap_w0
xfeed_12905 0 1 decap_w0
xfeed_12904 0 1 decap_w0
xfeed_12903 0 1 decap_w0
xfeed_12902 0 1 decap_w0
xfeed_12901 0 1 decap_w0
xfeed_12900 0 1 decap_w0
xfeed_7238 0 1 decap_w0
xfeed_7237 0 1 tie
xfeed_7235 0 1 decap_w0
xfeed_7234 0 1 decap_w0
xfeed_7233 0 1 decap_w0
xfeed_7232 0 1 decap_w0
xfeed_7231 0 1 decap_w0
xfeed_7230 0 1 decap_w0
xfeed_6709 0 1 decap_w0
xfeed_6708 0 1 decap_w0
xfeed_6707 0 1 decap_w0
xfeed_6706 0 1 decap_w0
xfeed_6705 0 1 tie
xfeed_6704 0 1 decap_w0
xfeed_6703 0 1 decap_w0
xfeed_6702 0 1 decap_w0
xfeed_6701 0 1 decap_w0
xfeed_6700 0 1 decap_w0
xsubckt_1163_nor4_x0 0 1 1398 2053 2052 2051 2050 nor4_x0
xsubckt_990_nand2_x0 0 1 1538 1944 1575 nand2_x0
xsubckt_469_nand2_x0 0 1 281 345 343 nand2_x0
xfeed_1789 0 1 decap_w0
xfeed_1788 0 1 decap_w0
xfeed_1787 0 1 decap_w0
xfeed_1786 0 1 decap_w0
xfeed_1785 0 1 decap_w0
xfeed_1784 0 1 decap_w0
xfeed_1783 0 1 decap_w0
xfeed_1782 0 1 decap_w0
xfeed_1781 0 1 decap_w0
xfeed_1780 0 1 decap_w0
xsubckt_1175_mux2_x1 0 1 1387 1388 485 1392 mux2_x1
xsubckt_722_nand2_x0 0 1 1742 600 1745 nand2_x0
xsubckt_1458_and3_x1 0 1 1138 779 756 548 and3_x1
xsubckt_1490_nand3_x0 0 1 1106 547 1745 1108 nand3_x0
xsubckt_1531_or21nand_x0 0 1 1062 1063 1065 1074 or21nand_x0
xspare_buffer_11 0 1 16 22 buf_x4
xspare_buffer_12 0 1 55 82 buf_x4
xspare_buffer_15 0 1 11 22 buf_x4
xspare_buffer_16 0 1 42 82 buf_x4
xspare_buffer_19 0 1 6 22 buf_x4
xfeed_290 0 1 decap_w0
xfeed_291 0 1 decap_w0
xfeed_292 0 1 decap_w0
xfeed_293 0 1 decap_w0
xfeed_294 0 1 decap_w0
xfeed_295 0 1 tie
xfeed_296 0 1 decap_w0
xfeed_298 0 1 decap_w0
xfeed_299 0 1 decap_w0
xfeed_13449 0 1 decap_w0
xfeed_13448 0 1 decap_w0
xfeed_13447 0 1 decap_w0
xfeed_13446 0 1 decap_w0
xfeed_13445 0 1 decap_w0
xfeed_13444 0 1 decap_w0
xfeed_13443 0 1 decap_w0
xfeed_13442 0 1 decap_w0
xfeed_13441 0 1 decap_w0
xfeed_13440 0 1 decap_w0
xfeed_12919 0 1 decap_w0
xfeed_12917 0 1 decap_w0
xfeed_12916 0 1 decap_w0
xfeed_12915 0 1 decap_w0
xfeed_12914 0 1 decap_w0
xfeed_12913 0 1 decap_w0
xfeed_12912 0 1 tie
xfeed_12911 0 1 decap_w0
xfeed_12910 0 1 decap_w0
xfeed_7249 0 1 decap_w0
xfeed_7248 0 1 decap_w0
xfeed_7247 0 1 decap_w0
xfeed_7246 0 1 decap_w0
xfeed_7245 0 1 decap_w0
xfeed_7244 0 1 decap_w0
xfeed_7243 0 1 decap_w0
xfeed_7242 0 1 decap_w0
xfeed_7241 0 1 decap_w0
xfeed_7240 0 1 decap_w0
xfeed_6716 0 1 decap_w0
xfeed_6715 0 1 decap_w0
xfeed_6714 0 1 decap_w0
xfeed_6713 0 1 decap_w0
xfeed_6712 0 1 decap_w0
xfeed_6711 0 1 decap_w0
xfeed_6710 0 1 decap_w0
xfeed_2409 0 1 decap_w0
xfeed_2408 0 1 tie
xfeed_2407 0 1 decap_w0
xfeed_2406 0 1 decap_w0
xfeed_2405 0 1 decap_w0
xfeed_2404 0 1 decap_w0
xfeed_2403 0 1 decap_w0
xfeed_2402 0 1 decap_w0
xfeed_2401 0 1 decap_w0
xfeed_2400 0 1 decap_w0
xsubckt_1222_nand3_x0 0 1 1342 1351 1346 1343 nand3_x0
xsubckt_896_nand3_x0 0 1 1591 1962 1964 2055 nand3_x0
xsubckt_597_and3_x1 0 1 158 164 160 159 and3_x1
xsubckt_1406_and2_x1 0 1 1186 1190 1187 and2_x1
xsubckt_1796_nexor2_x0 0 1 798 812 808 nexor2_x0
xfeed_6719 0 1 decap_w0
xfeed_6718 0 1 decap_w0
xfeed_6717 0 1 decap_w0
xfeed_1799 0 1 decap_w0
xfeed_1798 0 1 decap_w0
xfeed_1797 0 1 decap_w0
xfeed_1796 0 1 decap_w0
xfeed_1795 0 1 decap_w0
xfeed_1794 0 1 decap_w0
xfeed_1793 0 1 decap_w0
xfeed_1792 0 1 decap_w0
xfeed_1791 0 1 decap_w0
xfeed_1790 0 1 decap_w0
xsubckt_962_or21nand_x0 0 1 1872 1561 1562 1566 or21nand_x0
xsubckt_1484_and21nor_x0 0 1 1112 1113 1117 2046 and21nor_x0
xsubckt_1631_or21nand_x0 0 1 963 966 1122 129 or21nand_x0
xspare_buffer_20 0 1 80 81 buf_x4
xspare_buffer_21 0 1 79 81 buf_x4
xspare_buffer_22 0 1 78 81 buf_x4
xspare_buffer_23 0 1 20 21 buf_x4
xspare_buffer_24 0 1 77 81 buf_x4
xspare_buffer_25 0 1 76 81 buf_x4
xspare_buffer_26 0 1 75 81 buf_x4
xspare_buffer_27 0 1 19 21 buf_x4
xspare_buffer_28 0 1 74 81 buf_x4
xspare_buffer_29 0 1 73 81 buf_x4
xfeed_13459 0 1 decap_w0
xfeed_13458 0 1 decap_w0
xfeed_13457 0 1 decap_w0
xfeed_13456 0 1 decap_w0
xfeed_13455 0 1 decap_w0
xfeed_13454 0 1 decap_w0
xfeed_13453 0 1 decap_w0
xfeed_13452 0 1 decap_w0
xfeed_13451 0 1 decap_w0
xfeed_13450 0 1 decap_w0
xfeed_12929 0 1 tie
xfeed_12928 0 1 decap_w0
xfeed_12927 0 1 decap_w0
xfeed_12926 0 1 decap_w0
xfeed_12925 0 1 decap_w0
xfeed_12924 0 1 decap_w0
xfeed_12923 0 1 decap_w0
xfeed_12922 0 1 decap_w0
xfeed_12921 0 1 decap_w0
xfeed_12920 0 1 decap_w0
xfeed_7259 0 1 decap_w0
xfeed_7258 0 1 decap_w0
xfeed_7257 0 1 decap_w0
xfeed_7256 0 1 decap_w0
xfeed_7255 0 1 decap_w0
xfeed_7254 0 1 tie
xfeed_7253 0 1 decap_w0
xfeed_7252 0 1 decap_w0
xfeed_7250 0 1 decap_w0
xfeed_6723 0 1 decap_w0
xfeed_6722 0 1 decap_w0
xfeed_6721 0 1 decap_w0
xfeed_6720 0 1 decap_w0
xfeed_2419 0 1 decap_w0
xfeed_2418 0 1 decap_w0
xfeed_2417 0 1 decap_w0
xfeed_2416 0 1 decap_w0
xfeed_2415 0 1 tie
xfeed_2414 0 1 decap_w0
xfeed_2413 0 1 decap_w0
xfeed_2412 0 1 decap_w0
xfeed_2411 0 1 decap_w0
xfeed_2410 0 1 decap_w0
xsubckt_272_nand2_x0 0 1 476 678 490 nand2_x0
xsubckt_144_mux2_x1 0 1 624 1987 1996 1986 mux2_x1
xsubckt_1427_or21nand_x0 0 1 1801 1179 1170 1167 or21nand_x0
xcmpt_abc_11867_new_n583_hfns_0 0 1 490 488 buf_x4
xcmpt_abc_11867_new_n583_hfns_1 0 1 489 488 buf_x4
xfeed_6729 0 1 decap_w0
xfeed_6728 0 1 decap_w0
xfeed_6727 0 1 decap_w0
xfeed_6726 0 1 decap_w0
xfeed_6725 0 1 decap_w0
xfeed_6724 0 1 decap_w0
xsubckt_719_and21nor_x0 0 1 1745 468 581 608 and21nor_x0
xsubckt_427_and3_x1 0 1 322 330 329 327 and3_x1
xspare_buffer_30 0 1 72 81 buf_x4
xspare_buffer_31 0 1 18 21 buf_x4
xspare_buffer_32 0 1 71 81 buf_x4
xspare_buffer_33 0 1 70 81 buf_x4
xspare_buffer_34 0 1 69 81 buf_x4
xspare_buffer_35 0 1 17 21 buf_x4
xspare_buffer_36 0 1 67 68 buf_x4
xspare_buffer_37 0 1 66 68 buf_x4
xcmpt_abc_11867_new_n583_hfns_2 0 1 488 491 buf_x4
xfeed_13469 0 1 decap_w0
xfeed_13468 0 1 decap_w0
xfeed_13467 0 1 decap_w0
xfeed_13466 0 1 decap_w0
xfeed_13465 0 1 decap_w0
xfeed_13464 0 1 decap_w0
xfeed_13463 0 1 decap_w0
xfeed_13462 0 1 decap_w0
xfeed_13461 0 1 decap_w0
xfeed_13460 0 1 decap_w0
xfeed_12939 0 1 decap_w0
xfeed_12938 0 1 decap_w0
xfeed_12937 0 1 decap_w0
xfeed_12936 0 1 decap_w0
xfeed_12935 0 1 decap_w0
xfeed_12934 0 1 decap_w0
xfeed_12933 0 1 decap_w0
xfeed_12932 0 1 decap_w0
xfeed_12930 0 1 decap_w0
xfeed_7269 0 1 decap_w0
xfeed_7268 0 1 decap_w0
xfeed_7267 0 1 decap_w0
xfeed_7266 0 1 tie
xfeed_7265 0 1 decap_w0
xfeed_7264 0 1 decap_w0
xfeed_7263 0 1 decap_w0
xfeed_7262 0 1 decap_w0
xfeed_7261 0 1 decap_w0
xfeed_7260 0 1 decap_w0
xfeed_6730 0 1 decap_w0
xfeed_2429 0 1 decap_w0
xfeed_2428 0 1 decap_w0
xfeed_2427 0 1 decap_w0
xfeed_2426 0 1 decap_w0
xfeed_2425 0 1 decap_w0
xfeed_2424 0 1 decap_w0
xfeed_2423 0 1 decap_w0
xfeed_2422 0 1 tie
xfeed_2421 0 1 decap_w0
xfeed_2420 0 1 decap_w0
xsubckt_309_and4_x1 0 1 439 1927 713 681 589 and4_x1
xsubckt_178_nand3_x0 0 1 580 714 1928 674 nand3_x0
xsubckt_1296_and2_x1 0 1 1287 435 1288 and2_x1
xsubckt_1479_nand3_x0 0 1 1117 498 211 1763 nand3_x0
xspare_buffer_38 0 1 65 68 buf_x4
xspare_buffer_39 0 1 15 16 buf_x4
.ends arlet6502_cts_r
