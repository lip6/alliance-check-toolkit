* BulkConn_1000WNoUp
* BulkConn_1000WNoUp
.subckt BulkConn_1000WNoUp vdd vss iovdd iovss

.ends BulkConn_1000WNoUp
