* DP8TArray_128X32
* DP8TCell
.subckt DP8TCell vdd vss wl1 wl2 bl1 bl1_n bl2 bl2_n
Mpu1 vdd bit_n bit vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpu2 vdd bit bit_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpd1 vss bit_n bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpd2 vss bit bit_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg1 bl1 wl1 bit vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg1n bl1_n wl1 bit_n vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg2 bl2 wl2 bit vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg2n bl2_n wl2 bit_n vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
.ends DP8TCell
* DP8TArray_2X1
.subckt DP8TArray_2X1 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 vdd vss wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
Xinst1x0 vdd vss wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
.ends DP8TArray_2X1
* DP8TArray_2X2
.subckt DP8TArray_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TArray_2X1
Xinst0x1 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X1
.ends DP8TArray_2X2
* DP8TArray_4X2
.subckt DP8TArray_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
.ends DP8TArray_4X2
* DP8TArray_4X4
.subckt DP8TArray_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X2
.ends DP8TArray_4X4
* DP8TArray_8X4
.subckt DP8TArray_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X4
.ends DP8TArray_8X4
* DP8TArray_8X8
.subckt DP8TArray_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X4
.ends DP8TArray_8X8
* DP8TArray_16X8
.subckt DP8TArray_16X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X8
.ends DP8TArray_16X8
* DP8TArray_16X16
.subckt DP8TArray_16X16 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_16X8
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X8
.ends DP8TArray_16X16
* DP8TArray_32X16
.subckt DP8TArray_32X16 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X16
Xinst1x0 vss vdd wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X16
.ends DP8TArray_32X16
* DP8TArray_32X32
.subckt DP8TArray_32X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_32X16
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X16
.ends DP8TArray_32X32
* DP8TArray_64X32
.subckt DP8TArray_64X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X32
Xinst1x0 vss vdd wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X32
.ends DP8TArray_64X32
* DP8TArray_128X32
.subckt DP8TArray_128X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_64X32
Xinst1x0 vss vdd wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_64X32
.ends DP8TArray_128X32
