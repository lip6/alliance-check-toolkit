-- no model for dffnr_x1
