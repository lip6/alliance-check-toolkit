* nexor2_x0
.subckt nexor2_x0 vdd vss i0 i1 nq
Mi0_nmos0 i0_n i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi0_pmos0 i0_n i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi0_nmos1 vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi0_pmos1 vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi1_n_nmos _net0 i1_n nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi1_pmos0 _net1 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi0_n_nmos nq i0_n _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi0_n_pmos nq i0_n _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi1_nmos0 _net2 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi1_n_pmos _net1 i1_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi1_nmos1 vss i1 i1_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi1_pmos1 vdd i1 i1_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends nexor2_x0
