* GuardRing_P18000W3888HFT
* GuardRing_P18000W3888HFT
.subckt GuardRing_P18000W3888HFT conn

.ends GuardRing_P18000W3888HFT
