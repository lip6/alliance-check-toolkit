* Filler2000
* Filler2000
.subckt Filler2000 vss vdd iovss iovdd

.ends Filler2000
