* diode_ss
.param
+ sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult = 1.1178e+00    
+ sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult = 1.0401e+00    
+ sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult = 1.234       
+ sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult = 1.189     
+ sky130_fd_pr__nfet_01v8__ajunction_mult = 1.1505e+0
+ sky130_fd_pr__nfet_01v8__pjunction_mult = 1.1793e+0
+ sky130_fd_pr__pfet_01v8__ajunction_mult = 1.0625
+ sky130_fd_pr__pfet_01v8__pjunction_mult = 1.0675
