* fill
.subckt fill vdd vss

.ends fill
