* Spice description of oa2a2a23_x4
* Spice driver version -71684325
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:30

* INTERF i0 i1 i2 i3 i4 i5 q vdd vss 


.subckt oa2a2a23_x4 6 5 8 9 10 13 4 1 15 
* NET 1 = vdd
* NET 4 = q
* NET 5 = i1
* NET 6 = i0
* NET 8 = i2
* NET 9 = i3
* NET 10 = i4
* NET 13 = i5
* NET 15 = vss
Mtr_00016 1 12 4 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00015 4 12 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00014 1 6 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 2 5 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 12 13 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 3 8 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 2 9 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 3 10 12 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 15 12 4 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00007 4 12 15 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00006 7 5 12 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 15 8 11 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 14 13 15 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 15 6 7 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 11 9 12 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 12 10 14 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C15 1 15 4.28155e-15
C14 2 15 8.47842e-16
C13 3 15 7.92919e-16
C12 4 15 2.15173e-15
C11 5 15 1.45223e-15
C10 6 15 1.4431e-15
C8 8 15 1.45223e-15
C7 9 15 1.46135e-15
C6 10 15 1.75227e-15
C4 12 15 3.29941e-15
C3 13 15 1.46135e-15
C1 15 15 3.36701e-15
.ends oa2a2a23_x4

