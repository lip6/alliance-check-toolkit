* Spice description of ao2o22_x4
* Spice driver version -781979877
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:37

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt ao2o22_x4 9 8 6 5 4 3 7 
* NET 3 = vdd
* NET 4 = q
* NET 5 = i3
* NET 6 = i2
* NET 7 = vss
* NET 8 = i1
* NET 9 = i0
Mtr_00012 3 10 4 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 4 10 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 3 5 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00009 1 6 10 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00008 10 8 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00007 2 9 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00006 7 10 4 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 4 10 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 11 5 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00003 7 6 11 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00002 11 8 10 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00001 10 9 11 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
C9 3 7 3.58487e-15
C8 4 7 2.15173e-15
C7 5 7 1.96725e-15
C6 6 7 1.86548e-15
C5 7 7 2.90768e-15
C4 8 7 1.79868e-15
C3 9 7 1.49465e-15
C2 10 7 3.27621e-15
C1 11 7 7.92919e-16
.ends ao2o22_x4

