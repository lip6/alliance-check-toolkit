* This spice netlist for sff1r_x4 is made manually based on sff1_x4 extracted
* netlist.
* Inverter in master latch with y as output has been replaced with nand2.
*   orig: y <= NOT sff_m;
*    new: y <= NOT (sff_m and nrst);
* Tri-state inverter in slave latch has been replaced with tri-state nand2.
*   orig: sff_s <= NOT q WHEN nckr ELSE 'Z';
*    new: sff_s <= NOT (q and nrst) WHEN nckr ELSE 'Z'

* INTERF ck i nrst q vdd vss 


.subckt sff1_x4 ck i nrst q vdd vss 

Mtr_00014 nckr ck vdd vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00008 vss ck nckr vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 
Mtr_00015 vdd nckr ckr vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00001 ckr nckr vss vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 

Mtr_00023 u i vdd vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00009 vss i u vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 

Mtr_00024 vdd u 2 vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00016 2 ckr sff_m vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00002 11 u vss vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 
Mtr_00007 sff_m nckr 11 vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 

# NAND2; replaces INV
# - input: sff_m, nrst
# - output y
Mtr_00026 y sff_m vdd vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00026b y nrst vdd vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00012 y sff_m y2 vss tn L=0.05U W=0.44U AS=0.022P AD=0.022P PS=0.65U PD=0.65U 
Mtr_00012b y2 nrst vss vss tn L=0.05U W=0.44U AS=0.022P AD=0.022P PS=0.65U PD=0.65U 

Mtr_00017 3 y vdd vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00022 sff_m nckr 3 vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00013 vss y 9 vss tn L=0.05U W=0.22U AS=0.022P AD=0.022P PS=0.65U PD=0.65U 
Mtr_00003 9 ckr sff_m vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 

Mtr_00021 y nckr sff_s vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00004 sff_s ckr y vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 

Mtr_00025 q sff_s vdd vdd tp L=0.05U W=1U AS=0.1P AD=0.1P PS=2.2U PD=2.2U 
Mtr_00018 vdd sff_s q vdd tp L=0.05U W=1U AS=0.1P AD=0.1P PS=2.2U PD=2.2U 
Mtr_00011 q sff_s vss vss tn L=0.05U W=0.47U AS=0.047P AD=0.047P PS=1.15U PD=1.15U 
Mtr_00010 vss sff_s q vss tn L=0.05U W=0.47U AS=0.047P AD=0.047P PS=1.15U PD=1.15U 

# tri-state NAND2; replaces TRI-INV
# - input: q, nrst
# - enable: nckr
# - output: sff_s
Mtr_00019 sff_s_p q vdd vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00019b sff_s_p nrst vdd vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00020 sff_s ckr sff_s_p vdd tp L=0.05U W=0.5U AS=0.05P AD=0.05P PS=1.2U PD=1.2U 
Mtr_00005 sff_s_n nckr sff_s vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 
Mtr_00006 sff_s_n nrst sff_s_n2 vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 
Mtr_00006b sff_s_n2 q vss vss tn L=0.05U W=0.25U AS=0.025P AD=0.025P PS=0.7U PD=0.7U 

C14 vdd vss 9.25562e-16
C13 q vss 7.48882e-16
C11 sff_s vss 7.24108e-16
C10 y vss 4.62063e-16
C8 sff_m vss 6.08385e-16
C6 i vss 5.2061e-16
C5 u vss 5.95978e-16
C4 ck vss 5.56318e-16
C3 nckr vss 1.59449e-15
C2 vss vss 8.01335e-16
C1 ckr vss 1.31048e-15
.ends sff1_x4

