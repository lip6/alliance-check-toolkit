* Spice description of oa2a2a2a24_x2
* Spice driver version -2025853157
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:31

* INTERF i0 i1 i2 i3 i4 i5 i6 i7 q vdd vss 


.subckt oa2a2a2a24_x2 5 6 9 10 12 13 16 17 8 2 19 
* NET 2 = vdd
* NET 5 = i0
* NET 6 = i1
* NET 8 = q
* NET 9 = i2
* NET 10 = i3
* NET 12 = i4
* NET 13 = i5
* NET 16 = i6
* NET 17 = i7
* NET 19 = vss
Mtr_00018 8 15 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00017 4 16 15 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00016 2 5 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00015 1 6 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00014 3 9 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 1 10 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 3 12 4 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 4 13 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 15 17 4 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 8 15 19 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00008 15 16 18 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00007 19 5 7 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00006 7 6 15 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 19 9 11 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 11 10 15 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 15 12 14 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 14 13 19 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 18 17 19 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C19 1 19 7.71835e-16
C18 2 19 4.01809e-15
C17 3 19 1.05722e-15
C16 4 19 1.33673e-15
C15 5 19 1.69828e-15
C14 6 19 1.38512e-15
C12 8 19 1.9237e-15
C11 9 19 1.38512e-15
C10 10 19 1.39425e-15
C8 12 19 1.39425e-15
C7 13 19 1.38512e-15
C5 15 19 3.25034e-15
C4 16 19 1.49829e-15
C3 17 19 1.69828e-15
C1 19 19 3.58313e-15
.ends oa2a2a2a24_x2

