* Spice description of ao22_x4
* Spice driver version 1987985179
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:35

* INTERF i0 i1 i2 q vdd vss 


.subckt ao22_x4 7 6 4 3 2 5 
* NET 2 = vdd
* NET 3 = q
* NET 4 = i2
* NET 5 = vss
* NET 6 = i1
* NET 7 = i0
Mtr_00010 2 8 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 3 8 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 2 4 8 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 8 6 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 1 7 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00005 5 8 3 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00004 3 8 5 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00003 5 4 9 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00002 9 6 8 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00001 8 7 9 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
C8 2 5 3.74455e-15
C7 3 5 2.15173e-15
C6 4 5 2.15293e-15
C5 5 5 2.78442e-15
C4 6 5 1.69381e-15
C3 7 5 1.37606e-15
C2 8 5 2.27276e-15
C1 9 5 4.83008e-16
.ends ao22_x4

