* IOPadAnalog
.subckt IOPadAnalog vss vdd iovss iovdd pad padres
Xpad pad Pad_15800W12000H
Xnclamp iovss iovdd pad Clamp_N12N0D
Xpclamp iovss iovdd pad Clamp_P12N0D
Xsecondprot iovdd iovss pad padres SecondaryProtection
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadAnalog
