* Spice description of on12_x1
* Spice driver version -845959397
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:37

* INTERF i0 i1 q vdd vss 


.subckt on12_x1 2 5 3 1 7 
* NET 1 = vdd
* NET 2 = i0
* NET 3 = q
* NET 5 = i1
* NET 7 = vss
Mtr_00006 3 6 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00005 1 5 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00004 1 2 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00003 4 6 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00002 7 5 6 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00001 3 2 4 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
C7 1 7 1.46971e-15
C6 2 7 2.05116e-15
C5 3 7 2.28266e-15
C3 5 7 1.97952e-15
C2 6 7 1.48193e-15
C1 7 7 1.64625e-15
.ends on12_x1

