-- no model for buf_x4
