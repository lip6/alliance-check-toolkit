-- no model for dff_x1
