* Spice description of nmx2_x4
* Spice driver version 553643803
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:58

* INTERF cmd i0 i1 nq vdd vss 


.subckt nmx2_x4 11 7 5 4 3 13 
* NET 3 = vdd
* NET 4 = nq
* NET 5 = i1
* NET 7 = i0
* NET 11 = cmd
* NET 13 = vss
Mtr_00016 4 6 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00015 3 6 4 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00014 6 10 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.29U AS=0.5496P AD=0.5496P PS=5.07U PD=5.07U 
Mtr_00013 3 11 12 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.29U AS=0.5496P AD=0.5496P PS=5.07U PD=5.07U 
Mtr_00012 3 5 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.29U AS=0.5496P AD=0.5496P PS=5.07U PD=5.07U 
Mtr_00011 2 12 10 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.29U AS=0.5496P AD=0.5496P PS=5.07U PD=5.07U 
Mtr_00010 10 11 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.29U AS=0.5496P AD=0.5496P PS=5.07U PD=5.07U 
Mtr_00009 1 7 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.29U AS=0.5496P AD=0.5496P PS=5.07U PD=5.07U 
Mtr_00008 4 6 13 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00007 13 6 4 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00006 6 10 13 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00005 13 11 12 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00004 13 5 9 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00003 8 7 13 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00002 10 12 8 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00001 9 11 10 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
C11 3 13 4.50778e-15
C10 4 13 2.15173e-15
C9 5 13 2.42347e-15
C8 6 13 2.10853e-15
C7 7 13 2.1073e-15
C4 10 13 1.88346e-15
C3 11 13 2.95155e-15
C2 12 13 2.89635e-15
C1 13 13 3.69377e-15
.ends nmx2_x4

