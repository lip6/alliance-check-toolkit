-- no model for tie_diff_w2
