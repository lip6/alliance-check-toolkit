* Spice description of an12_x4
* Spice driver version 1982746395
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:33

* INTERF i0 i1 q vdd vss 


.subckt an12_x4 6 2 5 1 7 
* NET 1 = vdd
* NET 2 = i1
* NET 5 = q
* NET 6 = i0
* NET 7 = vss
Mtr_00010 1 4 5 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 5 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 1 2 4 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 4 8 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 1 6 8 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 7 4 5 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 5 4 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 7 2 3 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 3 8 4 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 7 6 8 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C8 1 7 2.99804e-15
C7 2 7 2.25616e-15
C5 4 7 2.00816e-15
C4 5 7 2.25814e-15
C3 6 7 1.90058e-15
C2 7 7 2.39685e-15
C1 8 7 1.86209e-15
.ends an12_x4

