-- no model for or21nand_x1
