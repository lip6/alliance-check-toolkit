* Spice description of oa3ao322_x4
* Spice driver version -2006802661
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:36

* INTERF i0 i1 i2 i3 i4 i5 i6 q vdd vss 


.subckt oa3ao322_x4 12 11 7 8 5 6 9 16 4 17 
* NET 4 = vdd
* NET 5 = i4
* NET 6 = i5
* NET 7 = i2
* NET 8 = i3
* NET 9 = i6
* NET 11 = i1
* NET 12 = i0
* NET 16 = q
* NET 17 = vss
Mtr_00018 15 9 3 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00017 3 7 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00016 4 11 3 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00015 3 12 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00014 4 15 16 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 16 15 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 2 8 15 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00011 3 6 1 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00010 1 5 2 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00009 15 7 14 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.36U AS=0.3264P AD=0.3264P PS=3.2U PD=3.2U 
Mtr_00008 10 5 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.68U AS=0.1632P AD=0.1632P PS=1.84U PD=1.84U 
Mtr_00007 17 6 10 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.68U AS=0.1632P AD=0.1632P PS=1.84U PD=1.84U 
Mtr_00006 17 8 10 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00005 10 9 15 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00004 14 11 13 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.36U AS=0.3264P AD=0.3264P PS=3.2U PD=3.2U 
Mtr_00003 13 12 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.36U AS=0.3264P AD=0.3264P PS=3.2U PD=3.2U 
Mtr_00002 16 15 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00001 17 15 16 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
C15 3 17 1.30977e-15
C14 4 17 4.28319e-15
C13 5 17 1.74392e-15
C12 6 17 1.7713e-15
C11 7 17 1.51898e-15
C10 8 17 1.7713e-15
C9 9 17 1.40032e-15
C8 10 17 5.74217e-16
C7 11 17 1.86578e-15
C6 12 17 1.86578e-15
C3 15 17 3.09325e-15
C2 16 17 2.15173e-15
C1 17 17 3.87031e-15
.ends oa3ao322_x4

