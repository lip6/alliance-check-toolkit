* Spice description of mx3_x4
* Spice driver version 311590683
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:47

* INTERF cmd0 cmd1 i0 i1 i2 q vdd vss 


.subckt mx3_x4 9 17 6 8 12 7 5 19 
* NET 5 = vdd
* NET 6 = i0
* NET 7 = q
* NET 8 = i1
* NET 9 = cmd0
* NET 12 = i2
* NET 17 = cmd1
* NET 19 = vss
Mtr_00022 5 15 7 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00021 5 9 10 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00020 7 15 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00019 4 8 3 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00018 15 6 1 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00017 3 16 15 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00016 5 10 4 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00015 1 9 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00014 2 12 4 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00013 16 17 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00012 15 17 2 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00011 19 15 7 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00010 19 9 10 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.51U AS=0.1224P AD=0.1224P PS=1.5U PD=1.5U 
Mtr_00009 7 15 19 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00008 11 10 19 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00007 16 17 19 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.68U AS=0.1632P AD=0.1632P PS=1.84U PD=1.84U 
Mtr_00006 14 12 18 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00005 15 16 14 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00004 13 17 15 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00003 18 8 13 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00002 15 6 11 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00001 19 9 18 19 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
C16 4 19 8.3264e-16
C15 5 19 4.93427e-15
C14 6 19 1.47501e-15
C13 7 19 2.41603e-15
C12 8 19 1.0671e-15
C11 9 19 1.95732e-15
C10 10 19 2.13754e-15
C8 12 19 1.08148e-15
C5 15 19 4.22605e-15
C4 16 19 1.81503e-15
C3 17 19 2.88805e-15
C2 18 19 8.02238e-16
C1 19 19 4.61847e-15
.ends mx3_x4

