* SP6TArray_2X1
* SP6TCell
.subckt SP6TCell vdd vss wl bl bl_n
Mpu1 vdd bit_n bit vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpu2 bit_n bit vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpd1 vss bit_n bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpd2 bit_n bit vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg1 bl wl bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg2 bl_n wl bit_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
.ends SP6TCell
* SP6TArray_2X1
.subckt SP6TArray_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 vdd vss wl[0] bl[0] bl_n[0] SP6TCell
Xinst1x0 vdd vss wl[1] bl[0] bl_n[0] SP6TCell
.ends SP6TArray_2X1
