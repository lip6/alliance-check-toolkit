* Spice description of noa2ao222_x4
* Spice driver version -90042597
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:14

* INTERF i0 i1 i2 i3 i4 nq vdd vss 


.subckt noa2ao222_x4 10 11 7 5 8 4 3 14 
* NET 3 = vdd
* NET 4 = nq
* NET 5 = i3
* NET 7 = i2
* NET 8 = i4
* NET 10 = i0
* NET 11 = i1
* NET 14 = vss
Mtr_00016 2 5 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00015 2 11 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00014 3 6 4 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 4 6 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 1 7 13 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 13 8 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 3 10 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00009 3 13 6 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00008 14 6 4 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 4 6 14 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 9 5 14 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00005 14 7 9 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00004 9 8 13 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00003 12 10 14 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00002 13 11 12 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00001 14 13 6 14 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C13 2 14 1.09695e-15
C12 3 14 4.29251e-15
C11 4 14 2.20321e-15
C10 5 14 1.06552e-15
C9 6 14 1.45604e-15
C8 7 14 1.36955e-15
C7 8 14 1.38512e-15
C6 9 14 7.41432e-16
C5 10 14 1.62526e-15
C4 11 14 1.71653e-15
C2 13 14 2.76159e-15
C1 14 14 4.56026e-15
.ends noa2ao222_x4

