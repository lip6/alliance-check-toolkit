-- no model for fill
