* tie_w4
* tie_w4
.subckt tie_w4 vdd vss

.ends tie_w4
