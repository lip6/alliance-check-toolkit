-- no model for tie_w2
