-- no model for nsnrlatch_x1
