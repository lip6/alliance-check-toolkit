* IOPadAnalog
.subckt IOPadAnalog vss vdd iovss iovdd pad padres
Xpad pad Pad_15800W12000H
Xnclamp iovss iovdd pad Clamp_N12N0D
Xpclamp iovss iovdd pad Clamp_P12N0D
Xbulkconn vdd vss iovdd iovss BulkConn_18000WUp
Xsecondprot iovdd iovss pad padres SecondaryProtection
.ends IOPadAnalog
