-- no model for or3_x1
