-- no model for tie_w4
