* Spice description of o2_x4
* Spice driver version 562732827
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:21

* INTERF i0 i1 q vdd vss 


.subckt o2_x4 3 5 4 1 6 
* NET 1 = vdd
* NET 3 = i0
* NET 4 = q
* NET 5 = i1
* NET 6 = vss
Mtr_00009 1 7 4 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 4 7 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 2 5 7 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00006 1 3 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00005 6 7 4 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 4 7 6 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 6 3 7 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 7 5 6 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 6 3 7 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C7 1 6 2.38589e-15
C5 3 6 2.33831e-15
C4 4 6 2.15173e-15
C3 5 6 1.81693e-15
C2 6 6 2.25839e-15
C1 7 6 2.18167e-15
.ends o2_x4

