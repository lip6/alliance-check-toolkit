* Spice description of oa22_x4
* Spice driver version 1499328283
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:26

* INTERF i0 i1 i2 q vdd vss 


.subckt oa22_x4 7 6 4 3 2 9 
* NET 2 = vdd
* NET 3 = q
* NET 4 = i2
* NET 6 = i1
* NET 7 = i0
* NET 9 = vss
Mtr_00010 3 5 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 2 5 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 1 6 5 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 2 4 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 5 7 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00005 9 5 3 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 3 5 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 8 7 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 5 6 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 9 4 5 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C9 1 9 4.9821e-16
C8 2 9 2.87563e-15
C7 3 9 2.15173e-15
C6 4 9 2.38394e-15
C5 5 9 2.16779e-15
C4 6 9 1.86716e-15
C3 7 9 1.90821e-15
C1 9 9 2.52011e-15
.ends oa22_x4

