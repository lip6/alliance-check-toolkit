* Gallery
.subckt Gallery vdd vss iovdd iopadin_pad iopadout_pad iopadtriout_pad iopadinout_pad iopadin_p2c iopadinout_p2c iopadout_c2p iopadtriout_c2p iopadinout_c2p iopadtriout_c2p_en iopadinout_c2p_en ana_out ana_outres
Xcorner vss vdd vss iovdd Corner
Xfiller200 vss vdd vss iovdd Filler200
Xfiller400 vss vdd vss iovdd Filler400
Xfiller1000 vss vdd vss iovdd Filler1000
Xfiller2000 vss vdd vss iovdd Filler2000
Xfiller4000 vss vdd vss iovdd Filler4000
Xfiller10000 vss vdd vss iovdd Filler10000
Xiopadvss vss vdd vss iovdd IOPadVss
Xiopadvdd vss vdd vss iovdd IOPadVdd
Xiopadin vss vdd vss iovdd iopadin_p2c iopadin_pad IOPadIn
Xiopadout vss vdd vss iovdd iopadout_c2p iopadout_pad IOPadOut
Xiopadtriout vss vdd vss iovdd iopadtriout_c2p iopadtriout_c2p_en iopadtriout_pad IOPadTriOut
Xiopadinout vss vdd vss iovdd iopadinout_p2c iopadinout_c2p iopadinout_c2p_en iopadinout_pad IOPadInOut
Xiopadiovss vss vdd vss iovdd IOPadIOVss
Xiopadiovdd vss vdd vss iovdd IOPadIOVdd
Xiopadanalog vss vdd vss iovdd ana_out ana_outres IOPadAnalog
Xcorner2 vss vdd vss iovdd Corner
.ends Gallery
