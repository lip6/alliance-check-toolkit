* Spice description of a4_x4
* Spice driver version 526434075
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:32

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt a4_x4 7 8 4 3 2 1 11 
* NET 1 = vdd
* NET 2 = q
* NET 3 = i3
* NET 4 = i2
* NET 7 = i0
* NET 8 = i1
* NET 11 = vss
Mtr_00012 1 5 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 1 3 5 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00010 5 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00009 1 8 5 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00008 5 7 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00007 2 5 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 11 5 2 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 2 5 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 5 3 6 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00003 6 4 10 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00002 9 7 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00001 10 8 9 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
C11 1 11 3.80192e-15
C10 2 11 2.15173e-15
C9 3 11 1.44901e-15
C8 4 11 1.75304e-15
C7 5 11 2.58332e-15
C5 7 11 1.40338e-15
C4 8 11 1.72566e-15
C1 11 11 2.73293e-15
.ends a4_x4

