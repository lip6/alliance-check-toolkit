* and2_x1
.subckt and2_x1 vdd vss q i0 i1
Mi0_nmos nq i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos _net0 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mn_pd vss nq q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mq_pu vdd nq q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends and2_x1
