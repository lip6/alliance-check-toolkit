* Spice description of no2_x4
* Spice driver version -1070620901
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:01

* INTERF i0 i1 nq vdd vss 


.subckt no2_x4 5 6 4 1 8 
* NET 1 = vdd
* NET 4 = nq
* NET 5 = i0
* NET 6 = i1
* NET 8 = vss
Mtr_00010 1 3 4 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 4 3 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 3 7 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 1 5 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 2 6 7 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 3 7 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00004 8 3 4 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 4 3 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 8 5 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 7 6 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C8 1 8 1.95945e-15
C6 3 8 1.93514e-15
C5 4 8 1.6579e-15
C4 5 8 1.78042e-15
C3 6 8 1.76217e-15
C2 7 8 2.78651e-15
C1 8 8 2.36645e-15
.ends no2_x4

