* Spice description of a2_x2
* Spice driver version -173076709
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:27

* INTERF i0 i1 q vdd vss 


.subckt a2_x2 5 2 3 1 4 
* NET 1 = vdd
* NET 2 = i1
* NET 3 = q
* NET 4 = vss
* NET 5 = i0
Mtr_00006 3 7 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 1 2 7 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00004 7 5 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00003 3 7 4 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 6 5 7 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 4 2 6 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C7 1 4 1.58611e-15
C6 2 4 2.49032e-15
C5 3 4 2.15173e-15
C4 4 4 1.33112e-15
C3 5 4 1.70216e-15
C1 7 4 1.83178e-15
.ends a2_x2

