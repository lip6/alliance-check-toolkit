-- no model for powmid_x0
