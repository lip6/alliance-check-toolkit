* Spice description of nao22_x4
* Spice driver version 1492225819
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:54

* INTERF i0 i1 i2 nq vdd vss 


.subckt nao22_x4 6 5 8 4 2 10 
* NET 2 = vdd
* NET 4 = nq
* NET 5 = i1
* NET 6 = i0
* NET 8 = i2
* NET 10 = vss
Mtr_00012 2 3 4 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 4 3 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 1 5 7 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00009 2 6 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00008 7 8 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 2 7 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 4 3 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 10 3 4 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 7 5 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00003 9 8 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 9 6 7 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 10 7 3 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C9 2 10 4.10186e-15
C8 3 10 1.78987e-15
C7 4 10 2.15173e-15
C6 5 10 1.6436e-15
C5 6 10 1.65894e-15
C4 7 10 2.73442e-15
C3 8 10 2.4615e-15
C2 9 10 5.28612e-16
C1 10 10 3.2126e-15
.ends nao22_x4

