* Spice description of oa2a2a23_x2
* Spice driver version -1686868197
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:29

* INTERF i0 i1 i2 i3 i4 i5 q vdd vss 


.subckt oa2a2a23_x2 5 6 8 10 9 13 4 1 15 
* NET 1 = vdd
* NET 4 = q
* NET 5 = i0
* NET 6 = i1
* NET 8 = i2
* NET 9 = i4
* NET 10 = i3
* NET 13 = i5
* NET 15 = vss
Mtr_00014 4 12 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 3 8 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 1 5 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 2 6 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 12 13 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 3 9 12 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 2 10 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 4 12 15 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00006 15 8 11 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 15 5 7 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 7 6 12 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 14 13 15 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 12 9 14 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 11 10 12 15 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C15 1 15 3.60092e-15
C14 2 15 8.47842e-16
C13 3 15 8.0812e-16
C12 4 15 2.21103e-15
C11 5 15 1.39425e-15
C10 6 15 1.38512e-15
C8 8 15 1.42809e-15
C7 9 15 1.69828e-15
C6 10 15 1.38512e-15
C4 12 15 3.04153e-15
C3 13 15 1.38512e-15
C1 15 15 3.0419e-15
.ends oa2a2a23_x2

