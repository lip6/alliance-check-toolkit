* Spice description of a3_x2
* Spice driver version -161280229
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:29

* INTERF i0 i1 i2 q vdd vss 


.subckt a3_x2 5 6 2 3 1 4 
* NET 1 = vdd
* NET 2 = i2
* NET 3 = q
* NET 4 = vss
* NET 5 = i0
* NET 6 = i1
Mtr_00008 3 9 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 1 2 9 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00006 9 6 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00005 1 5 9 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00004 3 9 4 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00003 4 2 8 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00002 7 5 9 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00001 8 6 7 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
C9 1 4 2.18239e-15
C8 2 4 1.34257e-15
C7 3 4 2.15173e-15
C6 4 4 1.71458e-15
C5 5 4 1.34257e-15
C4 6 4 1.36995e-15
C1 9 4 2.46382e-15
.ends a3_x2

