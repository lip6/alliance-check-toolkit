* Spice description of sff1r_x4
* Spice driver version -779358437
* Date ( dd/mm/yyyy hh:mm:ss ): 29/07/2024 at 18:03:57

* INTERF ck i nrst q vdd vss 


.subckt sff1r_x4 17 14 7 5 4 18 
* NET 4 = vdd
* NET 5 = q
* NET 7 = nrst
* NET 8 = sff_s
* NET 10 = y
* NET 11 = sff_m
* NET 14 = i
* NET 15 = ckr
* NET 17 = ck
* NET 18 = vss
* NET 19 = nckr
Mtr_00028 5 8 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_00027 8 15 1 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_00026 4 8 5 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_00025 1 5 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_00024 10 19 8 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_00023 4 7 10 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00022 11 19 3 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00021 3 10 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00020 10 11 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00019 2 15 11 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00018 4 16 2 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00017 16 14 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00016 4 19 15 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00015 19 17 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00014 18 8 5 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00013 5 8 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00012 18 5 6 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00011 6 19 8 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00010 8 15 10 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00009 10 7 9 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00008 9 11 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00007 18 10 12 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00006 12 15 11 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00005 11 19 13 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00004 13 16 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00003 18 17 19 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00002 15 19 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00001 18 14 16 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
.ends sff1r_x4

