(* blackbox = 1 *)
module spblock_512w64b8w(input [8:0] a,
			 input [63:0] d,
			 output [63:0] q,
			 input [7:0] we,
			 input clk);
endmodule // SPBlock_512W64B8W
