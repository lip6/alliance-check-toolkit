* Spice description of o4_x4
* Spice driver version -467919077
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:25

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt o4_x4 8 9 7 6 5 1 11 
* NET 1 = vdd
* NET 5 = q
* NET 6 = i3
* NET 7 = i2
* NET 8 = i0
* NET 9 = i1
* NET 11 = vss
Mtr_00012 5 10 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 1 10 5 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 1 6 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 2 7 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 3 8 4 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 4 9 10 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 5 10 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 11 10 5 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 11 6 10 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 10 7 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 11 8 10 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 10 9 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C11 1 11 2.67213e-15
C7 5 11 2.18213e-15
C6 6 11 1.71653e-15
C5 7 11 2.01143e-15
C4 8 11 2.00231e-15
C3 9 11 2.00231e-15
C2 10 11 3.20087e-15
C1 11 11 2.30729e-15
.ends o4_x4

