* SP6TWriteDriver_4M2B
* inv_x0
.subckt inv_x0 vdd vss i nq
Mn vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends inv_x0
* nor2_x0
.subckt nor2_x0 vdd vss nq i0 i1
Mn0 vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp0 vdd i0 int0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn1 nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp1 int0 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
.ends nor2_x0
* sff1_x4
.subckt sff1_x4 vdd ck vss i q
Mp_ck nckr ck vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_ck nckr ck vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ckr_1 _net1 ckr sff_m vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_ckr_2 y ckr sff_s vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_ckr_1 sff_m ckr _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ckr_2 sff_s ckr _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i u i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i u i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_2 sff_m nckr _net5 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_3 y nckr sff_s vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_1 vdd nckr ckr vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nckr_1 vss nckr ckr vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nckr_3 sff_s nckr _net6 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nckr_2 _net2 nckr sff_m vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_q_1 _net6 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_q_1 _net0 q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_sffm_1 vss sff_m y vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_sffm_1 vdd sff_m y vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_sffs_1 vdd sff_s q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_sffs_1 vss sff_s q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mn_sffs_2 q sff_s vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_sffs_2 q sff_s vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_u vss u _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_u vdd u _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_y_1 _net4 y vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_y_1 _net5 y vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends sff1_x4
* SP6TWriteDriver_4M2B
.subckt SP6TWriteDriver_4M2B vss vdd clk we_n bl[0] bl_n[0] d[0] bl[1] bl_n[1] d[1]
Xff[0] vdd clk vss d[0] d_latched[0] sff1_x4
Xff[1] vdd clk vss d[1] d_latched[1] sff1_x4
Xnora[0] vdd vss bl_drive[0] d_latched[0] we_n nor2_x0
Xnora[1] vdd vss bl_drive[1] d_latched[1] we_n nor2_x0
Xinv[0] vdd vss d_latched[0] d_n[0] inv_x0
Xinv[1] vdd vss d_latched[1] d_n[1] inv_x0
Xnorb[0] vdd vss bln_drive[0] d_n[0] we_n nor2_x0
Xnorb[1] vdd vss bln_drive[1] d_n[1] we_n nor2_x0
Mblpd[0] vss bl_drive[0] bl[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblpd[1] vss bl_drive[1] bl[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblnpd[0] bl_n[0] bln_drive[0] vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblnpd[1] bl_n[1] bln_drive[1] vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
.ends SP6TWriteDriver_4M2B
