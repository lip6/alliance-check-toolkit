* Spice description of noa22_x4
* Spice driver version -110084325
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:06

* INTERF i0 i1 i2 nq vdd vss 


.subckt noa22_x4 4 6 7 3 2 10 
* NET 2 = vdd
* NET 3 = nq
* NET 4 = i0
* NET 6 = i1
* NET 7 = i2
* NET 10 = vss
Mtr_00012 2 5 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 2 9 5 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00010 1 4 9 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00009 9 6 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00008 1 7 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00007 3 5 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 10 5 3 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 10 9 5 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00004 10 4 8 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3048P AD=0.3048P PS=3.03U PD=3.03U 
Mtr_00003 8 6 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3048P AD=0.3048P PS=3.03U PD=3.03U 
Mtr_00002 9 7 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3048P AD=0.3048P PS=3.03U PD=3.03U 
Mtr_00001 3 5 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C10 1 10 4.52605e-16
C9 2 10 3.57898e-15
C8 3 10 2.18213e-15
C7 4 10 1.9478e-15
C6 5 10 1.87148e-15
C5 6 10 2.01773e-15
C4 7 10 1.79868e-15
C2 9 10 2.32081e-15
C1 10 10 3.10817e-15
.ends noa22_x4

