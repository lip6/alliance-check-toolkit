* top_hitas_eldo.cir bench SARlogic
* 

*****************

.TEMP 25
.GLOBAL VDD VSS
Vsupply vdd 0  DC 1.8
Vground vss 0  DC 0

******************
* circuit model
* include standard cells
.INCLUDE /users/soft/techno/techno/pdkmaster/views/tsmc_c018/FlexLib/spice/FlexLib.spi

* include circuit netlist
.INCLUDE SARlogic_netlist.spi

*****************
* NET     0 = vss
* NET     1 = vdd
* NET     2 = rst
* NET    27 = res[7]
* NET    28 = res[6]
* NET    29 = res[5]
* NET    30 = res[4]
* NET    31 = res[3]
* NET    32 = res[2]
* NET    33 = res[1]
* NET    34 = res[0]
* NET    45 = cmp
* NET    46 = clk
* NET   144 = SOC
* NET   146 = SE
* NET   148 = EOC
* NET   157 = DAC_control[7]
* NET   158 = DAC_control[6]
* NET   159 = DAC_control[5]
* NET   160 = DAC_control[4]
* NET   161 = DAC_control[3]
* NET   162 = DAC_control[2]
* NET   163 = DAC_control[1]
* NET   164 = DAC_control[0]

*SARlogic 0 1 2 27 28 29 30 31 32 33 34 45 46 144 146 148 157 158 159 160 161 162 163 164

*load on outputs

.end
