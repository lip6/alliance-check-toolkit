* SP6TColumnBlock_128R64B4M8W
.subckt SP6TColumnBlock_128R64B4M8W vss vdd clk precharge_n we_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] mux[0] mux[1] mux[2] mux[3] we[0] q[0] d[0] q[1] d[1] q[2] d[2] q[3] d[3] q[4] d[4] q[5] d[5] q[6] d[6] q[7] d[7] we[1] q[8] d[8] q[9] d[9] q[10] d[10] q[11] d[11] q[12] d[12] q[13] d[13] q[14] d[14] q[15] d[15] we[2] q[16] d[16] q[17] d[17] q[18] d[18] q[19] d[19] q[20] d[20] q[21] d[21] q[22] d[22] q[23] d[23] we[3] q[24] d[24] q[25] d[25] q[26] d[26] q[27] d[27] q[28] d[28] q[29] d[29] q[30] d[30] q[31] d[31] we[4] q[32] d[32] q[33] d[33] q[34] d[34] q[35] d[35] q[36] d[36] q[37] d[37] q[38] d[38] q[39] d[39] we[5] q[40] d[40] q[41] d[41] q[42] d[42] q[43] d[43] q[44] d[44] q[45] d[45] q[46] d[46] q[47] d[47] we[6] q[48] d[48] q[49] d[49] q[50] d[50] q[51] d[51] q[52] d[52] q[53] d[53] q[54] d[54] q[55] d[55] we[7] q[56] d[56] q[57] d[57] q[58] d[58] q[59] d[59] q[60] d[60] q[61] d[61] q[62] d[62] q[63] d[63]
Xcolumn[0] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[0] d[0] q[1] d[1] q[2] d[2] q[3] d[3] q[4] d[4] q[5] d[5] q[6] d[6] q[7] d[7] we[0] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[1] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[8] d[8] q[9] d[9] q[10] d[10] q[11] d[11] q[12] d[12] q[13] d[13] q[14] d[14] q[15] d[15] we[1] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[2] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[16] d[16] q[17] d[17] q[18] d[18] q[19] d[19] q[20] d[20] q[21] d[21] q[22] d[22] q[23] d[23] we[2] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[3] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[24] d[24] q[25] d[25] q[26] d[26] q[27] d[27] q[28] d[28] q[29] d[29] q[30] d[30] q[31] d[31] we[3] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[4] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[32] d[32] q[33] d[33] q[34] d[34] q[35] d[35] q[36] d[36] q[37] d[37] q[38] d[38] q[39] d[39] we[4] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[5] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[40] d[40] q[41] d[41] q[42] d[42] q[43] d[43] q[44] d[44] q[45] d[45] q[46] d[46] q[47] d[47] we[5] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[6] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[48] d[48] q[49] d[49] q[50] d[50] q[51] d[51] q[52] d[52] q[53] d[53] q[54] d[54] q[55] d[55] we[6] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[7] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[56] d[56] q[57] d[57] q[58] d[58] q[59] d[59] q[60] d[60] q[61] d[61] q[62] d[62] q[63] d[63] we[7] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
.ends SP6TColumnBlock_128R64B4M8W
