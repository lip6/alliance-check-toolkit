* tie_poly
* tie_poly
.subckt tie_poly vdd vss

.ends tie_poly
