* GuardRing_P12310W3968HFT
* GuardRing_P12310W3968HFT
.subckt GuardRing_P12310W3968HFT conn

.ends GuardRing_P12310W3968HFT
