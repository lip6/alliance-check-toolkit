../rtl/cpu.vhdl