*
* sample.spi
* 
*.INCLUDE ./techno/bsim4_dummy.hsp
*.INCLUDE ./techno/bsim4_dummy.ng

.TEMP 125
Vground gnd 0 DC 0
Vsupply vdd 0 DC 1.62

.subckt inv a y vdd gnd
MM02 y   a   gnd gnd tn L=0.18U W=1.15U AS=0.414P AD=0.414P PS=3.02U PD=3.02U
MM03 y   a   vdd vdd tp L=0.18U W=2.23U AS=0.8028P AD=0.8028P PS=5.18U PD=5.18U
.ends

.subckt inv_chain in out vdd gnd
Xa in 1 vdd gnd inv
Xb 1  2 vdd gnd inv
Xc 2  3 vdd gnd inv
Xd 3  4 vdd gnd inv
Xe 4  out vdd gnd inv
.ends

Xch in out vdd gnd inv_chain
