* Spice description of na2_x1
* Spice driver version -93352165
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:48

* INTERF i0 i1 nq vdd vss 


.subckt na2_x1 4 2 3 1 6 
* NET 1 = vdd
* NET 2 = i1
* NET 3 = nq
* NET 4 = i0
* NET 6 = vss
Mtr_00004 1 2 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00003 3 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00002 3 2 5 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00001 5 4 6 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
C6 1 6 1.63184e-15
C5 2 6 1.80296e-15
C4 3 6 2.22185e-15
C3 4 6 1.84551e-15
C1 6 6 1.32537e-15
.ends na2_x1

