* nand3_x0
.subckt nand3_x0 vdd vss nq i0 i1 i2
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi1_nmos _net0 i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi2_nmos _net1 i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi2_pmos vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends nand3_x0
