* diode_fs
.param
+ sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult = 1.1756e+00    
+ sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult = 1.0618e+00    
+ sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult = 1.3319      
+ sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult = 1.280     
+ sky130_fd_pr__nfet_01v8__ajunction_mult = 1.2169e+0
+ sky130_fd_pr__nfet_01v8__pjunction_mult = 1.2474e+0
+ sky130_fd_pr__pfet_01v8__ajunction_mult = 0.90161
+ sky130_fd_pr__pfet_01v8__pjunction_mult = 0.90587
