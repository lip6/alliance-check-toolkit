* MacroLib

* PNP_05v5_W3u40L3u40
.subckt PNP_05v5_W3u40L3u40 collector base emitter
Xpnp collector base emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
.ends PNP_05v5_W3u40L3u40
