* test bench for functional verification of flop with reset
.LIB 'mm0355v.l' TT
* The extracted netlist
.INCLUDE 'check/sff1r_x4.spi'

.PARAM VVDD = 3.3
.PARAM VNRST = 0

XFF clk d nrst q vdd vss sff1r_x4

VVDD vdd vss DC VVDD
VVSS vss 0 DC 0

VD d vss PWL(0 0 2NS 0 2.1NS VVDD)
VCLK clk vss PWL(0 0 1.0NS 0 1.1NS VVDD 2NS VVDD 2.1NS 0 3.0NS 0 3.1NS VVDD 4.5NS VVDD 4.6NS 0)
VNRST nrst vss PWL(0 VVDD 5.0NS VVDD 5.1NS 0)
CQ q vss 10f

.TRAN 0.01NS 6NS
.SAVE ALL
.END
