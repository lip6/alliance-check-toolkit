* Spice description of no4_x1
* Spice driver version -82268389
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:03

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt no4_x1 7 8 6 5 9 1 10 
* NET 1 = vdd
* NET 5 = i3
* NET 6 = i2
* NET 7 = i0
* NET 8 = i1
* NET 9 = nq
* NET 10 = vss
Mtr_00008 3 6 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 2 7 4 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 4 8 9 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 1 5 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00004 10 5 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00003 9 6 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 10 7 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 9 8 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C10 1 10 1.66309e-15
C6 5 10 2.05116e-15
C5 6 10 1.74315e-15
C4 7 10 1.75626e-15
C3 8 10 1.74659e-15
C2 9 10 2.65925e-15
C1 10 10 2.20691e-15
.ends no4_x1

