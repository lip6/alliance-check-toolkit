-- no model for buf_x2
