* using
* Coriolis Structural SPICE Driver
* Generated on Oct 21, 2022, 15:40
* Cell/Subckt "sarlogic_r".
* 
* top_r_hitas_eldo.cir bench SARlogic
* 

*****************

.TEMP 25
.GLOBAL VDD VSS
Vsupply vdd 0  DC 1.8
Vground vss 0  DC 0

******************
* circuit model
* include standard cells
.INCLUDE /users/soft/techno/techno/pdkmaster/views/tsmc_c018/FlexLib/spice/FlexLib.spi
.INCLUDE /users/soft/techno/techno/pdkmaster/views/tsmc_c018/FlexLib/spice/tiepoly_x0.spi

* include circuit netlist
*.subckt sarlogic_r 0 1 2 4 5 30 31 32 33 34 35 36 37 49 58 59 60 61 62 63 64 65 66 67
.INCLUDE sarlogic_r_netlist.spi

* Interface
* INTERF vss
* INTERF vdd
* INTERF soc
* INTERF se
* INTERF rst
* INTERF res[7]
* INTERF res[6]
* INTERF res[5]
* INTERF res[4]
* INTERF res[3]
* INTERF res[2]
* INTERF res[1]
* INTERF res[0]
* INTERF eoc
* INTERF dac_control[7]
* INTERF dac_control[6]
* INTERF dac_control[5]
* INTERF dac_control[4]
* INTERF dac_control[3]
* INTERF dac_control[2]
* INTERF dac_control[1]
* INTERF dac_control[0]
* INTERF cmp
* INTERF clk

* NET     0 = vss
* NET     1 = vdd
* NET     2 = soc
* NET     4 = se
* NET     5 = rst
* NET    30 = res[7]
* NET    31 = res[6]
* NET    32 = res[5]
* NET    33 = res[4]
* NET    34 = res[3]
* NET    35 = res[2]
* NET    36 = res[1]
* NET    37 = res[0]
* NET    49 = eoc
* NET    58 = dac_control[7]
* NET    59 = dac_control[6]
* NET    60 = dac_control[5]
* NET    61 = dac_control[4]
* NET    62 = dac_control[3]
* NET    63 = dac_control[2]
* NET    64 = dac_control[1]
* NET    65 = dac_control[0]
* NET    66 = cmp
* NET    67 = clk
.end
