*.include /users/cao/aoudrhiri/coriolis-2.x/src/alliance-check-toolkit/pdkmaster/C4M.Sky130/libs.ref/StdCellLib/spice/StdCellLib.spi
* Spice driver version -182784229
* Date ( dd/mm/yyyy hh:mm:ss ):  2/07/2024 at 13:54:53

* INTERF adrs[0] adrs[1] adrs[2] adrs[3] adrs[4] adrs[5] adrs[6] adrs[7] 
* INTERF adrs[8] adrs[9] adrs[10] adrs[11] adrs[12] adrs[13] adrs[14] 
* INTERF adrs[15] data[0] data[1] data[2] data[3] data[4] data[5] data[6] 
* INTERF data[7] datao[0] datao[1] datao[2] datao[3] datao[4] datao[5] 
* INTERF datao[6] datao[7] debug[0] debug[1] debug[2] debug[3] debug[4] 
* INTERF debug[5] debug[6] debug[7] debug[8] debug[9] debug[10] debug[11] 
* INTERF debug[12] debug[13] debug[14] debug[15] irq m_clock nmi p_reset rd 
* INTERF rdy start sync vdd vss wt 


.subckt m65_cts_r_ext 6571 6376 6522 6165 5936 5501 5039 5268 3946 3709 3547 3546 3382 3376 3379 3560 6727 6265 5902 5372 5262 5243 4308 5272 6491 6024 5585 5168 5325 4465 4021 3614 6906 6893 6885 6874 6850 6820 6740 6591 6807 6905 6665 5670 5524 5026 4918 4914 6243 m_clock 6261 6976 3655 6440 6728 5907 vdd vss 4720 
* NET 29 = subckt_1623_sff1_x4.sff_m
* NET 30 = subckt_1623_sff1_x4.ckr
* NET 34 = subckt_1624_sff1_x4.sff_m
* NET 35 = subckt_1624_sff1_x4.ckr
* NET 39 = subckt_1632_sff1_x4.sff_m
* NET 40 = subckt_1632_sff1_x4.ckr
* NET 43 = subckt_1634_sff1_x4.sff_m
* NET 45 = subckt_1634_sff1_x4.ckr
* NET 48 = subckt_1619_sff1_x4.sff_m
* NET 50 = subckt_1619_sff1_x4.ckr
* NET 54 = subckt_1627_sff1_x4.sff_m
* NET 55 = subckt_1627_sff1_x4.ckr
* NET 69 = abc_8311_new_n932
* NET 81 = abc_8311_new_n950
* NET 86 = abc_8311_new_n945
* NET 95 = subckt_1623_sff1_x4.sff_s
* NET 99 = subckt_1623_sff1_x4.nckr
* NET 101 = subckt_1624_sff1_x4.sff_s
* NET 105 = subckt_1624_sff1_x4.nckr
* NET 107 = subckt_1632_sff1_x4.sff_s
* NET 111 = subckt_1632_sff1_x4.nckr
* NET 115 = subckt_1634_sff1_x4.sff_s
* NET 120 = subckt_1634_sff1_x4.nckr
* NET 121 = subckt_1619_sff1_x4.sff_s
* NET 124 = subckt_1619_sff1_x4.nckr
* NET 126 = subckt_1627_sff1_x4.sff_s
* NET 131 = subckt_1627_sff1_x4.nckr
* NET 133 = abc_8311_new_n605
* NET 138 = abc_8311_new_n604
* NET 191 = abc_8311_new_n1094
* NET 196 = abc_8311_new_n1081
* NET 200 = abc_8311_new_n1093
* NET 209 = abc_8311_new_n948
* NET 210 = abc_8311_new_n942
* NET 212 = abc_8311_new_n946
* NET 214 = abc_8311_new_n944
* NET 216 = abc_8311_new_n940
* NET 222 = abc_8311_auto_rtlil_cc_2693_muxgate_8270
* NET 225 = abc_8311_auto_rtlil_cc_2693_muxgate_8272
* NET 228 = subckt_1631_sff1_x4.sff_s
* NET 231 = subckt_1631_sff1_x4.sff_m
* NET 233 = subckt_1631_sff1_x4.ckr
* NET 235 = subckt_1631_sff1_x4.nckr
* NET 237 = abc_8311_auto_rtlil_cc_2693_muxgate_8286
* NET 239 = abc_8311_auto_rtlil_cc_2693_muxgate_8288
* NET 243 = abc_8311_auto_rtlil_cc_2693_muxgate_8292
* NET 246 = subckt_1626_sff1_x4.sff_s
* NET 249 = subckt_1626_sff1_x4.sff_m
* NET 251 = subckt_1626_sff1_x4.ckr
* NET 254 = subckt_1626_sff1_x4.nckr
* NET 255 = abc_8311_auto_rtlil_cc_2693_muxgate_8262
* NET 258 = abc_8311_auto_rtlil_cc_2693_muxgate_8278
* NET 261 = abc_8311_new_n1726
* NET 263 = abc_8311_new_n618
* NET 264 = abc_8311_new_n620
* NET 265 = abc_8311_new_n622
* NET 301 = abc_8311_new_n1090
* NET 302 = abc_8311_new_n1088
* NET 305 = abc_8311_new_n1089
* NET 307 = abc_8311_new_n1073
* NET 310 = abc_8311_new_n1015
* NET 312 = abc_8311_new_n1087
* NET 314 = abc_8311_new_n1074
* NET 319 = abc_8311_new_n941
* NET 320 = abc_8311_new_n947
* NET 322 = abc_8311_new_n1092
* NET 323 = abc_8311_new_n1016
* NET 328 = abc_8311_new_n1011
* NET 332 = abc_8311_new_n1009
* NET 335 = abc_8311_new_n1008
* NET 342 = subckt_1622_sff1_x4.sff_s
* NET 345 = subckt_1622_sff1_x4.sff_m
* NET 348 = subckt_1622_sff1_x4.ckr
* NET 349 = subckt_1622_sff1_x4.nckr
* NET 350 = abc_8311_auto_rtlil_cc_2693_muxgate_8268
* NET 355 = subckt_1630_sff1_x4.sff_s
* NET 358 = subckt_1630_sff1_x4.sff_m
* NET 362 = subckt_1630_sff1_x4.ckr
* NET 363 = subckt_1630_sff1_x4.nckr
* NET 364 = abc_8311_auto_rtlil_cc_2693_muxgate_8284
* NET 369 = subckt_1633_sff1_x4.sff_s
* NET 372 = subckt_1633_sff1_x4.sff_m
* NET 376 = subckt_1633_sff1_x4.nckr
* NET 377 = subckt_1633_sff1_x4.ckr
* NET 379 = subckt_1625_sff1_x4.sff_s
* NET 382 = subckt_1625_sff1_x4.sff_m
* NET 384 = subckt_1625_sff1_x4.ckr
* NET 386 = subckt_1625_sff1_x4.nckr
* NET 387 = abc_8311_auto_rtlil_cc_2693_muxgate_8276
* NET 392 = ry[7]
* NET 395 = abc_8311_new_n623
* NET 399 = abc_8311_new_n1725
* NET 402 = abc_8311_new_n631
* NET 405 = abc_8311_new_n603
* NET 461 = abc_8311_new_n1097
* NET 466 = abc_8311_new_n1125
* NET 470 = abc_8311_new_n1077
* NET 473 = abc_8311_new_n1078
* NET 476 = abc_8311_new_n1069
* NET 477 = abc_8311_new_n1014
* NET 478 = abc_8311_new_n1012
* NET 480 = abc_8311_new_n1017
* NET 482 = abc_8311_new_n1013
* NET 486 = abc_8311_new_n949
* NET 488 = abc_8311_new_n1007
* NET 489 = abc_8311_new_n1010
* NET 491 = abc_8311_new_n943
* NET 493 = abc_8311_new_n939
* NET 494 = abc_8311_new_n1006
* NET 500 = ry[4]
* NET 502 = ry[3]
* NET 504 = ry[5]
* NET 509 = subckt_1607_sff1_x4.sff_s
* NET 513 = subckt_1607_sff1_x4.sff_m
* NET 514 = subckt_1607_sff1_x4.ckr
* NET 516 = subckt_1607_sff1_x4.nckr
* NET 517 = abc_8311_auto_rtlil_cc_2693_muxgate_8274
* NET 522 = rx[7]
* NET 525 = rx[0]
* NET 527 = ry[0]
* NET 530 = subckt_1603_sff1_x4.sff_s
* NET 534 = subckt_1603_sff1_x4.sff_m
* NET 536 = subckt_1603_sff1_x4.ckr
* NET 537 = subckt_1603_sff1_x4.nckr
* NET 569 = abc_8311_new_n1086
* NET 571 = abc_8311_new_n1095
* NET 573 = abc_8311_new_n1126
* NET 576 = abc_8311_new_n1096
* NET 579 = abc_8311_new_n1098
* NET 581 = abc_8311_new_n1084
* NET 586 = abc_8311_new_n1083
* NET 588 = abc_8311_new_n1079
* NET 589 = abc_8311_new_n1076
* NET 591 = abc_8311_new_n1082
* NET 592 = abc_8311_new_n1080
* NET 596 = abc_8311_new_n1042
* NET 598 = abc_8311_new_n1068
* NET 603 = abc_8311_new_n1070
* NET 607 = abc_8311_new_n1071
* NET 611 = abc_8311_new_n1072
* NET 615 = abc_8311_new_n938
* NET 619 = abc_8311_new_n1067
* NET 624 = abc_8311_new_n897
* NET 625 = abc_8311_new_n895
* NET 629 = abc_8311_new_n957
* NET 633 = rx[4]
* NET 636 = rx[5]
* NET 640 = abc_8311_new_n1066
* NET 641 = abc_8311_new_n959
* NET 643 = subckt_1608_sff1_x4.sff_s
* NET 646 = subckt_1608_sff1_x4.sff_m
* NET 650 = subckt_1608_sff1_x4.ckr
* NET 651 = subckt_1608_sff1_x4.nckr
* NET 652 = abc_8311_auto_rtlil_cc_2693_muxgate_8208
* NET 657 = abc_8311_auto_rtlil_cc_2693_muxgate_8206
* NET 661 = abc_8311_auto_rtlil_cc_2693_muxgate_8290
* NET 663 = ry[6]
* NET 669 = subckt_1628_sff1_x4.sff_s
* NET 673 = subckt_1628_sff1_x4.sff_m
* NET 675 = subckt_1628_sff1_x4.ckr
* NET 676 = subckt_1628_sff1_x4.nckr
* NET 677 = abc_8311_auto_rtlil_cc_2693_muxgate_8198
* NET 682 = abc_8311_new_n607
* NET 686 = abc_8311_new_n498
* NET 690 = abc_8311_new_n1181
* NET 766 = abc_8311_new_n1018
* NET 769 = abc_8311_new_n833
* NET 770 = abc_8311_new_n812
* NET 772 = abc_8311_new_n931
* NET 774 = abc_8311_new_n1041
* NET 776 = abc_8311_new_n1128
* NET 779 = abc_8311_new_n1005
* NET 784 = abc_8311_new_n1004
* NET 787 = abc_8311_new_n937
* NET 791 = abc_8311_new_n982
* NET 793 = abc_8311_new_n983
* NET 794 = abc_8311_new_n935
* NET 801 = abc_8311_new_n914
* NET 803 = subckt_1629_sff1_x4.sff_s
* NET 806 = subckt_1629_sff1_x4.sff_m
* NET 809 = subckt_1629_sff1_x4.ckr
* NET 810 = abc_8311_auto_rtlil_cc_2693_muxgate_8282
* NET 811 = subckt_1629_sff1_x4.nckr
* NET 817 = subckt_1621_sff1_x4.sff_s
* NET 821 = subckt_1621_sff1_x4.sff_m
* NET 823 = subckt_1621_sff1_x4.ckr
* NET 824 = subckt_1621_sff1_x4.nckr
* NET 825 = rx[6]
* NET 828 = abc_8311_auto_rtlil_cc_2693_muxgate_8280
* NET 829 = ry[1]
* NET 830 = abc_8311_new_n1727
* NET 836 = subckt_1610_sff1_x4.sff_s
* NET 840 = subckt_1610_sff1_x4.sff_m
* NET 842 = subckt_1610_sff1_x4.ckr
* NET 843 = subckt_1610_sff1_x4.nckr
* NET 844 = abc_8311_new_n611
* NET 845 = abc_8311_new_n472
* NET 849 = abc_8311_new_n477
* NET 851 = abc_8311_new_n500
* NET 857 = abc_8311_new_n471
* NET 859 = abc_8311_new_n610
* NET 860 = abc_8311_new_n499
* NET 863 = abc_8311_new_n245
* NET 870 = abc_8311_new_n1127
* NET 911 = abc_8311_new_n742
* NET 914 = abc_8311_new_n989
* NET 917 = abc_8311_new_n1117
* NET 918 = abc_8311_new_n894
* NET 919 = abc_8311_new_n896
* NET 923 = subckt_1620_sff1_x4.sff_m
* NET 924 = subckt_1620_sff1_x4.ckr
* NET 925 = subckt_1620_sff1_x4.nckr
* NET 933 = abc_8311_new_n813
* NET 936 = abc_8311_new_n831
* NET 938 = abc_8311_new_n810
* NET 941 = abc_8311_new_n811
* NET 943 = abc_8311_new_n805
* NET 946 = abc_8311_new_n600
* NET 947 = abc_8311_new_n806
* NET 953 = abc_8311_new_n1091
* NET 961 = abc_8311_new_n1019
* NET 965 = abc_8311_new_n953
* NET 968 = abc_8311_new_n986
* NET 973 = abc_8311_new_n984
* NET 975 = abc_8311_new_n1104
* NET 980 = abc_8311_new_n1105
* NET 981 = abc_8311_new_n1002
* NET 982 = abc_8311_new_n976
* NET 986 = abc_8311_new_n626
* NET 987 = abc_8311_new_n617
* NET 988 = ry[2]
* NET 990 = abc_8311_auto_rtlil_cc_2693_muxgate_8266
* NET 998 = subckt_1620_sff1_x4.sff_s
* NET 1001 = abc_8311_auto_rtlil_cc_2693_muxgate_8264
* NET 1002 = rx[1]
* NET 1004 = abc_8311_new_n1716
* NET 1007 = abc_8311_auto_rtlil_cc_2693_muxgate_8212
* NET 1029 = abc_8311_new_n473
* NET 1031 = abc_8311_new_n488
* NET 1033 = abc_8311_new_n382
* NET 1035 = abc_8311_new_n1715
* NET 1038 = abc_8311_new_n608
* NET 1039 = abc_8311_new_n632
* NET 1138 = subckt_1575_sff1_x4.sff_s
* NET 1142 = subckt_1575_sff1_x4.sff_m
* NET 1143 = subckt_1575_sff1_x4.ckr
* NET 1145 = subckt_1575_sff1_x4.nckr
* NET 1146 = abc_8311_new_n809
* NET 1151 = abc_8311_new_n885
* NET 1156 = abc_8311_new_n801
* NET 1158 = abc_8311_new_n770
* NET 1163 = abc_8311_new_n1153
* NET 1165 = abc_8311_new_n1100
* NET 1169 = abc_8311_new_n737
* NET 1171 = abc_8311_new_n740
* NET 1172 = abc_8311_new_n985
* NET 1175 = abc_8311_new_n936
* NET 1176 = abc_8311_new_n915
* NET 1177 = abc_8311_new_n954
* NET 1178 = abc_8311_new_n981
* NET 1182 = rx[3]
* NET 1186 = abc_8311_new_n977
* NET 1188 = abc_8311_new_n956
* NET 1189 = abc_8311_new_n958
* NET 1190 = abc_8311_new_n606
* NET 1191 = rx[2]
* NET 1194 = abc_8311_new_n612
* NET 1196 = abc_8311_new_n1145
* NET 1198 = subckt_1609_sff1_x4.sff_s
* NET 1200 = subckt_1609_sff1_x4.sff_m
* NET 1203 = abc_8311_auto_rtlil_cc_2693_muxgate_8210
* NET 1204 = subckt_1609_sff1_x4.ckr
* NET 1206 = subckt_1609_sff1_x4.nckr
* NET 1208 = abc_8311_new_n1173
* NET 1209 = abc_8311_new_n739
* NET 1210 = abc_8311_new_n581
* NET 1212 = abc_8311_new_n1193
* NET 1214 = abc_8311_new_n580
* NET 1215 = abc_8311_new_n578
* NET 1218 = abc_8311_new_n389
* NET 1221 = abc_8311_new_n570
* NET 1223 = abc_8311_new_n385
* NET 1224 = abc_8311_new_n567
* NET 1229 = abc_8311_new_n1186
* NET 1231 = abc_8311_new_n384
* NET 1232 = abc_8311_new_n569
* NET 1233 = abc_8311_new_n496
* NET 1234 = abc_8311_new_n534
* NET 1235 = abc_8311_new_n1185
* NET 1236 = abc_8311_new_n568
* NET 1239 = abc_8311_new_n301
* NET 1280 = abc_8311_new_n820
* NET 1287 = abc_8311_new_n818
* NET 1289 = abc_8311_new_n804
* NET 1292 = abc_8311_new_n815
* NET 1298 = abc_8311_new_n769
* NET 1300 = abc_8311_new_n1101
* NET 1304 = abc_8311_new_n1129
* NET 1306 = abc_8311_new_n1154
* NET 1309 = abc_8311_new_n1156
* NET 1312 = abc_8311_new_n1085
* NET 1313 = abc_8311_new_n1099
* NET 1315 = spare_buffer_18.q
* NET 1317 = abc_8311_new_n1050
* NET 1320 = abc_8311_new_n768
* NET 1322 = abc_8311_new_n583
* NET 1323 = abc_8311_new_n1003
* NET 1326 = abc_8311_new_n1112
* NET 1328 = abc_8311_new_n1106
* NET 1329 = abc_8311_new_n1107
* NET 1330 = abc_8311_new_n1113
* NET 1332 = abc_8311_new_n980
* NET 1333 = abc_8311_new_n978
* NET 1338 = abc_8311_new_n1109
* NET 1339 = abc_8311_new_n1111
* NET 1340 = abc_8311_new_n975
* NET 1343 = abc_8311_new_n1110
* NET 1345 = abc_8311_new_n1029
* NET 1346 = abc_8311_new_n1028
* NET 1353 = abc_8311_new_n680
* NET 1356 = abc_8311_new_n682
* NET 1360 = abc_8311_new_n503
* NET 1365 = abc_8311_new_n571
* NET 1367 = abc_8311_new_n736
* NET 1370 = spare_buffer_14.q
* NET 1372 = abc_8311_new_n1745
* NET 1379 = abc_8311_new_n566
* NET 1380 = abc_8311_new_n1184
* NET 1381 = abc_8311_new_n1694
* NET 1385 = abc_8311_new_n497
* NET 1389 = abc_8311_new_n609
* NET 1390 = abc_8311_new_n493
* NET 1394 = abc_8311_new_n369
* NET 1395 = abc_8311_new_n494
* NET 1478 = abc_8311_new_n819
* NET 1479 = abc_8311_new_n830
* NET 1480 = abc_8311_new_n816
* NET 1482 = abc_8311_new_n796
* NET 1483 = abc_8311_new_n802
* NET 1484 = abc_8311_new_n817
* NET 1485 = abc_8311_new_n807
* NET 1488 = abc_8311_new_n795
* NET 1490 = abc_8311_new_n803
* NET 1491 = abc_8311_new_n814
* NET 1492 = abc_8311_new_n799
* NET 1498 = abc_8311_new_n794
* NET 1501 = abc_8311_new_n748
* NET 1505 = abc_8311_new_n1026
* NET 1508 = abc_8311_new_n1027
* NET 1510 = spare_buffer_17.q
* NET 1513 = abc_8311_new_n1049
* NET 1517 = abc_8311_new_n1114
* NET 1518 = abc_8311_new_n1103
* NET 1521 = abc_8311_new_n917
* NET 1524 = abc_8311_new_n955
* NET 1527 = abc_8311_new_n916
* NET 1530 = abc_8311_new_n979
* NET 1533 = abc_8311_new_n1108
* NET 1534 = abc_8311_new_n913
* NET 1541 = abc_8311_new_n668
* NET 1542 = abc_8311_new_n666
* NET 1544 = subckt_1606_sff1_x4.sff_s
* NET 1548 = subckt_1606_sff1_x4.sff_m
* NET 1549 = abc_8311_auto_rtlil_cc_2693_muxgate_8204
* NET 1551 = subckt_1606_sff1_x4.ckr
* NET 1552 = subckt_1606_sff1_x4.nckr
* NET 1553 = abc_8311_new_n476
* NET 1558 = abc_8311_new_n1194
* NET 1559 = abc_8311_new_n629
* NET 1560 = abc_8311_new_n449
* NET 1562 = abc_8311_new_n483
* NET 1563 = abc_8311_new_n478
* NET 1564 = abc_8311_new_n735
* NET 1565 = abc_8311_new_n1760
* NET 1569 = spare_buffer_13.q
* NET 1572 = abc_8311_new_n1182
* NET 1575 = abc_8311_new_n1766
* NET 1576 = abc_8311_new_n257
* NET 1578 = abc_8311_new_n639
* NET 1579 = abc_8311_new_n317
* NET 1580 = abc_8311_new_n318
* NET 1582 = abc_8311_new_n383
* NET 1583 = abc_8311_new_n621
* NET 1587 = abc_8311_new_n596
* NET 1588 = abc_8311_new_n327
* NET 1620 = abc_8311_new_n829
* NET 1627 = abc_8311_new_n808
* NET 1632 = abc_8311_new_n822
* NET 1635 = abc_8311_new_n800
* NET 1640 = abc_8311_new_n601
* NET 1641 = abc_8311_new_n792
* NET 1645 = abc_8311_new_n793
* NET 1647 = abc_8311_new_n749
* NET 1649 = abc_8311_new_n951
* NET 1652 = abc_8311_new_n1040
* NET 1655 = abc_8311_new_n1075
* NET 1661 = abc_8311_new_n1192
* NET 1662 = abc_8311_new_n1241
* NET 1667 = abc_8311_new_n747
* NET 1669 = abc_8311_new_n918
* NET 1670 = abc_8311_new_n892
* NET 1676 = abc_8311_new_n767
* NET 1679 = abc_8311_new_n751
* NET 1682 = abc_8311_new_n766
* NET 1687 = abc_8311_new_n764
* NET 1688 = abc_8311_new_n753
* NET 1694 = abc_8311_new_n1131
* NET 1695 = abc_8311_new_n1242
* NET 1699 = abc_8311_new_n1136
* NET 1700 = abc_8311_new_n1138
* NET 1703 = abc_8311_new_n688
* NET 1704 = abc_8311_new_n1137
* NET 1706 = abc_8311_new_n1166
* NET 1708 = abc_8311_new_n1168
* NET 1716 = abc_8311_new_n1167
* NET 1722 = abc_8311_new_n1191
* NET 1724 = abc_8311_new_n1195
* NET 1727 = abc_8311_new_n564
* NET 1728 = abc_8311_new_n1196
* NET 1730 = abc_8311_new_n577
* NET 1732 = abc_8311_new_n559
* NET 1735 = abc_8311_new_n1761
* NET 1737 = abc_8311_new_n597
* NET 1740 = abc_8311_new_n598
* NET 1744 = abc_8311_new_n484
* NET 1745 = abc_8311_new_n560
* NET 1746 = abc_8311_new_n390
* NET 1749 = abc_8311_new_n310
* NET 1757 = abc_8311_new_n625
* NET 1758 = abc_8311_new_n591
* NET 1760 = abc_8311_new_n387
* NET 1778 = abc_8311_new_n533
* NET 1779 = abc_8311_new_n300
* NET 1875 = abc_8311_new_n828
* NET 1876 = abc_8311_new_n738
* NET 1877 = abc_8311_new_n832
* NET 1880 = abc_8311_new_n825
* NET 1882 = abc_8311_new_n797
* NET 1883 = abc_8311_new_n824
* NET 1884 = abc_8311_new_n798
* NET 1885 = abc_8311_new_n722
* NET 1886 = abc_8311_new_n821
* NET 1888 = abc_8311_new_n719
* NET 1891 = abc_8311_new_n730
* NET 1893 = abc_8311_new_n777
* NET 1900 = abc_8311_new_n510
* NET 1904 = abc_8311_new_n563
* NET 1905 = abc_8311_new_n574
* NET 1911 = abc_8311_new_n746
* NET 1913 = abc_8311_new_n890
* NET 1914 = abc_8311_new_n889
* NET 1918 = abc_8311_new_n765
* NET 1919 = abc_8311_new_n750
* NET 1925 = abc_8311_new_n1142
* NET 1929 = abc_8311_new_n1064
* NET 1931 = abc_8311_new_n780
* NET 1933 = abc_8311_new_n779
* NET 1944 = abc_8311_new_n1243
* NET 1945 = abc_8311_new_n1162
* NET 1946 = abc_8311_new_n562
* NET 1947 = abc_8311_new_n1762
* NET 1950 = abc_8311_new_n1765
* NET 1953 = abc_8311_new_n328
* NET 1956 = subckt_1641_sff1r_x4.sff_s
* NET 1959 = abc_8311_auto_rtlil_cc_2693_muxgate_8310
* NET 1960 = subckt_1641_sff1r_x4.sff_m
* NET 1963 = subckt_1641_sff1r_x4.ckr
* NET 1964 = subckt_1641_sff1r_x4.nckr
* NET 1965 = abc_8311_new_n531
* NET 1967 = abc_8311_new_n594
* NET 1968 = abc_8311_new_n687
* NET 1971 = abc_8311_new_n686
* NET 1972 = abc_8311_new_n685
* NET 1973 = abc_8311_new_n684
* NET 1975 = abc_8311_new_n595
* NET 1979 = abc_8311_new_n324
* NET 1982 = abc_8311_new_n592
* NET 1985 = abc_8311_new_n320
* NET 1986 = abc_8311_new_n319
* NET 1988 = abc_8311_new_n391
* NET 1989 = abc_8311_new_n388
* NET 1990 = abc_8311_new_n386
* NET 1991 = abc_8311_new_n326
* NET 1992 = abc_8311_new_n380
* NET 2044 = abc_8311_new_n891
* NET 2045 = abc_8311_new_n919
* NET 2046 = abc_8311_new_n893
* NET 2048 = abc_8311_new_n923
* NET 2050 = abc_8311_new_n1163
* NET 2051 = abc_8311_new_n1164
* NET 2052 = abc_8311_new_n1169
* NET 2057 = abc_8311_new_n1763
* NET 2058 = abc_8311_new_n546
* NET 2065 = subckt_1635_sff1_x4.sff_m
* NET 2067 = subckt_1635_sff1_x4.ckr
* NET 2068 = subckt_1635_sff1_x4.nckr
* NET 2070 = abc_8311_new_n630
* NET 2074 = abc_8311_new_n1188
* NET 2080 = abc_8311_new_n858
* NET 2086 = abc_8311_new_n558
* NET 2088 = abc_8311_new_n727
* NET 2092 = abc_8311_new_n731
* NET 2095 = abc_8311_new_n720
* NET 2097 = abc_8311_new_n778
* NET 2102 = abc_8311_new_n721
* NET 2106 = abc_8311_new_n557
* NET 2107 = abc_8311_new_n662
* NET 2109 = abc_8311_new_n697
* NET 2111 = abc_8311_new_n588
* NET 2116 = abc_8311_new_n696
* NET 2117 = abc_8311_new_n695
* NET 2122 = abc_8311_new_n694
* NET 2124 = abc_8311_new_n448
* NET 2125 = abc_8311_new_n323
* NET 2128 = abc_8311_new_n1133
* NET 2129 = abc_8311_new_n1140
* NET 2135 = abc_8311_new_n1048
* NET 2136 = abc_8311_new_n1065
* NET 2138 = abc_8311_new_n1157
* NET 2139 = abc_8311_new_n1170
* NET 2142 = abc_8311_new_n1051
* NET 2144 = abc_8311_new_n1132
* NET 2146 = abc_8311_new_n1165
* NET 2154 = abc_8311_new_n1161
* NET 2155 = abc_8311_new_n576
* NET 2156 = abc_8311_new_n1197
* NET 2157 = abc_8311_new_n613
* NET 2161 = abc_8311_new_n556
* NET 2165 = abc_8311_new_n627
* NET 2167 = subckt_1635_sff1_x4.sff_s
* NET 2170 = abc_8311_new_n481
* NET 2173 = abc_8311_new_n482
* NET 2174 = abc_8311_new_n644
* NET 2180 = abc_8311_new_n329
* NET 2182 = abc_8311_new_n304
* NET 2183 = abc_8311_new_n309
* NET 2184 = abc_8311_new_n645
* NET 2188 = abc_8311_new_n619
* NET 2193 = abc_8311_new_n322
* NET 2194 = abc_8311_new_n377
* NET 2195 = abc_8311_new_n370
* NET 2196 = abc_8311_new_n393
* NET 2198 = abc_8311_new_n325
* NET 2202 = abc_8311_new_n395
* NET 2207 = abc_8311_new_n330
* NET 2208 = abc_8311_new_n313
* NET 2286 = abc_8311_new_n859
* NET 2291 = abc_8311_new_n732
* NET 2292 = abc_8311_new_n728
* NET 2298 = abc_8311_new_n725
* NET 2299 = abc_8311_new_n717
* NET 2301 = abc_8311_new_n711
* NET 2303 = abc_8311_new_n723
* NET 2304 = abc_8311_new_n726
* NET 2306 = abc_8311_new_n718
* NET 2307 = abc_8311_new_n724
* NET 2308 = abc_8311_new_n729
* NET 2314 = abc_8311_new_n602
* NET 2319 = abc_8311_new_n575
* NET 2320 = abc_8311_new_n659
* NET 2323 = abc_8311_new_n692
* NET 2325 = abc_8311_new_n1240
* NET 2326 = abc_8311_new_n743
* NET 2329 = abc_8311_new_n665
* NET 2331 = abc_8311_new_n663
* NET 2333 = abc_8311_new_n744
* NET 2336 = abc_8311_new_n870
* NET 2340 = abc_8311_new_n1134
* NET 2342 = abc_8311_new_n869
* NET 2344 = abc_8311_new_n1139
* NET 2345 = abc_8311_new_n1135
* NET 2346 = abc_8311_new_n1141
* NET 2347 = abc_8311_new_n752
* NET 2349 = abc_8311_new_n689
* NET 2350 = abc_8311_new_n683
* NET 2352 = abc_8311_new_n367
* NET 2353 = abc_8311_new_n690
* NET 2355 = abc_8311_new_n664
* NET 2356 = abc_8311_new_n1025
* NET 2360 = abc_8311_new_n1764
* NET 2361 = abc_8311_new_n1159
* NET 2364 = subckt_1605_sff1_x4.sff_s
* NET 2367 = subckt_1605_sff1_x4.sff_m
* NET 2369 = subckt_1605_sff1_x4.ckr
* NET 2371 = abc_8311_new_n508
* NET 2372 = subckt_1605_sff1_x4.nckr
* NET 2375 = abc_8311_new_n545
* NET 2379 = abc_8311_new_n572
* NET 2381 = abc_8311_new_n565
* NET 2382 = abc_8311_new_n573
* NET 2384 = abc_8311_new_n505
* NET 2386 = abc_8311_new_n701
* NET 2387 = abc_8311_new_n459
* NET 2389 = abc_8311_new_n479
* NET 2392 = abc_8311_new_n480
* NET 2394 = abc_8311_new_n475
* NET 2396 = abc_8311_new_n1183
* NET 2399 = abc_8311_new_n638
* NET 2400 = abc_8311_new_n495
* NET 2404 = abc_8311_new_n451
* NET 2406 = abc_8311_new_n298
* NET 2407 = abc_8311_new_n312
* NET 2408 = abc_8311_new_n399
* NET 2409 = abc_8311_new_n321
* NET 2411 = abc_8311_new_n381
* NET 2412 = abc_8311_new_n302
* NET 2415 = abc_8311_new_n373
* NET 2418 = abc_8311_new_n343
* NET 2461 = subckt_1571_sff1_x4.sff_s
* NET 2465 = subckt_1571_sff1_x4.sff_m
* NET 2468 = subckt_1571_sff1_x4.ckr
* NET 2469 = subckt_1571_sff1_x4.nckr
* NET 2479 = abc_8311_new_n657
* NET 2483 = abc_8311_new_n660
* NET 2485 = abc_8311_new_n658
* NET 2487 = abc_8311_new_n656
* NET 2489 = abc_8311_new_n716
* NET 2492 = abc_8311_new_n715
* NET 2495 = abc_8311_new_n771
* NET 2498 = abc_8311_new_n599
* NET 2499 = abc_8311_new_n661
* NET 2501 = abc_8311_new_n506
* NET 2506 = abc_8311_new_n561
* NET 2507 = abc_8311_new_n888
* NET 2508 = abc_8311_new_n920
* NET 2511 = abc_8311_new_n714
* NET 2512 = abc_8311_new_n678
* NET 2513 = abc_8311_new_n840
* NET 2514 = abc_8311_new_n693
* NET 2517 = abc_8311_new_n691
* NET 2518 = abc_8311_new_n842
* NET 2519 = abc_8311_new_n844
* NET 2520 = abc_8311_new_n655
* NET 2521 = abc_8311_new_n681
* NET 2522 = abc_8311_new_n843
* NET 2525 = abc_8311_new_n865
* NET 2526 = abc_8311_new_n866
* NET 2530 = abc_8311_new_n1045
* NET 2532 = abc_8311_new_n1047
* NET 2534 = abc_8311_new_n679
* NET 2535 = abc_8311_new_n791
* NET 2536 = abc_8311_new_n845
* NET 2537 = abc_8311_new_n912
* NET 2542 = abc_8311_new_n781
* NET 2544 = abc_8311_new_n1063
* NET 2545 = abc_8311_new_n1053
* NET 2546 = abc_8311_new_n1052
* NET 2550 = abc_8311_new_n667
* NET 2551 = abc_8311_new_n1160
* NET 2553 = abc_8311_new_n1039
* NET 2560 = abc_8311_auto_rtlil_cc_2693_muxgate_8202
* NET 2562 = abc_8311_new_n616
* NET 2567 = subckt_1604_sff1_x4.sff_s
* NET 2570 = subckt_1604_sff1_x4.sff_m
* NET 2573 = subckt_1604_sff1_x4.ckr
* NET 2574 = subckt_1604_sff1_x4.nckr
* NET 2578 = abc_8311_new_n641
* NET 2582 = abc_8311_auto_rtlil_cc_2693_muxgate_8294
* NET 2583 = tc
* NET 2587 = abc_8311_new_n457
* NET 2591 = subckt_1538_sff1r_x4.sff_s
* NET 2594 = subckt_1538_sff1r_x4.sff_m
* NET 2598 = subckt_1538_sff1r_x4.nckr
* NET 2599 = subckt_1538_sff1r_x4.ckr
* NET 2600 = abc_8311_new_n1198
* NET 2601 = abc_8311_auto_rtlil_cc_2693_muxgate_8068
* NET 2603 = abc_8311_new_n1189
* NET 2604 = abc_8311_new_n1187
* NET 2607 = abc_8311_new_n633
* NET 2610 = abc_8311_new_n635
* NET 2615 = abc_8311_new_n368
* NET 2622 = abc_8311_new_n394
* NET 2623 = abc_8311_new_n392
* NET 2625 = abc_8311_new_n374
* NET 2628 = abc_8311_new_n375
* NET 2629 = abc_8311_new_n308
* NET 2632 = abc_8311_new_n306
* NET 2705 = subckt_1574_sff1_x4.sff_s
* NET 2708 = subckt_1574_sff1_x4.sff_m
* NET 2710 = subckt_1574_sff1_x4.ckr
* NET 2712 = abc_8311_new_n883
* NET 2713 = subckt_1574_sff1_x4.nckr
* NET 2716 = abc_8311_new_n861
* NET 2717 = abc_8311_new_n860
* NET 2720 = abc_8311_new_n836
* NET 2723 = abc_8311_new_n734
* NET 2727 = abc_8311_new_n741
* NET 2728 = abc_8311_new_n834
* NET 2730 = abc_8311_new_n590
* NET 2733 = abc_8311_new_n587
* NET 2734 = abc_8311_new_n589
* NET 2736 = abc_8311_new_n776
* NET 2737 = abc_8311_new_n775
* NET 2739 = abc_8311_new_n712
* NET 2740 = abc_8311_new_n586
* NET 2741 = abc_8311_new_n875
* NET 2742 = abc_8311_new_n1239
* NET 2744 = abc_8311_new_n1238
* NET 2746 = abc_8311_new_n288
* NET 2747 = abc_8311_new_n1001
* NET 2749 = abc_8311_new_n868
* NET 2750 = abc_8311_new_n871
* NET 2752 = abc_8311_new_n867
* NET 2755 = abc_8311_new_n1046
* NET 2758 = abc_8311_new_n1044
* NET 2763 = abc_8311_new_n1144
* NET 2766 = abc_8311_new_n1038
* NET 2770 = abc_8311_new_n974
* NET 2773 = abc_8311_new_n642
* NET 2775 = abc_8311_new_n1236
* NET 2778 = abc_8311_new_n1037
* NET 2779 = abc_8311_new_n1237
* NET 2782 = abc_8311_new_n504
* NET 2787 = abc_8311_new_n474
* NET 2788 = abc_8311_new_n491
* NET 2790 = abc_8311_new_n507
* NET 2792 = abc_8311_auto_rtlil_cc_2693_muxgate_8200
* NET 2793 = abc_8311_new_n850
* NET 2797 = abc_8311_new_n1695
* NET 2799 = abc_8311_new_n247
* NET 2801 = abc_8311_new_n1768
* NET 2803 = abc_8311_new_n1767
* NET 2807 = abc_8311_new_n409
* NET 2809 = subckt_1639_sff1r_x4.sff_s
* NET 2812 = subckt_1639_sff1r_x4.sff_m
* NET 2815 = subckt_1639_sff1r_x4.ckr
* NET 2816 = subckt_1639_sff1r_x4.nckr
* NET 2817 = abc_8311_new_n1204
* NET 2820 = abc_8311_new_n1203
* NET 2823 = abc_8311_new_n1190
* NET 2824 = abc_8311_new_n1753
* NET 2826 = abc_8311_auto_rtlil_cc_2693_muxgate_8306
* NET 2827 = abc_8311_new_n1312
* NET 2830 = abc_8311_new_n452
* NET 2833 = abc_8311_new_n376
* NET 2834 = abc_8311_new_n371
* NET 2836 = abc_8311_new_n397
* NET 2837 = abc_8311_new_n378
* NET 2842 = subckt_1579_sff1_x4.sff_s
* NET 2846 = subckt_1579_sff1_x4.sff_m
* NET 2849 = subckt_1579_sff1_x4.nckr
* NET 2850 = subckt_1579_sff1_x4.ckr
* NET 2851 = abc_8311_auto_rtlil_cc_2693_muxgate_8150
* NET 2852 = op[0]
* NET 2895 = abc_8311_new_n827
* NET 2896 = abc_8311_new_n826
* NET 2897 = abc_8311_new_n823
* NET 2901 = subckt_1576_sff1_x4.sff_s
* NET 2903 = subckt_1576_sff1_x4.sff_m
* NET 2907 = subckt_1576_sff1_x4.ckr
* NET 2908 = subckt_1576_sff1_x4.nckr
* NET 2909 = abc_8311_new_n884
* NET 2913 = abc_8311_new_n886
* NET 2915 = abc_8311_new_n837
* NET 2919 = abc_8311_new_n862
* NET 2921 = abc_8311_new_n733
* NET 2924 = abc_8311_new_n835
* NET 2928 = subckt_1578_sff1_x4.sff_s
* NET 2931 = subckt_1578_sff1_x4.sff_m
* NET 2933 = subckt_1578_sff1_x4.ckr
* NET 2935 = subckt_1578_sff1_x4.nckr
* NET 2936 = abc_8311_new_n772
* NET 2938 = abc_8311_new_n864
* NET 2940 = abc_8311_new_n872
* NET 2944 = abc_8311_new_n584
* NET 2946 = abc_8311_new_n1023
* NET 2950 = abc_8311_new_n1020
* NET 2951 = abc_8311_new_n1024
* NET 2952 = abc_8311_new_n1021
* NET 2953 = abc_8311_new_n1022
* NET 2958 = subckt_1617_sff1r_x4.sff_s
* NET 2961 = abc_8311_auto_rtlil_cc_2693_muxgate_8254
* NET 2962 = subckt_1617_sff1r_x4.sff_m
* NET 2965 = subckt_1617_sff1r_x4.ckr
* NET 2966 = subckt_1617_sff1r_x4.nckr
* NET 2970 = subckt_1618_sff1r_x4.sff_s
* NET 2973 = subckt_1618_sff1r_x4.sff_m
* NET 2976 = subckt_1618_sff1r_x4.ckr
* NET 2977 = abc_8311_auto_rtlil_cc_2693_muxgate_8260
* NET 2978 = subckt_1618_sff1r_x4.nckr
* NET 2979 = abc_8311_auto_ff_cc_704_flip_bits_8255
* NET 2981 = abc_8311_new_n1172
* NET 2986 = abc_8311_new_n677
* NET 2987 = abc_8311_new_n669
* NET 2990 = abc_8311_new_n1030
* NET 2993 = abc_8311_new_n1036
* NET 2996 = abc_8311_new_n1031
* NET 2997 = abc_8311_new_n1247
* NET 2998 = abc_8311_new_n1248
* NET 2999 = abc_8311_new_n1155
* NET 3003 = abc_8311_new_n637
* NET 3004 = abc_8311_new_n654
* NET 3006 = abc_8311_new_n544
* NET 3010 = abc_8311_new_n542
* NET 3015 = abc_8311_new_n541
* NET 3021 = abc_8311_new_n463
* NET 3023 = abc_8311_new_n461
* NET 3029 = subckt_1638_sff1r_x4.sff_s
* NET 3032 = subckt_1638_sff1r_x4.sff_m
* NET 3035 = subckt_1638_sff1r_x4.nckr
* NET 3036 = subckt_1638_sff1r_x4.ckr
* NET 3037 = abc_8311_new_n256
* NET 3039 = abc_8311_auto_rtlil_cc_2693_muxgate_8304
* NET 3040 = abc_8311_new_n258
* NET 3042 = abc_8311_new_n1746
* NET 3044 = abc_8311_new_n1750
* NET 3046 = abc_8311_new_n1201
* NET 3049 = abc_8311_new_n437
* NET 3051 = abc_8311_new_n634
* NET 3060 = abc_8311_new_n303
* NET 3062 = abc_8311_new_n314
* NET 3069 = subckt_1583_sff1_x4.sff_s
* NET 3073 = subckt_1583_sff1_x4.sff_m
* NET 3075 = subckt_1583_sff1_x4.ckr
* NET 3076 = subckt_1583_sff1_x4.nckr
* NET 3144 = subckt_1572_sff1_x4.sff_s
* NET 3147 = subckt_1572_sff1_x4.sff_m
* NET 3150 = subckt_1572_sff1_x4.ckr
* NET 3151 = subckt_1572_sff1_x4.nckr
* NET 3152 = abc_8311_auto_rtlil_cc_2693_muxgate_8144
* NET 3153 = subckt_1577_sff1_x4.sff_s
* NET 3158 = subckt_1577_sff1_x4.sff_m
* NET 3160 = m_clock_root_tr_0
* NET 3161 = subckt_1577_sff1_x4.ckr
* NET 3162 = subckt_1577_sff1_x4.nckr
* NET 3163 = abc_8311_auto_rtlil_cc_2693_muxgate_8146
* NET 3165 = abc_8311_new_n1607
* NET 3167 = abc_8311_new_n774
* NET 3172 = abc_8311_new_n773
* NET 3174 = abc_8311_new_n839
* NET 3178 = abc_8311_new_n988
* NET 3182 = abc_8311_new_n847
* NET 3183 = abc_8311_new_n841
* NET 3184 = abc_8311_new_n846
* NET 3186 = abc_8311_new_n470
* NET 3187 = abc_8311_new_n933
* NET 3188 = abc_8311_new_n934
* NET 3190 = abc_8311_auto_ff_cc_704_flip_bits_8249
* NET 3191 = abc_8311_new_n1000
* NET 3193 = abc_8311_new_n910
* NET 3195 = abc_8311_new_n972
* NET 3197 = abc_8311_new_n898
* NET 3199 = abc_8311_new_n615
* NET 3201 = abc_8311_new_n960
* NET 3202 = abc_8311_new_n909
* NET 3204 = abc_8311_new_n900
* NET 3208 = abc_8311_new_n790
* NET 3210 = abc_8311_new_n911
* NET 3212 = abc_8311_new_n899
* NET 3217 = abc_8311_new_n554
* NET 3218 = abc_8311_new_n513
* NET 3221 = abc_8311_new_n1704
* NET 3225 = abc_8311_new_n1705
* NET 3226 = abc_8311_new_n468
* NET 3227 = abc_8311_new_n540
* NET 3229 = abc_8311_new_n535
* NET 3231 = abc_8311_new_n539
* NET 3233 = abc_8311_new_n538
* NET 3234 = abc_8311_new_n530
* NET 3236 = abc_8311_new_n1202
* NET 3238 = abc_8311_new_n1752
* NET 3242 = abc_8311_new_n1200
* NET 3245 = abc_8311_new_n1749
* NET 3246 = abc_8311_new_n1748
* NET 3248 = abc_8311_new_n1747
* NET 3252 = subckt_1580_sff1_x4.sff_s
* NET 3257 = subckt_1580_sff1_x4.sff_m
* NET 3259 = m_clock_root_tl_0
* NET 3260 = subckt_1580_sff1_x4.nckr
* NET 3261 = subckt_1580_sff1_x4.ckr
* NET 3262 = abc_8311_auto_rtlil_cc_2693_muxgate_8158
* NET 3263 = op[4]
* NET 3312 = subckt_1573_sff1_x4.sff_m
* NET 3313 = subckt_1573_sff1_x4.ckr
* NET 3314 = subckt_1573_sff1_x4.nckr
* NET 3315 = abc_8311_auto_rtlil_cc_2693_muxgate_8142
* NET 3317 = abc_8311_new_n1595
* NET 3318 = abc_8311_auto_rtlil_cc_2693_muxgate_8140
* NET 3326 = subckt_1614_sff1r_x4.sff_m
* NET 3328 = subckt_1614_sff1r_x4.ckr
* NET 3329 = subckt_1614_sff1r_x4.nckr
* NET 3335 = subckt_1615_sff1r_x4.sff_m
* NET 3337 = abc_8311_auto_rtlil_cc_2693_muxgate_8242
* NET 3339 = subckt_1615_sff1r_x4.ckr
* NET 3340 = subckt_1615_sff1r_x4.nckr
* NET 3347 = subckt_1616_sff1r_x4.sff_m
* NET 3349 = subckt_1616_sff1r_x4.nckr
* NET 3350 = subckt_1616_sff1r_x4.ckr
* NET 3360 = subckt_1640_sff1r_x4.sff_m
* NET 3363 = subckt_1640_sff1r_x4.nckr
* NET 3364 = subckt_1640_sff1r_x4.ckr
* NET 3369 = abc_8311_new_n406
* NET 3371 = abc_8311_new_n366
* NET 3373 = subckt_1573_sff1_x4.sff_s
* NET 3376 = adrs[13]
* NET 3379 = adrs[14]
* NET 3382 = adrs[12]
* NET 3385 = subckt_1614_sff1r_x4.sff_s
* NET 3388 = subckt_1615_sff1r_x4.sff_s
* NET 3391 = abc_8311_new_n745
* NET 3395 = abc_8311_auto_ff_cc_704_flip_bits_8237
* NET 3396 = subckt_1616_sff1r_x4.sff_s
* NET 3397 = abc_8311_auto_rtlil_cc_2693_muxgate_8248
* NET 3401 = abc_8311_new_n1116
* NET 3403 = abc_8311_auto_ff_cc_704_flip_bits_8243
* NET 3404 = abc_8311_new_n961
* NET 3408 = abc_8311_new_n973
* NET 3413 = abc_8311_new_n636
* NET 3414 = abc_8311_new_n628
* NET 3416 = abc_8311_new_n782
* NET m_clock = m_clock
* NET 3421 = ra[2]
* NET 3423 = ra[7]
* NET 3424 = abc_8311_new_n469
* NET 3429 = abc_8311_new_n653
* NET 3430 = abc_8311_new_n647
* NET 3434 = ra[0]
* NET 3438 = abc_8311_new_n526
* NET 3442 = abc_8311_new_n331
* NET 3445 = subckt_1640_sff1r_x4.sff_s
* NET 3449 = abc_8311_new_n398
* NET 3451 = abc_8311_new_n408
* NET 3452 = abc_8311_new_n364
* NET 3453 = abc_8311_new_n413
* NET 3455 = abc_8311_new_n400
* NET 3456 = abc_8311_new_n379
* NET 3457 = abc_8311_new_n396
* NET 3458 = abc_8311_new_n410
* NET 3459 = abc_8311_auto_rtlil_cc_2693_muxgate_8152
* NET 3460 = op[1]
* NET 3546 = adrs[11]
* NET 3547 = adrs[10]
* NET 3548 = abc_8311_auto_rtlil_cc_2693_muxgate_8138
* NET 3549 = abc_8311_new_n1599
* NET 3550 = abc_8311_new_n1597
* NET 3552 = abc_8311_new_n1611
* NET 3553 = abc_8311_new_n1609
* NET 3555 = abc_8311_new_n1617
* NET 3556 = abc_8311_new_n1615
* NET 3558 = abc_8311_new_n1589
* NET 3560 = adrs[15]
* NET 3561 = abc_8311_new_n1601
* NET 3563 = abc_8311_auto_rtlil_cc_2693_muxgate_8148
* NET 3565 = abc_8311_auto_rtlil_cc_2693_muxgate_8236
* NET 3566 = abc_8311_new_n922
* NET 3570 = abc_8311_new_n849
* NET 3572 = abc_8311_new_n585
* NET 3573 = abc_8311_auto_ff_cc_704_flip_bits_8231
* NET 3576 = subckt_1611_sff1r_x4.sff_s
* NET 3579 = subckt_1611_sff1r_x4.sff_m
* NET 3582 = subckt_1611_sff1r_x4.ckr
* NET 3583 = subckt_1611_sff1r_x4.nckr
* NET 3586 = abc_8311_new_n1043
* NET 3589 = abc_8311_new_n962
* NET 3591 = abc_8311_new_n971
* NET 3592 = abc_8311_new_n968
* NET 3593 = abc_8311_new_n763
* NET 3595 = abc_8311_new_n754
* NET 3596 = abc_8311_new_n908
* NET 3598 = abc_8311_new_n907
* NET 3600 = abc_8311_new_n1054
* NET 3602 = abc_8311_new_n1062
* NET 3604 = ra[3]
* NET 3606 = abc_8311_new_n906
* NET 3607 = ra[4]
* NET 3608 = abc_8311_new_n901
* NET 3610 = abc_8311_new_n676
* NET 3613 = abc_8311_new_n1174
* NET 3614 = datao[7]
* NET 3616 = abc_8311_new_n671
* NET 3617 = abc_8311_new_n490
* NET 3618 = abc_8311_new_n516
* NET 3621 = abc_8311_new_n1636
* NET 3622 = abc_8311_new_n1270
* NET 3624 = abc_8311_new_n403
* NET 3625 = abc_8311_new_n462
* NET 3629 = abc_8311_new_n525
* NET 3631 = abc_8311_new_n614
* NET 3632 = abc_8311_new_n315
* NET 3634 = abc_8311_new_n254
* NET 3636 = abc_8311_new_n537
* NET 3637 = abc_8311_new_n431
* NET 3639 = abc_8311_new_n455
* NET 3640 = abc_8311_auto_rtlil_cc_2693_muxgate_8308
* NET 3641 = abc_8311_new_n269
* NET 3645 = abc_8311_new_n1758
* NET 3648 = abc_8311_new_n1757
* NET 3649 = abc_8311_new_n453
* NET 3652 = abc_8311_new_n414
* NET 3653 = abc_8311_new_n415
* NET 3654 = abc_8311_new_n454
* NET 3655 = rd
* NET 3658 = abc_8311_new_n342
* NET 3660 = abc_8311_new_n624
* NET 3662 = abc_8311_new_n1756
* NET 3663 = abc_8311_new_n1755
* NET 3664 = abc_8311_new_n246
* NET 3709 = adrs[9]
* NET 3712 = abc_8311_auto_rtlil_cc_2693_muxgate_8136
* NET 3714 = abc_8311_new_n1593
* NET 3715 = abc_8311_new_n1591
* NET 3717 = abc_8311_new_n1605
* NET 3720 = abc_8311_new_n1603
* NET 3725 = abc_8311_new_n1583
* NET 3727 = abc_8311_new_n1623
* NET 3728 = abc_8311_new_n1621
* NET 3734 = abc_8311_new_n1604
* NET 3736 = abc_8311_new_n1613
* NET 3737 = abc_8311_new_n582
* NET 3738 = abc_8311_new_n509
* NET 3740 = abc_8311_new_n555
* NET 3741 = abc_8311_new_n713
* NET 3746 = subckt_1612_sff1r_x4.sff_s
* NET 3748 = subckt_1612_sff1r_x4.sff_m
* NET 3750 = abc_8311_auto_rtlil_cc_2693_muxgate_8224
* NET 3753 = subckt_1612_sff1r_x4.ckr
* NET 3754 = subckt_1612_sff1r_x4.nckr
* NET 3757 = abc_8311_new_n1610
* NET 3758 = abc_8311_auto_rtlil_cc_2693_muxgate_8218
* NET 3759 = abc_8311_auto_ff_cc_704_flip_bits_8213
* NET 3761 = abc_8311_new_n700
* NET 3766 = abc_8311_new_n1616
* NET 3769 = subckt_1589_sff1_x4.sff_s
* NET 3772 = subckt_1589_sff1_x4.sff_m
* NET 3774 = subckt_1589_sff1_x4.ckr
* NET 3776 = abc_8311_new_n970
* NET 3777 = subckt_1589_sff1_x4.nckr
* NET 3781 = abc_8311_new_n969
* NET 3783 = abc_8311_new_n1061
* NET 3788 = abc_8311_new_n963
* NET 3789 = abc_8311_new_n643
* NET 3790 = ra[6]
* NET 3792 = abc_8311_new_n646
* NET 3793 = abc_8311_new_n579
* NET 3795 = abc_8311_new_n1056
* NET 3796 = ra[5]
* NET 3797 = abc_8311_new_n1578
* NET 3798 = abc_8311_new_n512
* NET 3800 = abc_8311_new_n282
* NET 3802 = ra[1]
* NET 3805 = abc_8311_new_n407
* NET 3813 = abc_8311_new_n502
* NET 3814 = abc_8311_new_n511
* NET 3816 = abc_8311_new_n517
* NET 3818 = abc_8311_new_n365
* NET 3819 = abc_8311_new_n402
* NET 3821 = abc_8311_new_n467
* NET 3827 = abc_8311_new_n520
* NET 3831 = abc_8311_new_n523
* NET 3836 = abc_8311_new_n250
* NET 3849 = abc_8311_new_n299
* NET 3853 = abc_8311_new_n354
* NET 3856 = abc_8311_new_n1319
* NET 3863 = abc_8311_new_n412
* NET 3866 = abc_8311_new_n305
* NET 3868 = subckt_1586_sff1_x4.sff_s
* NET 3870 = subckt_1586_sff1_x4.sff_m
* NET 3873 = subckt_1586_sff1_x4.ckr
* NET 3875 = subckt_1586_sff1_x4.nckr
* NET 3946 = adrs[8]
* NET 3947 = abc_8311_new_n1579
* NET 3948 = abc_8311_new_n1571
* NET 3949 = abc_8311_auto_rtlil_cc_2693_muxgate_8134
* NET 3950 = abc_8311_new_n1587
* NET 3951 = abc_8311_new_n1585
* NET 3953 = abc_8311_new_n1608
* NET 3957 = abc_8311_new_n1614
* NET 3962 = abc_8311_new_n1425
* NET 3964 = abc_8311_new_n1598
* NET 3967 = abc_8311_new_n1592
* NET 3969 = abc_8311_new_n1570
* NET 3971 = abc_8311_new_n1619
* NET 3972 = abc_8311_auto_ff_cc_704_flip_bits_8219
* NET 3975 = abc_8311_new_n874
* NET 3976 = abc_8311_new_n1706
* NET 3979 = abc_8311_auto_ff_cc_704_flip_bits_8225
* NET 3981 = subckt_1613_sff1r_x4.sff_s
* NET 3985 = subckt_1613_sff1r_x4.sff_m
* NET 3986 = abc_8311_auto_rtlil_cc_2693_muxgate_8230
* NET 3987 = subckt_1613_sff1r_x4.ckr
* NET 3989 = subckt_1613_sff1r_x4.nckr
* NET 3991 = abc_8311_new_n1574
* NET 3993 = subckt_1593_sff1_x4.sff_s
* NET 3997 = subckt_1593_sff1_x4.sff_m
* NET 4000 = subckt_1593_sff1_x4.ckr
* NET 4001 = subckt_1593_sff1_x4.nckr
* NET 4002 = abc_8311_auto_rtlil_cc_2693_muxgate_8178
* NET 4008 = abc_8311_new_n762
* NET 4009 = abc_8311_new_n761
* NET 4010 = abc_8311_new_n755
* NET 4013 = abc_8311_new_n1577
* NET 4014 = abc_8311_new_n789
* NET 4015 = abc_8311_new_n784
* NET 4016 = abc_8311_new_n783
* NET 4018 = abc_8311_new_n670
* NET 4020 = abc_8311_new_n1146
* NET 4021 = datao[6]
* NET 4024 = abc_8311_new_n279
* NET 4028 = abc_8311_new_n268
* NET 4032 = abc_8311_new_n285
* NET 4038 = abc_8311_new_n528
* NET 4042 = abc_8311_new_n1445
* NET 4043 = abc_8311_new_n265
* NET 4048 = abc_8311_new_n543
* NET 4051 = abc_8311_new_n492
* NET 4052 = abc_8311_new_n1254
* NET 4053 = abc_8311_new_n435
* NET 4059 = abc_8311_new_n263
* NET 4062 = abc_8311_new_n466
* NET 4066 = abc_8311_new_n1635
* NET 4068 = abc_8311_new_n532
* NET 4071 = abc_8311_new_n251
* NET 4072 = abc_8311_new_n1633
* NET 4075 = abc_8311_new_n1740
* NET 4079 = abc_8311_new_n416
* NET 4080 = abc_8311_new_n450
* NET 4082 = abc_8311_new_n430
* NET 4083 = abc_8311_new_n1199
* NET 4086 = abc_8311_new_n446
* NET 4087 = abc_8311_new_n340
* NET 4088 = abc_8311_new_n372
* NET 4089 = abc_8311_new_n341
* NET 4091 = abc_8311_new_n411
* NET 4093 = abc_8311_auto_rtlil_cc_2693_muxgate_8164
* NET 4094 = op[7]
* NET 4150 = abc_8311_new_n1576
* NET 4151 = abc_8311_new_n1581
* NET 4153 = abc_8311_new_n1580
* NET 4157 = abc_8311_new_n1414
* NET 4160 = abc_8311_new_n1428
* NET 4163 = abc_8311_new_n280
* NET 4171 = abc_8311_new_n1586
* NET 4175 = abc_8311_new_n1422
* NET 4176 = abc_8311_new_n289
* NET 4181 = abc_8311_new_n1622
* NET 4183 = subckt_1590_sff1_x4.sff_s
* NET 4186 = subckt_1590_sff1_x4.sff_m
* NET 4189 = subckt_1590_sff1_x4.ckr
* NET 4190 = subckt_1590_sff1_x4.nckr
* NET 4191 = abc_8311_auto_rtlil_cc_2693_muxgate_8172
* NET 4200 = abc_8311_auto_rtlil_cc_2693_muxgate_8170
* NET 4205 = abc_8311_new_n236
* NET 4212 = abc_8311_new_n527
* NET 4213 = abc_8311_new_n640
* NET 4215 = abc_8311_new_n1055
* NET 4217 = abc_8311_new_n1573
* NET 4220 = abc_8311_new_n464
* NET 4224 = abc_8311_new_n272
* NET 4226 = abc_8311_new_n1179
* NET 4228 = abc_8311_new_n1178
* NET 4233 = abc_8311_new_n456
* NET 4235 = fn
* NET 4238 = abc_8311_new_n1175
* NET 4239 = fd
* NET 4241 = fv
* NET 4250 = abc_8311_new_n518
* NET 4253 = abc_8311_new_n521
* NET 4254 = abc_8311_new_n432
* NET 4257 = abc_8311_new_n1634
* NET 4258 = abc_8311_new_n529
* NET 4261 = abc_8311_new_n252
* NET 4265 = abc_8311_new_n417
* NET 4273 = abc_8311_new_n1320
* NET 4275 = abc_8311_new_n249
* NET 4276 = abc_8311_new_n339
* NET 4280 = abc_8311_new_n255
* NET 4281 = abc_8311_new_n349
* NET 4282 = abc_8311_new_n260
* NET 4285 = abc_8311_new_n418
* NET 4286 = abc_8311_new_n307
* NET 4287 = abc_8311_new_n355
* NET 4290 = subckt_1581_sff1_x4.sff_s
* NET 4293 = subckt_1581_sff1_x4.sff_m
* NET 4297 = subckt_1581_sff1_x4.ckr
* NET 4298 = subckt_1581_sff1_x4.nckr
* NET 4299 = op[2]
* NET 4300 = abc_8311_auto_rtlil_cc_2693_muxgate_8154
* NET 4308 = data[6]
* NET 4386 = subckt_1560_sff1_x4.sff_s
* NET 4390 = subckt_1560_sff1_x4.sff_m
* NET 4392 = subckt_1560_sff1_x4.ckr
* NET 4393 = subckt_1560_sff1_x4.nckr
* NET 4394 = abc_8311_new_n1411
* NET 4395 = abc_8311_auto_rtlil_cc_2693_muxgate_8112
* NET 4396 = abc_8311_new_n1420
* NET 4397 = abc_8311_new_n1419
* NET 4399 = abc_8311_new_n1620
* NET 4401 = abc_8311_new_n1435
* NET 4405 = subckt_1561_sff1_x4.sff_s
* NET 4409 = subckt_1561_sff1_x4.sff_m
* NET 4410 = abc_8311_auto_rtlil_cc_2693_muxgate_8114
* NET 4412 = subckt_1561_sff1_x4.ckr
* NET 4413 = subckt_1561_sff1_x4.nckr
* NET 4414 = abc_8311_new_n1431
* NET 4418 = subckt_1570_sff1_x4.sff_s
* NET 4421 = subckt_1570_sff1_x4.sff_m
* NET 4424 = subckt_1570_sff1_x4.ckr
* NET 4425 = subckt_1570_sff1_x4.nckr
* NET 4429 = subckt_1592_sff1_x4.sff_s
* NET 4432 = subckt_1592_sff1_x4.sff_m
* NET 4434 = abc_8311_auto_rtlil_cc_2693_muxgate_8176
* NET 4435 = subckt_1592_sff1_x4.ckr
* NET 4437 = subckt_1592_sff1_x4.nckr
* NET 4438 = abc_8311_new_n235
* NET 4441 = abc_8311_new_n233
* NET 4444 = abc_8311_new_n1565
* NET 4447 = abc_8311_new_n1564
* NET 4452 = abc_8311_new_n1575
* NET 4453 = abc_8311_new_n1446
* NET 4455 = abc_8311_new_n1271
* NET 4456 = abc_8311_new_n549
* NET 4460 = abc_8311_new_n1449
* NET 4461 = abc_8311_new_n1151
* NET 4462 = abc_8311_new_n1147
* NET 4463 = abc_8311_new_n1150
* NET 4465 = datao[5]
* NET 4466 = abc_8311_new_n995
* NET 4469 = abc_8311_new_n1121
* NET 4470 = abc_8311_new_n704
* NET 4471 = abc_8311_new_n1255
* NET 4472 = abc_8311_new_n465
* NET 4477 = abc_8311_new_n547
* NET 4482 = abc_8311_new_n1246
* NET 4483 = abc_8311_new_n1251
* NET 4485 = abc_8311_new_n460
* NET 4488 = abc_8311_new_n1265
* NET 4489 = abc_8311_new_n1259
* NET 4491 = abc_8311_new_n426
* NET 4492 = abc_8311_new_n522
* NET 4496 = abc_8311_new_n1264
* NET 4497 = abc_8311_new_n1260
* NET 4499 = abc_8311_new_n1263
* NET 4501 = abc_8311_new_n248
* NET 4502 = abc_8311_new_n1324
* NET 4503 = abc_8311_new_n1321
* NET 4505 = abc_8311_new_n429
* NET 4506 = abc_8311_new_n444
* NET 4507 = abc_8311_new_n433
* NET 4509 = abc_8311_new_n311
* NET 4510 = abc_8311_new_n1323
* NET 4512 = abc_8311_new_n1742
* NET 4515 = abc_8311_new_n425
* NET 4517 = abc_8311_new_n420
* NET 4518 = abc_8311_new_n1739
* NET 4520 = abc_8311_new_n1741
* NET 4521 = abc_8311_new_n1743
* NET 4523 = abc_8311_new_n316
* NET 4524 = op[6]
* NET 4525 = subckt_1585_sff1_x4.sff_s
* NET 4530 = subckt_1585_sff1_x4.sff_m
* NET 4531 = abc_8311_auto_rtlil_cc_2693_muxgate_8162
* NET 4533 = subckt_1585_sff1_x4.nckr
* NET 4534 = subckt_1585_sff1_x4.ckr
* NET 4572 = abc_8311_new_n519
* NET 4584 = subckt_1562_sff1_x4.sff_m
* NET 4585 = subckt_1562_sff1_x4.ckr
* NET 4586 = subckt_1562_sff1_x4.nckr
* NET 4587 = abc_8311_new_n1433
* NET 4589 = abc_8311_auto_rtlil_cc_2693_muxgate_8132
* NET 4591 = abc_8311_new_n1542
* NET 4604 = abc_8311_new_n1060
* NET 4608 = abc_8311_new_n1035
* NET 4609 = abc_8311_new_n1122
* NET 4610 = abc_8311_new_n1123
* NET 4611 = abc_8311_new_n1272
* NET 4612 = abc_8311_new_n1274
* NET 4613 = abc_8311_new_n348
* NET 4616 = abc_8311_new_n353
* NET 4618 = abc_8311_new_n1325
* NET 4622 = abc_8311_new_n424
* NET 4629 = subckt_1637_sff1r_x4.sff_m
* NET 4630 = abc_8311_auto_rtlil_cc_2693_muxgate_8302
* NET 4633 = subckt_1637_sff1r_x4.ckr
* NET 4634 = subckt_1637_sff1r_x4.nckr
* NET 4638 = subckt_1584_sff1_x4.sff_m
* NET 4639 = subckt_1584_sff1_x4.ckr
* NET 4640 = subckt_1584_sff1_x4.nckr
* NET 4643 = abc_8311_new_n1417
* NET 4649 = abc_8311_new_n1415
* NET 4653 = abc_8311_new_n1436
* NET 4658 = abc_8311_new_n1426
* NET 4664 = subckt_1562_sff1_x4.sff_s
* NET 4665 = abc_8311_auto_rtlil_cc_2693_muxgate_8116
* NET 4668 = abc_8311_new_n1423
* NET 4671 = abc_8311_new_n1171
* NET 4672 = abc_8311_new_n1556
* NET 4673 = abc_8311_new_n1158
* NET 4675 = abc_8311_new_n1430
* NET 4676 = abc_8311_new_n290
* NET 4679 = abc_8311_new_n1566
* NET 4682 = abc_8311_new_n1563
* NET 4685 = abc_8311_new_n1536
* NET 4687 = abc_8311_new_n234
* NET 4688 = abc_8311_new_n1551
* NET 4689 = abc_8311_new_n1550
* NET 4692 = abc_8311_new_n1535
* NET 4695 = abc_8311_new_n1058
* NET 4696 = abc_8311_new_n240
* NET 4699 = abc_8311_new_n1033
* NET 4701 = abc_8311_new_n1148
* NET 4703 = abc_8311_new_n1177
* NET 4704 = abc_8311_new_n1120
* NET 4708 = abc_8311_new_n356
* NET 4709 = abc_8311_new_n548
* NET 4715 = abc_8311_new_n514
* NET 4720 = wt
* NET 4722 = abc_8311_new_n362
* NET 4725 = abc_8311_new_n524
* NET 4726 = abc_8311_new_n428
* NET 4731 = abc_8311_new_n357
* NET 4732 = abc_8311_new_n1317
* NET 4733 = abc_8311_new_n427
* NET 4737 = abc_8311_new_n1249
* NET 4744 = abc_8311_new_n423
* NET 4745 = abc_8311_new_n422
* NET 4747 = subckt_1637_sff1r_x4.sff_s
* NET 4748 = op[5]
* NET 4749 = subckt_1584_sff1_x4.sff_s
* NET 4751 = abc_8311_auto_rtlil_cc_2693_muxgate_8160
* NET 4836 = abc_8311_new_n277
* NET 4838 = abc_8311_new_n1590
* NET 4839 = abc_8311_new_n1384
* NET 4843 = abc_8311_new_n1602
* NET 4847 = abc_8311_new_n1416
* NET 4849 = abc_8311_new_n1418
* NET 4850 = abc_8311_new_n1413
* NET 4853 = abc_8311_new_n283
* NET 4854 = abc_8311_new_n1424
* NET 4855 = abc_8311_new_n1427
* NET 4857 = abc_8311_new_n1437
* NET 4859 = abc_8311_new_n1434
* NET 4862 = abc_8311_new_n1441
* NET 4863 = abc_8311_new_n1438
* NET 4865 = abc_8311_new_n1429
* NET 4866 = abc_8311_new_n1439
* NET 4868 = subckt_1569_sff1_x4.sff_s
* NET 4872 = subckt_1569_sff1_x4.sff_m
* NET 4873 = abc_8311_auto_rtlil_cc_2693_muxgate_8130
* NET 4875 = subckt_1569_sff1_x4.ckr
* NET 4876 = abc_8311_new_n1568
* NET 4877 = subckt_1569_sff1_x4.nckr
* NET 4878 = abc_8311_new_n1567
* NET 4880 = abc_8311_new_n1130
* NET 4881 = abc_8311_new_n1143
* NET 4883 = abc_8311_new_n1537
* NET 4886 = abc_8311_new_n1538
* NET 4887 = abc_8311_new_n1552
* NET 4889 = abc_8311_new_n1549
* NET 4892 = abc_8311_new_n1523
* NET 4895 = abc_8311_new_n1505
* NET 4896 = abc_8311_new_n1506
* NET 4897 = abc_8311_new_n237
* NET 4899 = abc_8311_new_n1522
* NET 4903 = abc_8311_new_n1460
* NET 4906 = abc_8311_new_n1461
* NET 4909 = abc_8311_new_n967
* NET 4911 = abc_8311_new_n964
* NET 4914 = debug[15]
* NET 4916 = abc_8311_new_n1032
* NET 4918 = debug[14]
* NET 4919 = abc_8311_new_n1057
* NET 4921 = abc_8311_new_n1034
* NET 4925 = abc_8311_new_n1176
* NET 4927 = abc_8311_new_n927
* NET 4928 = abc_8311_new_n925
* NET 4929 = abc_8311_new_n928
* NET 4935 = fz
* NET 4937 = fc
* NET 4939 = abc_8311_new_n1333
* NET 4941 = abc_8311_new_n344
* NET 4942 = abc_8311_new_n404
* NET 4945 = abc_8311_new_n1327
* NET 4946 = abc_8311_new_n1313
* NET 4947 = abc_8311_new_n332
* NET 4948 = abc_8311_new_n1326
* NET 4952 = abc_8311_new_n1256
* NET 4953 = abc_8311_new_n1257
* NET 4954 = abc_8311_new_n1290
* NET 4955 = subckt_1548_sff1_x4.sff_s
* NET 4960 = subckt_1548_sff1_x4.sff_m
* NET 4961 = abc_8311_auto_rtlil_cc_2693_muxgate_8088
* NET 4963 = subckt_1548_sff1_x4.nckr
* NET 4964 = subckt_1548_sff1_x4.ckr
* NET 5003 = abc_8311_new_n1596
* NET 5004 = abc_8311_new_n1395
* NET 5008 = abc_8311_new_n1392
* NET 5011 = abc_8311_new_n1381
* NET 5014 = abc_8311_new_n1404
* NET 5017 = abc_8311_new_n1403
* NET 5019 = abc_8311_new_n1394
* NET 5022 = abc_8311_new_n1391
* NET 5025 = abc_8311_new_n1412
* NET 5026 = debug[13]
* NET 5029 = abc_8311_new_n1440
* NET 5034 = abc_8311_new_n1554
* NET 5036 = abc_8311_new_n1553
* NET 5039 = adrs[6]
* NET 5041 = abc_8311_new_n1548
* NET 5044 = abc_8311_new_n1102
* NET 5045 = abc_8311_new_n1115
* NET 5048 = subckt_1591_sff1_x4.sff_s
* NET 5050 = subckt_1591_sff1_x4.sff_m
* NET 5054 = m_clock_root_br_2
* NET 5055 = subckt_1591_sff1_x4.ckr
* NET 5056 = subckt_1591_sff1_x4.nckr
* NET 5057 = abc_8311_auto_rtlil_cc_2693_muxgate_8174
* NET 5062 = abc_8311_new_n1493
* NET 5064 = abc_8311_new_n238
* NET 5065 = abc_8311_new_n1492
* NET 5068 = abc_8311_new_n405
* NET 5069 = abc_8311_new_n401
* NET 5075 = subckt_1587_sff1_x4.sff_s
* NET 5077 = subckt_1587_sff1_x4.sff_m
* NET 5081 = subckt_1587_sff1_x4.nckr
* NET 5082 = subckt_1587_sff1_x4.ckr
* NET 5084 = abc_8311_new_n966
* NET 5088 = abc_8311_new_n1118
* NET 5089 = abc_8311_new_n1059
* NET 5094 = abc_8311_new_n1119
* NET 5097 = abc_8311_new_n1149
* NET 5102 = abc_8311_new_n501
* NET 5104 = abc_8311_new_n924
* NET 5106 = abc_8311_new_n929
* NET 5112 = abc_8311_new_n703
* NET 5113 = abc_8311_new_n360
* NET 5115 = abc_8311_new_n1315
* NET 5116 = abc_8311_new_n515
* NET 5121 = spare_buffer_6.q
* NET 5125 = abc_8311_new_n1250
* NET 5127 = abc_8311_new_n1275
* NET 5132 = abc_8311_new_n1277
* NET 5133 = abc_8311_new_n489
* NET 5134 = abc_8311_new_n232
* NET 5140 = abc_8311_new_n1258
* NET 5141 = abc_8311_new_n1279
* NET 5144 = ex_st[4]
* NET 5146 = subckt_1547_sff1_x4.sff_s
* NET 5149 = subckt_1547_sff1_x4.sff_m
* NET 5151 = abc_8311_auto_rtlil_cc_2693_muxgate_8086
* NET 5153 = subckt_1547_sff1_x4.ckr
* NET 5154 = abc_8311_new_n1252
* NET 5155 = subckt_1547_sff1_x4.nckr
* NET 5157 = op[3]
* NET 5159 = subckt_1582_sff1_x4.sff_s
* NET 5162 = subckt_1582_sff1_x4.sff_m
* NET 5164 = abc_8311_auto_rtlil_cc_2693_muxgate_8156
* NET 5166 = subckt_1582_sff1_x4.ckr
* NET 5167 = subckt_1582_sff1_x4.nckr
* NET 5168 = datao[3]
* NET 5243 = data[5]
* NET 5244 = abc_8311_new_n270
* NET 5245 = abc_8311_new_n1382
* NET 5250 = abc_8311_new_n1406
* NET 5254 = abc_8311_new_n1402
* NET 5258 = abc_8311_new_n1409
* NET 5259 = abc_8311_new_n1408
* NET 5261 = abc_8311_new_n1401
* NET 5262 = data[4]
* NET 5263 = abc_8311_new_n1407
* NET 5264 = abc_8311_new_n1361
* NET 5265 = abc_8311_new_n1528
* NET 5268 = adrs[7]
* NET 5269 = abc_8311_new_n1562
* NET 5270 = abc_8311_new_n1692
* NET 5272 = data[7]
* NET 5277 = abc_8311_new_n1509
* NET 5279 = abc_8311_new_n1510
* NET 5283 = subckt_1588_sff1_x4.sff_s
* NET 5286 = subckt_1588_sff1_x4.sff_m
* NET 5290 = subckt_1588_sff1_x4.ckr
* NET 5291 = subckt_1588_sff1_x4.nckr
* NET 5292 = abc_8311_auto_rtlil_cc_2693_muxgate_8168
* NET 5297 = abc_8311_new_n965
* NET 5299 = abc_8311_new_n239
* NET 5300 = abc_8311_new_n550
* NET 5305 = abc_8311_new_n788
* NET 5306 = abc_8311_auto_rtlil_cc_2693_muxgate_8166
* NET 5309 = abc_8311_new_n1637
* NET 5312 = abc_8311_new_n785
* NET 5315 = abc_8311_new_n786
* NET 5319 = abc_8311_new_n877
* NET 5320 = abc_8311_new_n879
* NET 5321 = abc_8311_new_n880
* NET 5322 = abc_8311_new_n878
* NET 5324 = abc_8311_new_n990
* NET 5325 = datao[4]
* NET 5326 = abc_8311_new_n852
* NET 5327 = abc_8311_new_n855
* NET 5329 = abc_8311_new_n1356
* NET 5331 = abc_8311_new_n1262
* NET 5332 = spare_buffer_5.q
* NET 5334 = blockagenet
* NET 5336 = abc_8311_new_n1328
* NET 5337 = abc_8311_new_n1276
* NET 5338 = abc_8311_new_n1329
* NET 5341 = abc_8311_new_n345
* NET 5342 = abc_8311_new_n1266
* NET 5343 = abc_8311_new_n1267
* NET 5345 = abc_8311_new_n443
* NET 5346 = abc_8311_new_n434
* NET 5348 = abc_8311_new_n1282
* NET 5349 = ex_st[0]
* NET 5351 = subckt_1543_sff1_x4.sff_s
* NET 5354 = abc_8311_auto_rtlil_cc_2693_muxgate_8078
* NET 5355 = subckt_1543_sff1_x4.sff_m
* NET 5357 = subckt_1543_sff1_x4.ckr
* NET 5359 = ex_st[5]
* NET 5360 = subckt_1543_sff1_x4.nckr
* NET 5361 = abc_8311_new_n1292
* NET 5363 = ex
* NET 5364 = subckt_1542_sff1r_x4.sff_s
* NET 5367 = subckt_1542_sff1r_x4.sff_m
* NET 5369 = abc_8311_auto_rtlil_cc_2693_muxgate_8076
* NET 5371 = subckt_1542_sff1r_x4.ckr
* NET 5372 = data[3]
* NET 5373 = subckt_1542_sff1r_x4.nckr
* NET 5417 = subckt_1557_sff1_x4.sff_s
* NET 5421 = subckt_1557_sff1_x4.sff_m
* NET 5424 = subckt_1557_sff1_x4.ckr
* NET 5425 = subckt_1557_sff1_x4.nckr
* NET 5426 = subckt_1559_sff1_x4.sff_s
* NET 5430 = subckt_1559_sff1_x4.sff_m
* NET 5431 = abc_8311_auto_rtlil_cc_2693_muxgate_8110
* NET 5434 = subckt_1559_sff1_x4.ckr
* NET 5435 = subckt_1559_sff1_x4.nckr
* NET 5436 = abc_8311_new_n1396
* NET 5440 = abc_8311_new_n1397
* NET 5442 = abc_8311_new_n1390
* NET 5444 = abc_8311_new_n1400
* NET 5448 = subckt_1568_sff1_x4.sff_s
* NET 5452 = subckt_1568_sff1_x4.sff_m
* NET 5453 = abc_8311_auto_rtlil_cc_2693_muxgate_8128
* NET 5454 = subckt_1568_sff1_x4.ckr
* NET 5456 = abc_8311_new_n1561
* NET 5457 = subckt_1568_sff1_x4.nckr
* NET 5465 = subckt_1602_sff1_x4.sff_s
* NET 5468 = abc_8311_auto_rtlil_cc_2693_muxgate_8196
* NET 5469 = subckt_1602_sff1_x4.sff_m
* NET 5471 = subckt_1602_sff1_x4.ckr
* NET 5473 = subckt_1602_sff1_x4.nckr
* NET 5474 = abc_8311_new_n1691
* NET 5478 = abc_8311_new_n1524
* NET 5483 = abc_8311_new_n1521
* NET 5485 = abc_8311_new_n1508
* NET 5489 = abc_8311_new_n1489
* NET 5490 = abc_8311_new_n1494
* NET 5493 = abc_8311_new_n1476
* NET 5496 = abc_8311_new_n1477
* NET 5498 = abc_8311_new_n758
* NET 5500 = abc_8311_new_n760
* NET 5501 = adrs[5]
* NET 5502 = abc_8311_new_n1253
* NET 5504 = abc_8311_new_n1462
* NET 5505 = abc_8311_new_n1459
* NET 5508 = abc_8311_new_n756
* NET 5510 = abc_8311_new_n759
* NET 5518 = abc_8311_new_n926
* NET 5521 = abc_8311_new_n991
* NET 5523 = abc_8311_new_n998
* NET 5524 = debug[12]
* NET 5525 = abc_8311_new_n992
* NET 5528 = abc_8311_new_n881
* NET 5531 = abc_8311_new_n702
* NET 5533 = abc_8311_new_n709
* NET 5534 = abc_8311_new_n705
* NET 5538 = abc_8311_new_n708
* NET 5540 = abc_8311_new_n706
* NET 5544 = abc_8311_new_n487
* NET 5545 = abc_8311_new_n486
* NET 5548 = abc_8311_new_n1273
* NET 5549 = abc_8311_new_n1332
* NET 5551 = abc_8311_new_n1211
* NET 5552 = abc_8311_new_n1314
* NET 5556 = abc_8311_new_n1286
* NET 5557 = abc_8311_new_n1268
* NET 5559 = abc_8311_new_n442
* NET 5561 = abc_8311_new_n1278
* NET 5564 = abc_8311_new_n1284
* NET 5567 = abc_8311_new_n253
* NET 5569 = abc_8311_new_n1288
* NET 5570 = abc_8311_new_n1280
* NET 5573 = abc_8311_new_n1305
* NET 5575 = ex_st[3]
* NET 5577 = subckt_1546_sff1_x4.sff_s
* NET 5580 = abc_8311_auto_rtlil_cc_2693_muxgate_8084
* NET 5581 = subckt_1546_sff1_x4.sff_m
* NET 5583 = subckt_1546_sff1_x4.ckr
* NET 5585 = datao[2]
* NET 5586 = subckt_1546_sff1_x4.nckr
* NET 5666 = abc_8311_new_n1584
* NET 5670 = debug[11]
* NET 5671 = subckt_1558_sff1_x4.sff_s
* NET 5674 = subckt_1558_sff1_x4.sff_m
* NET 5678 = subckt_1558_sff1_x4.ckr
* NET 5679 = subckt_1558_sff1_x4.nckr
* NET 5680 = abc_8311_new_n1398
* NET 5681 = abc_8311_new_n1389
* NET 5682 = abc_8311_auto_rtlil_cc_2693_muxgate_8108
* NET 5684 = subckt_1567_sff1_x4.sff_s
* NET 5689 = subckt_1567_sff1_x4.sff_m
* NET 5691 = subckt_1567_sff1_x4.ckr
* NET 5692 = subckt_1567_sff1_x4.nckr
* NET 5695 = abc_8311_new_n1560
* NET 5699 = abc_8311_new_n1558
* NET 5700 = abc_8311_new_n1529
* NET 5701 = abc_8311_new_n1540
* NET 5702 = abc_8311_new_n1539
* NET 5705 = abc_8311_new_n284
* NET 5708 = abc_8311_new_n1687
* NET 5709 = subckt_1594_sff1_x4.sff_s
* NET 5714 = subckt_1594_sff1_x4.sff_m
* NET 5715 = abc_8311_auto_rtlil_cc_2693_muxgate_8180
* NET 5717 = subckt_1594_sff1_x4.ckr
* NET 5718 = subckt_1594_sff1_x4.nckr
* NET 5721 = abc_8311_new_n921
* NET 5723 = abc_8311_new_n887
* NET 5725 = dl[6]
* NET 5727 = abc_8311_new_n1473
* NET 5728 = abc_8311_new_n1478
* NET 5730 = abc_8311_new_n757
* NET 5733 = abc_8311_new_n902
* NET 5735 = abc_8311_new_n903
* NET 5737 = abc_8311_new_n905
* NET 5738 = abc_8311_new_n904
* NET 5742 = dl[0]
* NET 5745 = abc_8311_new_n675
* NET 5746 = abc_8311_new_n672
* NET 5748 = abc_8311_new_n485
* NET 5749 = abc_8311_new_n436
* NET 5750 = abc_8311_new_n674
* NET 5753 = abc_8311_new_n352
* NET 5755 = abc_8311_new_n707
* NET 5756 = abc_8311_new_n536
* NET 5758 = abc_8311_new_n648
* NET 5759 = abc_8311_new_n652
* NET 5761 = abc_8311_new_n854
* NET 5762 = abc_8311_new_n856
* NET 5763 = abc_8311_new_n649
* NET 5766 = abc_8311_new_n651
* NET 5767 = abc_8311_new_n350
* NET 5770 = abc_8311_new_n1357
* NET 5772 = abc_8311_new_n336
* NET 5773 = ex_st[1]
* NET 5775 = subckt_1544_sff1_x4.sff_s
* NET 5778 = abc_8311_auto_rtlil_cc_2693_muxgate_8080
* NET 5779 = subckt_1544_sff1_x4.sff_m
* NET 5782 = subckt_1544_sff1_x4.ckr
* NET 5783 = subckt_1544_sff1_x4.nckr
* NET 5784 = abc_8311_new_n441
* NET 5787 = abc_8311_new_n440
* NET 5788 = abc_8311_new_n1245
* NET 5789 = abc_8311_new_n1234
* NET 5791 = abc_8311_new_n1235
* NET 5792 = abc_8311_new_n1244
* NET 5794 = subckt_1551_sff1r_x4.sff_s
* NET 5797 = subckt_1551_sff1r_x4.sff_m
* NET 5800 = abc_8311_auto_rtlil_cc_2693_muxgate_8094
* NET 5802 = subckt_1551_sff1r_x4.ckr
* NET 5803 = subckt_1551_sff1r_x4.nckr
* NET 5804 = dl[1]
* NET 5805 = abc_8311_new_n593
* NET 5856 = abc_8311_new_n1378
* NET 5857 = abc_8311_auto_rtlil_cc_2693_muxgate_8106
* NET 5859 = abc_8311_new_n1514
* NET 5861 = abc_8311_auto_rtlil_cc_2693_muxgate_8126
* NET 5862 = abc_8311_new_n1498
* NET 5864 = abc_8311_new_n1677
* NET 5867 = abc_8311_new_n1690
* NET 5877 = abc_8311_new_n445
* NET 5880 = abc_8311_new_n996
* NET 5884 = subckt_1545_sff1_x4.sff_m
* NET 5885 = subckt_1545_sff1_x4.ckr
* NET 5886 = subckt_1545_sff1_x4.nckr
* NET 5889 = abc_8311_new_n421
* NET 5893 = abc_8311_new_n296
* NET 5900 = subckt_1549_sff1r_x4.sff_m
* NET 5902 = data[2]
* NET 5903 = abc_8311_auto_rtlil_cc_2693_muxgate_8090
* NET 5905 = subckt_1549_sff1r_x4.ckr
* NET 5906 = subckt_1549_sff1r_x4.nckr
* NET 5907 = sync
* NET 5910 = abc_8311_new_n266
* NET 5914 = abc_8311_new_n1371
* NET 5915 = abc_8311_new_n1370
* NET 5918 = abc_8311_new_n1387
* NET 5919 = abc_8311_new_n1385
* NET 5925 = abc_8311_new_n1379
* NET 5927 = abc_8311_new_n1316
* NET 5931 = abc_8311_new_n1526
* NET 5932 = abc_8311_new_n1525
* NET 5936 = adrs[4]
* NET 5937 = abc_8311_new_n1515
* NET 5942 = abc_8311_new_n1547
* NET 5943 = abc_8311_new_n1544
* NET 5947 = abc_8311_new_n987
* NET 5948 = abc_8311_new_n1444
* NET 5949 = abc_8311_new_n952
* NET 5951 = abc_8311_new_n1559
* NET 5952 = abc_8311_new_n1557
* NET 5953 = dl[7]
* NET 5954 = abc_8311_new_n1359
* NET 5955 = abc_8311_new_n1689
* NET 5958 = dl[4]
* NET 5959 = dl[5]
* NET 5963 = dl[2]
* NET 5964 = abc_8311_new_n333
* NET 5965 = abc_8311_new_n1447
* NET 5967 = abc_8311_new_n698
* NET 5969 = abc_8311_new_n1448
* NET 5971 = abc_8311_new_n787
* NET 5972 = abc_8311_new_n1464
* NET 5973 = abc_8311_new_n1454
* NET 5975 = abc_8311_new_n1463
* NET 5978 = abc_8311_new_n876
* NET 5983 = abc_8311_new_n997
* NET 5985 = abc_8311_new_n853
* NET 5986 = abc_8311_new_n347
* NET 5987 = abc_8311_new_n553
* NET 5991 = subckt_1545_sff1_x4.sff_s
* NET 5992 = ex_st[2]
* NET 5993 = abc_8311_new_n699
* NET 5994 = abc_8311_auto_rtlil_cc_2693_muxgate_8082
* NET 5998 = abc_8311_new_n650
* NET 5999 = abc_8311_new_n447
* NET 6000 = abc_8311_new_n419
* NET 6004 = abc_8311_new_n1210
* NET 6011 = abc_8311_new_n1322
* NET 6013 = abc_8311_new_n1216
* NET 6014 = abc_8311_new_n1213
* NET 6015 = abc_8311_new_n1737
* NET 6019 = subckt_1549_sff1r_x4.sff_s
* NET 6023 = abc_8311_new_n292
* NET 6024 = datao[1]
* NET 6025 = abc_8311_new_n293
* NET 6112 = abc_8311_new_n275
* NET 6115 = abc_8311_new_n1405
* NET 6116 = abc_8311_new_n1393
* NET 6118 = abc_8311_new_n1572
* NET 6119 = abc_8311_new_n1353
* NET 6123 = abc_8311_new_n1343
* NET 6127 = abc_8311_new_n1380
* NET 6128 = abc_8311_new_n1383
* NET 6129 = abc_8311_new_n1386
* NET 6132 = abc_8311_new_n1331
* NET 6133 = subckt_1566_sff1_x4.sff_s
* NET 6137 = subckt_1566_sff1_x4.sff_m
* NET 6139 = abc_8311_auto_rtlil_cc_2693_muxgate_8124
* NET 6141 = subckt_1566_sff1_x4.ckr
* NET 6142 = subckt_1566_sff1_x4.nckr
* NET 6143 = abc_8311_new_n1482
* NET 6144 = abc_8311_new_n1466
* NET 6145 = subckt_1600_sff1_x4.sff_s
* NET 6148 = subckt_1600_sff1_x4.sff_m
* NET 6150 = abc_8311_auto_rtlil_cc_2693_muxgate_8192
* NET 6153 = subckt_1600_sff1_x4.ckr
* NET 6154 = subckt_1600_sff1_x4.nckr
* NET 6156 = subckt_1601_sff1_x4.sff_s
* NET 6158 = subckt_1601_sff1_x4.sff_m
* NET 6160 = abc_8311_auto_rtlil_cc_2693_muxgate_8194
* NET 6163 = subckt_1601_sff1_x4.ckr
* NET 6164 = subckt_1601_sff1_x4.nckr
* NET 6165 = adrs[3]
* NET 6166 = abc_8311_new_n1686
* NET 6167 = abc_8311_new_n1685
* NET 6169 = abc_8311_new_n1480
* NET 6170 = abc_8311_new_n1479
* NET 6172 = abc_8311_new_n863
* NET 6173 = abc_8311_new_n873
* NET 6175 = abc_8311_new_n1496
* NET 6176 = abc_8311_new_n1495
* NET 6177 = abc_8311_new_n1488
* NET 6178 = abc_8311_new_n1669
* NET 6180 = abc_8311_new_n1668
* NET 6182 = abc_8311_new_n1358
* NET 6183 = abc_8311_new_n1261
* NET 6184 = abc_8311_new_n1667
* NET 6186 = abc_8311_new_n1206
* NET 6187 = dl[3]
* NET 6188 = abc_8311_new_n1443
* NET 6190 = abc_8311_new_n838
* NET 6191 = abc_8311_new_n848
* NET 6194 = subckt_1563_sff1_x4.sff_s
* NET 6197 = abc_8311_auto_rtlil_cc_2693_muxgate_8118
* NET 6200 = subckt_1563_sff1_x4.sff_m
* NET 6201 = subckt_1563_sff1_x4.ckr
* NET 6202 = subckt_1563_sff1_x4.nckr
* NET 6203 = abc_8311_new_n1653
* NET 6204 = abc_8311_new_n1657
* NET 6205 = abc_8311_new_n1655
* NET 6207 = abc_8311_new_n1654
* NET 6208 = abc_8311_new_n1455
* NET 6209 = abc_8311_new_n1458
* NET 6211 = abc_8311_new_n1452
* NET 6212 = abc_8311_new_n673
* NET 6214 = abc_8311_new_n337
* NET 6216 = abc_8311_new_n994
* NET 6219 = abc_8311_new_n552
* NET 6220 = abc_8311_new_n1218
* NET 6221 = abc_8311_new_n346
* NET 6222 = abc_8311_new_n1336
* NET 6224 = abc_8311_new_n259
* NET 6225 = abc_8311_new_n1304
* NET 6226 = abc_8311_new_n294
* NET 6229 = subckt_1554_sff1r_x4.sff_s
* NET 6232 = abc_8311_auto_rtlil_cc_2693_muxgate_8100
* NET 6233 = subckt_1554_sff1r_x4.sff_m
* NET 6235 = subckt_1554_sff1r_x4.ckr
* NET 6237 = subckt_1554_sff1r_x4.nckr
* NET 6238 = abc_8311_new_n1208
* NET 6242 = abc_8311_auto_ff_cc_704_flip_bits_8297
* NET 6243 = irq
* NET 6245 = abc_8311_new_n1294
* NET 6247 = abc_8311_new_n1296
* NET 6250 = abc_8311_new_n1300
* NET 6252 = subckt_1636_sff1r_x4.sff_s
* NET 6254 = subckt_1636_sff1r_x4.sff_m
* NET 6256 = abc_8311_auto_rtlil_cc_2693_muxgate_8296
* NET 6259 = subckt_1636_sff1r_x4.ckr
* NET 6260 = subckt_1636_sff1r_x4.nckr
* NET 6261 = nmi
* NET 6263 = nm1
* NET 6265 = data[1]
* NET 6310 = abc_8311_new_n264
* NET 6322 = subckt_1565_sff1_x4.sff_s
* NET 6326 = abc_8311_auto_rtlil_cc_2693_muxgate_8122
* NET 6327 = subckt_1565_sff1_x4.sff_m
* NET 6330 = subckt_1565_sff1_x4.ckr
* NET 6331 = subckt_1565_sff1_x4.nckr
* NET 6332 = subckt_1564_sff1_x4.sff_s
* NET 6336 = abc_8311_auto_rtlil_cc_2693_muxgate_8120
* NET 6338 = subckt_1564_sff1_x4.sff_m
* NET 6340 = subckt_1564_sff1_x4.ckr
* NET 6341 = subckt_1564_sff1_x4.nckr
* NET 6342 = abc_8311_new_n1534
* NET 6347 = abc_8311_new_n1520
* NET 6348 = abc_8311_new_n1517
* NET 6352 = abc_8311_new_n281
* NET 6357 = abc_8311_new_n1675
* NET 6359 = abc_8311_new_n1545
* NET 6360 = abc_8311_new_n1684
* NET 6362 = abc_8311_new_n1512
* NET 6363 = abc_8311_new_n1504
* NET 6364 = abc_8311_new_n1511
* NET 6371 = abc_8311_new_n1683
* NET 6372 = abc_8311_new_n1467
* NET 6374 = abc_8311_new_n1453
* NET 6375 = abc_8311_new_n1450
* NET 6376 = adrs[1]
* NET 6381 = subckt_1598_sff1_x4.sff_s
* NET 6384 = abc_8311_auto_rtlil_cc_2693_muxgate_8188
* NET 6385 = subckt_1598_sff1_x4.sff_m
* NET 6387 = subckt_1598_sff1_x4.ckr
* NET 6389 = subckt_1598_sff1_x4.nckr
* NET 6390 = abc_8311_new_n1666
* NET 6393 = abc_8311_new_n1487
* NET 6398 = abc_8311_new_n1659
* NET 6400 = abc_8311_new_n1663
* NET 6401 = abc_8311_new_n1661
* NET 6405 = abc_8311_new_n1662
* NET 6410 = abc_8311_new_n1647
* NET 6413 = abc_8311_new_n1648
* NET 6414 = abc_8311_new_n1649
* NET 6417 = abc_8311_new_n1651
* NET 6418 = abc_8311_new_n1650
* NET 6420 = abc_8311_new_n1334
* NET 6421 = abc_8311_new_n1341
* NET 6422 = abc_8311_new_n1269
* NET 6423 = abc_8311_new_n1451
* NET 6424 = abc_8311_new_n1457
* NET 6426 = abc_8311_new_n1475
* NET 6430 = abc_8311_new_n993
* NET 6431 = abc_8311_new_n1507
* NET 6434 = abc_8311_new_n438
* NET 6440 = rdy
* NET 6442 = ift_run
* NET 6447 = abc_8311_new_n291
* NET 6448 = abc_8311_new_n551
* NET 6449 = abc_8311_new_n1215
* NET 6455 = subckt_1553_sff1r_x4.sff_s
* NET 6457 = subckt_1553_sff1r_x4.sff_m
* NET 6461 = subckt_1553_sff1r_x4.ckr
* NET 6462 = subckt_1553_sff1r_x4.nckr
* NET 6463 = abc_8311_auto_rtlil_cc_2693_muxgate_8098
* NET 6464 = abc_8311_new_n1308
* NET 6466 = abc_8311_new_n1295
* NET 6469 = abc_8311_new_n244
* NET 6471 = abc_8311_new_n295
* NET 6473 = abc_8311_new_n1297
* NET 6475 = abc_8311_new_n1299
* NET 6476 = abc_8311_new_n243
* NET 6477 = abc_8311_new_n1223
* NET 6480 = do_res
* NET 6483 = subckt_1550_sff1r_x4.sff_s
* NET 6487 = subckt_1550_sff1r_x4.sff_m
* NET 6490 = subckt_1550_sff1r_x4.ckr
* NET 6491 = datao[0]
* NET 6492 = subckt_1550_sff1r_x4.nckr
* NET 6522 = adrs[2]
* NET 6571 = adrs[0]
* NET 6573 = subckt_1556_sff1_x4.sff_s
* NET 6575 = subckt_1556_sff1_x4.sff_m
* NET 6578 = subckt_1556_sff1_x4.ckr
* NET 6580 = m_clock_root_br_1
* NET 6581 = abc_8311_new_n261
* NET 6582 = subckt_1556_sff1_x4.nckr
* NET 6585 = abc_8311_new_n1372
* NET 6586 = abc_8311_new_n1369
* NET 6588 = abc_8311_new_n1367
* NET 6589 = abc_8311_auto_rtlil_cc_2693_muxgate_8104
* NET 6590 = abc_8311_new_n1350
* NET 6591 = debug[7]
* NET 6593 = abc_8311_new_n1376
* NET 6594 = abc_8311_new_n1374
* NET 6596 = abc_8311_new_n1375
* NET 6598 = abc_8311_new_n287
* NET 6600 = abc_8311_new_n1360
* NET 6601 = abc_8311_new_n1207
* NET 6603 = abc_8311_new_n286
* NET 6607 = abc_8311_new_n1533
* NET 6609 = abc_8311_new_n1531
* NET 6613 = abc_8311_new_n1519
* NET 6616 = abc_8311_new_n1349
* NET 6619 = abc_8311_new_n1546
* NET 6622 = abc_8311_new_n1348
* NET 6624 = abc_8311_new_n1543
* NET 6627 = abc_8311_new_n1678
* NET 6628 = abc_8311_new_n1681
* NET 6629 = abc_8311_new_n1679
* NET 6631 = abc_8311_new_n1646
* NET 6632 = abc_8311_new_n1503
* NET 6636 = abc_8311_new_n1472
* NET 6637 = abc_8311_new_n1337
* NET 6640 = abc_8311_new_n1469
* NET 6644 = abc_8311_new_n1471
* NET 6648 = abc_8311_new_n1484
* NET 6650 = subckt_1597_sff1_x4.sff_s
* NET 6652 = abc_8311_auto_rtlil_cc_2693_muxgate_8186
* NET 6655 = subckt_1597_sff1_x4.sff_m
* NET 6657 = subckt_1597_sff1_x4.ckr
* NET 6658 = subckt_1597_sff1_x4.nckr
* NET 6660 = abc_8311_new_n1660
* NET 6661 = abc_8311_new_n1483
* NET 6665 = debug[10]
* NET 6667 = abc_8311_new_n1656
* NET 6668 = abc_8311_new_n1470
* NET 6675 = abc_8311_new_n1456
* NET 6676 = abc_8311_new_n1468
* NET 6678 = abc_8311_new_n1335
* NET 6680 = abc_8311_new_n1474
* NET 6682 = do_brk
* NET 6685 = abc_8311_new_n1491
* NET 6688 = abc_8311_new_n1490
* NET 6690 = abc_8311_new_n1224
* NET 6691 = abc_8311_new_n1222
* NET 6692 = abc_8311_new_n1307
* NET 6694 = do_nmi
* NET 6695 = abc_8311_new_n274
* NET 6696 = abc_8311_new_n1309
* NET 6700 = abc_8311_new_n351
* NET 6701 = abc_8311_new_n1217
* NET 6702 = abc_8311_new_n1214
* NET 6703 = abc_8311_new_n338
* NET 6704 = abc_8311_new_n1212
* NET 6705 = abc_8311_new_n1221
* NET 6706 = abc_8311_new_n1298
* NET 6707 = abc_8311_new_n1228
* NET 6711 = abc_8311_new_n335
* NET 6713 = abc_8311_new_n1209
* NET 6714 = int_req
* NET 6715 = abc_8311_new_n439
* NET 6717 = subckt_1541_sff1r_x4.sff_s
* NET 6720 = subckt_1541_sff1r_x4.sff_m
* NET 6723 = subckt_1541_sff1r_x4.ckr
* NET 6724 = subckt_1541_sff1r_x4.nckr
* NET 6725 = abc_8311_new_n1302
* NET 6726 = abc_8311_auto_rtlil_cc_2693_muxgate_8092
* NET 6727 = data[0]
* NET 6728 = start
* NET 6740 = debug[6]
* NET 6748 = abc_8311_new_n851
* NET vdd = vdd
* NET 6777 = abc_8311_new_n1373
* NET 6778 = abc_8311_new_n1351
* NET 6781 = subckt_1555_sff1_x4.sff_s
* NET 6784 = subckt_1555_sff1_x4.sff_m
* NET 6786 = abc_8311_auto_rtlil_cc_2693_muxgate_8102
* NET 6789 = subckt_1555_sff1_x4.ckr
* NET 6790 = subckt_1555_sff1_x4.nckr
* NET 6791 = abc_8311_new_n1340
* NET 6792 = abc_8311_new_n1352
* NET 6794 = abc_8311_new_n1342
* NET 6798 = abc_8311_new_n1368
* NET 6800 = abc_8311_new_n1365
* NET 6801 = abc_8311_new_n1364
* NET 6802 = abc_8311_new_n1354
* NET 6806 = abc_8311_new_n1355
* NET 6807 = debug[8]
* NET 6808 = abc_8311_new_n1363
* NET 6811 = abc_8311_new_n278
* NET 6814 = abc_8311_new_n1347
* NET 6817 = abc_8311_new_n1532
* NET 6819 = abc_8311_new_n1680
* NET 6820 = debug[5]
* NET 6821 = abc_8311_new_n1530
* NET 6825 = subckt_1599_sff1_x4.sff_s
* NET 6827 = subckt_1599_sff1_x4.sff_m
* NET 6830 = abc_8311_auto_rtlil_cc_2693_muxgate_8190
* NET 6832 = m_clock_root_br_0
* NET 6833 = subckt_1599_sff1_x4.ckr
* NET 6834 = subckt_1599_sff1_x4.nckr
* NET 6835 = abc_8311_new_n276
* NET 6839 = abc_8311_new_n1346
* NET 6841 = abc_8311_new_n1674
* NET 6842 = abc_8311_new_n1672
* NET 6843 = abc_8311_new_n1673
* NET 6847 = abc_8311_new_n1518
* NET 6849 = abc_8311_new_n1671
* NET 6850 = debug[4]
* NET 6851 = abc_8311_new_n1516
* NET 6855 = abc_8311_new_n1500
* NET 6858 = abc_8311_new_n1502
* NET 6861 = abc_8311_new_n271
* NET 6866 = abc_8311_new_n1501
* NET 6867 = abc_8311_new_n1338
* NET 6869 = abc_8311_new_n1665
* NET 6870 = abc_8311_new_n1345
* NET 6874 = debug[3]
* NET 6875 = abc_8311_new_n1499
* NET 6876 = abc_8311_new_n1339
* NET 6877 = abc_8311_new_n1318
* NET 6883 = abc_8311_new_n1486
* NET 6885 = debug[2]
* NET 6886 = abc_8311_new_n267
* NET 6889 = abc_8311_new_n1485
* NET 6890 = abc_8311_new_n1344
* NET 6893 = debug[1]
* NET 6895 = subckt_1596_sff1_x4.sff_s
* NET 6898 = subckt_1596_sff1_x4.sff_m
* NET 6900 = abc_8311_auto_rtlil_cc_2693_muxgate_8184
* NET 6901 = subckt_1596_sff1_x4.ckr
* NET 6903 = abc_8311_new_n262
* NET 6904 = subckt_1596_sff1_x4.nckr
* NET 6905 = debug[9]
* NET 6906 = debug[0]
* NET 6908 = subckt_1595_sff1_x4.sff_s
* NET 6910 = abc_8311_new_n1362
* NET 6912 = subckt_1595_sff1_x4.sff_m
* NET 6914 = abc_8311_auto_rtlil_cc_2693_muxgate_8182
* NET 6916 = subckt_1595_sff1_x4.ckr
* NET 6917 = abc_8311_new_n334
* NET 6918 = subckt_1595_sff1_x4.nckr
* NET 6919 = abc_8311_new_n358
* NET 6921 = abc_8311_new_n242
* NET 6923 = subckt_1552_sff1r_x4.sff_s
* NET 6928 = subckt_1552_sff1r_x4.sff_m
* NET 6930 = abc_8311_auto_rtlil_cc_2693_muxgate_8096
* NET 6932 = subckt_1552_sff1r_x4.ckr
* NET 6933 = subckt_1552_sff1r_x4.nckr
* NET 6934 = do_irq
* NET 6935 = abc_8311_new_n273
* NET 6939 = subckt_1539_sff1r_x4.sff_s
* NET 6942 = subckt_1539_sff1r_x4.sff_m
* NET 6945 = subckt_1539_sff1r_x4.ckr
* NET 6946 = abc_8311_auto_rtlil_cc_2693_muxgate_8070
* NET 6947 = subckt_1539_sff1r_x4.nckr
* NET 6948 = abc_8311_new_n1220
* NET 6951 = abc_8311_new_n361
* NET 6952 = reg_762[2]
* NET 6956 = abc_8311_new_n241
* NET 6957 = abc_8311_new_n1219
* NET 6959 = abc_8311_new_n1225
* NET 6962 = abc_8311_new_n359
* NET 6963 = reg_762[0]
* NET 6966 = abc_8311_new_n1232
* NET 6967 = abc_8311_auto_rtlil_cc_2693_muxgate_8074
* NET 6968 = abc_8311_new_n1231
* NET 6970 = abc_8311_new_n1229
* NET 6972 = abc_8311_new_n1227
* NET 6974 = reg_762[1]
* NET 6976 = p_reset
* NET 6978 = subckt_1540_sff1r_x4.sff_s
* NET 6981 = abc_8311_auto_rtlil_cc_2693_muxgate_8072
* NET 6982 = subckt_1540_sff1r_x4.sff_m
* NET 6984 = m_clock_root_bl_0
* NET 6986 = subckt_1540_sff1r_x4.ckr
* NET vss = vss
* NET 6988 = subckt_1540_sff1r_x4.nckr
Mtr_13918 6766 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13917 6855 6877 6766 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13916 vdd 6874 6855 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13915 214 2314 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13914 214 493 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13913 vdd 615 214 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13912 210 2314 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13911 210 493 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13910 vdd 787 210 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13909 6699 6952 6917 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13908 6698 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13907 vdd 6698 6699 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13906 6443 6934 6297 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13905 6297 6694 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13904 vdd 6442 6443 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13903 6449 6443 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13902 4036 4275 4035 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13901 4033 4032 4036 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13900 4034 4708 4033 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13899 vdd 6224 4034 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13898 4228 4035 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13897 861 2195 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13896 1039 2194 861 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13895 vdd 1033 1039 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13894 vdd 5068 4448 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13893 4448 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13892 4448 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13891 vdd 5272 4448 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13890 4447 4448 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13889 6763 6817 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13888 6819 6821 6763 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13887 vdd 6867 6819 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13886 vdd 6740 6617 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13885 6617 6839 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13884 6617 6820 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13883 vdd 6850 6617 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13882 6616 6617 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13881 1180 1339 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13880 vdd 1329 1180 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13879 1326 1180 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13878 5677 5676 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13877 5672 5678 5671 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13876 vdd 5670 5672 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13875 5674 5678 5677 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13874 5675 5679 5674 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13873 vdd 5673 5675 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13872 5673 5674 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13871 5671 5679 5673 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13870 vdd 5671 5670 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13869 5670 5671 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13868 vdd 6580 5679 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13867 5678 5679 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13866 vdd 5682 5676 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13865 vdd 4649 4162 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13864 4160 4918 4120 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13863 4120 4649 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13862 4120 4162 4160 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13861 vdd 4158 4120 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13860 4158 4918 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13859 vdd 489 211 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13858 211 209 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13857 vdd 210 211 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13856 477 211 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13855 vdd 6430 6217 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13854 6217 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13853 vdd 6917 6217 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13852 6216 6217 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13851 1211 1210 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13850 vdd 1360 1211 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13849 1322 1211 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13848 262 265 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13847 vdd 263 262 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13846 395 262 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13845 3181 3184 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13844 vdd 3183 3181 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13843 3182 3181 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13842 2528 2526 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13841 vdd 2525 2528 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13840 2752 2528 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13839 6654 6656 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13838 6649 6657 6650 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13837 vdd 6885 6649 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13836 6655 6657 6654 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13835 6653 6658 6655 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13834 vdd 6651 6653 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13833 6651 6655 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13832 6650 6658 6651 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13831 vdd 6650 6885 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13830 6885 6650 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13829 vdd 6984 6658 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13828 6657 6658 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13827 vdd 6652 6656 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13826 3000 2997 2874 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13825 2874 2999 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13824 vdd 2998 3000 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13823 4737 3000 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13822 2835 2833 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13821 vdd 2834 2835 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13820 2837 2835 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13819 5989 6219 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13818 vdd 6917 5989 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13817 5987 5989 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13816 5757 5805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13815 5763 5756 5757 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13814 vdd 6807 5763 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13813 vdd 5305 4017 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13812 4017 4015 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13811 vdd 4016 4017 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13810 4014 4017 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13809 vdd 6434 3669 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13808 3669 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13807 3734 5262 3669 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13806 3668 4217 3734 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13805 3669 5502 3668 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13804 4541 4666 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13803 4539 4585 4664 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13802 vdd 4914 4539 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13801 4584 4585 4541 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13800 4540 4586 4584 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13799 vdd 4582 4540 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13798 4582 4584 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13797 4664 4586 4582 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13796 vdd 4664 4914 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13795 4914 4664 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13794 vdd 6580 4586 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13793 4585 4586 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13792 vdd 4665 4666 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13791 2018 2046 2508 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13790 2017 2045 2018 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13789 vdd 2044 2017 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13788 4251 4491 4110 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13787 4110 4250 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13786 vdd 5349 4251 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13785 4572 4251 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13784 vdd 4941 4070 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13783 4070 4287 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13782 4070 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13781 vdd 4524 4070 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13780 4265 4070 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13779 2490 3741 2424 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13778 vdd 2733 2424 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13777 2424 2739 2490 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13776 2489 2490 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13775 vdd 5761 5328 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13774 5328 5327 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13773 5328 5985 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13772 vdd 5326 5328 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13771 5762 5328 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13770 vdd 5334 5033 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13769 5054 5033 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13768 vdd 5033 5054 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13767 vdd 5033 5054 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13766 5054 5033 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13765 vdd 5334 1571 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13764 3259 1571 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13763 vdd 1571 3259 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13762 vdd 1571 3259 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13761 3259 1571 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13760 vdd 5334 1570 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13759 1569 1570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13758 vdd 1570 1569 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13757 vdd 1570 1569 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13756 1569 1570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13755 vdd 5334 1371 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13754 1370 1371 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13753 vdd 1371 1370 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13752 vdd 1371 1370 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13751 1370 1371 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13750 vdd 5334 1512 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13749 3160 1512 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13748 vdd 1512 3160 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13747 vdd 1512 3160 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13746 3160 1512 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13745 vdd 5334 1511 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13744 1510 1511 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13743 vdd 1511 1510 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13742 vdd 1511 1510 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13741 1510 1511 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13740 vdd 5334 1316 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13739 1315 1316 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13738 vdd 1316 1315 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13737 vdd 1316 1315 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13736 1315 1316 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13735 vdd 6890 6891 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13734 6889 6886 6771 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13733 6771 6890 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13732 6771 6891 6889 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13731 vdd 6887 6771 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13730 6887 6886 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13729 6674 6877 6675 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13728 6673 6876 6674 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13727 vdd 6903 6673 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13726 vdd 4089 1762 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13725 1762 2352 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13724 1762 4087 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13723 vdd 4299 1762 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13722 1760 1762 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13721 2978 3160 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13720 vdd 2978 2976 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13719 2975 2977 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13718 vdd 2975 2870 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13717 2870 2976 2973 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13716 2973 2978 2869 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13715 2868 2979 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13714 vdd 2970 2979 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13713 2979 2970 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13712 2869 2971 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13711 2971 2973 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13710 vdd 6976 2971 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13709 2970 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13708 2970 2976 2868 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13707 2971 2978 2970 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13706 4177 6600 4099 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13705 4099 4176 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13704 vdd 6601 4177 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13703 4397 4177 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13702 6126 6877 6125 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13701 6125 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13700 vdd 6665 6126 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13699 6127 6126 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13698 5168 5106 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13697 vdd 5104 5168 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13696 5754 5753 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13695 5755 5767 5754 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13694 vdd 6807 5755 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13693 4976 5044 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13692 5265 5045 4976 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13691 vdd 5965 5265 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13690 6197 5972 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13689 vdd 5969 6197 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13688 2048 2508 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13687 vdd 2507 2048 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13686 3550 3546 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13685 3550 3947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13684 vdd 6423 3550 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13683 260 261 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13682 vdd 399 260 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13681 830 260 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13680 4143 4501 4274 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13679 4142 4275 4143 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13678 vdd 4273 4142 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13677 4512 4274 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13676 4575 6469 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13675 6877 4733 4575 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13674 vdd 4731 6877 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13673 570 569 542 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13672 542 579 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13671 vdd 2727 570 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13670 1313 570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13669 3592 4909 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13668 vdd 3788 3592 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13667 vdd 3460 2457 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13666 2458 4299 4941 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13665 2456 5157 2458 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13664 2457 2852 2456 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13663 2379 1365 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13662 vdd 3226 2379 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13661 1730 1732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13660 vdd 1760 1730 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13659 5792 2138 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13658 5792 1944 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13657 vdd 2139 5792 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13656 6477 6952 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13655 6477 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13654 vdd 6714 6477 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13653 vdd 6963 6477 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13652 vdd 5880 5843 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13651 5843 6216 5984 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13650 5983 5984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13649 vdd 3964 3551 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13648 3551 3550 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13647 vdd 5003 3551 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13646 3549 3551 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13645 4066 4953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13644 4066 4257 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13643 vdd 4072 4066 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13642 5309 3424 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13641 5309 3621 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13640 vdd 3622 5309 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13639 5693 5723 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13638 5862 5721 5693 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13637 vdd 5965 5862 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13636 vdd 4502 4504 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13635 4504 4510 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13634 vdd 4503 4504 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13633 4618 4504 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13632 2345 2331 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13631 2345 2136 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13630 vdd 2135 2345 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13629 5748 2173 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13628 5748 1744 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13627 vdd 1562 5748 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13626 vdd 1563 5748 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13625 vdd 4235 2389 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13624 vdd 4748 2390 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13623 2389 2390 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13622 1044 1991 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13621 vdd 5363 1044 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13620 1953 1044 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13619 vdd 5068 4907 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13618 4907 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13617 4907 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13616 vdd 6727 4907 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13615 4906 4907 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13614 2144 2532 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13613 2144 2544 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13612 vdd 2142 2144 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13611 1494 1891 1493 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13610 1493 1885 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13609 vdd 1882 1494 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13608 1492 1494 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13607 4841 5011 4842 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13606 4842 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13605 vdd 6678 4842 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13604 4838 4841 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13603 4840 6637 4841 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13602 4842 4839 4840 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13601 vdd 5115 5118 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13600 5118 5770 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13599 5118 5331 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13598 vdd 5116 5118 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13597 6910 5118 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13596 3294 4477 3420 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13595 3293 4456 3294 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13594 vdd 5987 3293 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13593 3740 3420 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13592 1641 3217 1598 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13591 1598 2535 1641 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13590 vdd 1640 1598 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13589 5683 6172 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13588 5856 6173 5683 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13587 vdd 5927 5856 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13586 1692 1925 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13585 vdd 1694 1692 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13584 2763 1692 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13583 2130 2128 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13582 vdd 2144 2130 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13581 2340 2130 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13580 1901 2501 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13579 vdd 2782 1901 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13578 1900 1901 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13577 3157 3159 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13576 3154 3161 3153 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13575 vdd 3379 3154 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13574 3158 3161 3157 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13573 3155 3162 3158 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13572 vdd 3156 3155 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13571 3156 3158 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13570 3153 3162 3156 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13569 vdd 3153 3379 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13568 3379 3153 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13567 vdd 3160 3162 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13566 3161 3162 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13565 vdd 3163 3159 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13564 vdd 6778 6779 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13563 6777 6905 6759 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13562 6759 6778 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13561 6759 6779 6777 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13560 vdd 6775 6759 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13559 6775 6905 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13558 1927 2122 1928 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13557 1928 2124 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13556 vdd 2125 1928 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13555 2128 1927 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13554 1926 1929 1927 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13553 1928 2532 1926 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13552 3219 3792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13551 3430 3793 3219 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13550 vdd 3434 3430 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13549 4113 4296 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13548 4111 4297 4290 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13547 vdd 4299 4111 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13546 4293 4297 4113 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13545 4112 4298 4293 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13544 vdd 4292 4112 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13543 4292 4293 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13542 4290 4298 4292 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13541 vdd 4290 4299 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13540 4299 4290 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13539 vdd 6984 4298 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13538 4297 4298 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13537 vdd 4300 4296 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13536 1259 1338 1339 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13535 1258 1343 1259 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13534 vdd 1533 1258 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13533 vdd 5341 4244 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13532 4244 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13531 vdd 6440 4244 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13530 4477 4244 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13529 862 1390 864 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13528 864 863 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13527 vdd 3263 862 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13526 860 862 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13525 vdd 2194 1349 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13524 1349 1553 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13523 1349 1953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13522 vdd 3836 1349 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13521 2122 1349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13520 2103 2314 2012 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13519 2012 2511 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13518 vdd 2111 2012 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13517 2102 2103 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13516 2011 3740 2103 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13515 2012 2512 2011 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13514 vdd 4009 4011 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13513 4011 5500 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13512 vdd 4010 4011 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13511 4008 4011 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13510 5698 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13509 5699 6877 5698 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13508 vdd 6591 5699 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13507 5743 6182 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13506 6413 6183 5743 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13505 vdd 5742 6413 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13504 3806 3805 3697 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13503 3697 3819 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13502 vdd 5102 3806 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13501 4611 3806 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13500 4050 5502 4471 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13499 4049 4052 4050 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13498 vdd 4048 4049 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13497 vdd 5069 2388 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13496 2388 2807 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13495 2388 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13494 vdd 6440 2388 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13493 2387 2388 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13492 2428 2514 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_13491 3183 2513 2428 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_13490 2427 2512 3183 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_13489 vdd 2511 2427 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_13488 3163 3555 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13487 vdd 3736 3163 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13486 3349 5054 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13485 vdd 3349 3350 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13484 3348 3397 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13483 vdd 3348 3275 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13482 3275 3350 3347 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13481 3347 3349 3276 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13480 3283 3403 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13479 vdd 3396 3403 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13478 3403 3396 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13477 3276 3344 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13476 3344 3347 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13475 vdd 6976 3344 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13474 3396 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13473 3396 3350 3283 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13472 3344 3349 3396 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13471 12 119 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13470 10 45 115 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13469 vdd 392 10 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13468 43 45 12 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13467 11 120 43 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13466 vdd 42 11 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13465 42 43 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13464 115 120 42 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13463 vdd 115 392 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13462 392 115 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13461 vdd 3259 120 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13460 45 120 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13459 vdd 243 119 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13458 5261 5524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13457 5261 6910 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13456 vdd 6806 5261 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13455 vdd 6480 5849 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13454 5849 6682 6012 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13453 6464 6012 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13452 3622 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13451 vdd 4233 3622 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13450 1506 2950 1507 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13449 1507 2946 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13448 vdd 2111 1506 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13447 1505 1506 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13446 1361 4051 1270 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13445 1270 2799 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13444 vdd 3813 1361 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13443 1360 1361 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13442 4938 5112 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13441 5534 5113 4938 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13440 vdd 4937 5534 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13439 3152 3552 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13438 vdd 3165 3152 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13437 5832 6182 6631 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13436 5831 6188 5832 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13435 vdd 6183 5831 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13434 4858 4857 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13433 4863 4859 4858 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13432 vdd 6867 4863 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13431 6602 6600 6604 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13430 6604 6603 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13429 vdd 6601 6602 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13428 6801 6602 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13427 917 1517 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13426 vdd 1518 917 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13425 1330 1339 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13424 vdd 1329 1330 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13423 1653 2553 1591 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13422 1591 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13421 vdd 2314 1653 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13420 1652 1653 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13419 3814 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13418 3814 2807 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13417 vdd 5069 3814 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13416 3456 2833 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13415 vdd 2834 3456 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13414 2303 2299 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13413 vdd 2489 2303 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13412 2307 2306 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13411 vdd 2492 2307 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13410 5402 5510 5500 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13409 5499 5498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13408 vdd 5499 5402 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13407 5700 6375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13406 5700 6374 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13405 vdd 6423 5700 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13404 vdd 5501 5700 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13403 6900 6204 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13402 vdd 6203 6900 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13401 4866 4914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13400 4866 6910 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13399 vdd 6806 4866 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13398 308 307 270 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13397 270 598 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13396 vdd 470 308 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13395 588 308 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13394 2194 2628 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13393 vdd 2625 2194 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13392 6823 6877 6735 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13391 6735 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13390 vdd 6820 6823 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13389 6821 6823 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13388 6914 6417 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13387 vdd 6418 6914 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13386 5492 5490 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13385 vdd 5489 5492 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13384 6176 5492 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13383 5142 5141 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13382 vdd 5140 5142 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13381 5570 5142 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13380 4498 5341 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13379 vdd 5773 4498 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13378 4497 4498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13377 4021 4461 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13376 vdd 4020 4021 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13375 1670 2331 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13374 1670 1676 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13373 vdd 1667 1670 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13372 3813 3818 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13371 3813 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13370 vdd 5069 3813 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13369 vdd 6819 6630 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13368 6630 6629 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13367 vdd 6627 6630 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13366 6628 6630 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13365 vdd 5867 5477 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13364 5477 5955 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13363 vdd 5485 5477 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13362 5474 5477 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13361 vdd 6129 5920 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13360 5920 5919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13359 vdd 5925 5920 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13358 5918 5920 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13357 2512 2550 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13356 2512 2986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13355 vdd 1541 2512 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13354 vdd 1542 2512 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13353 5269 6375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13352 5269 6374 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13351 vdd 6423 5269 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13350 vdd 5268 5269 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13349 vdd 6691 6693 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13348 6693 6692 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13347 6693 6695 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13346 vdd 6921 6693 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13345 6696 6693 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13344 1342 3408 1260 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13343 1260 1340 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13342 vdd 2521 1342 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13341 1699 1342 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13340 vdd 488 331 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13339 328 779 275 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13338 275 488 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13337 275 331 328 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13336 vdd 329 275 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13335 329 779 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13334 vdd 4456 4130 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13333 4130 4477 4223 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13332 5300 4223 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13331 2839 3263 4088 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13330 2838 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13329 vdd 2838 2839 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13328 6212 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13327 6212 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13326 vdd 6376 6212 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13325 vdd 6440 6212 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13324 5750 6893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13323 5750 5748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13322 vdd 5749 5750 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13321 vdd 6440 5750 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13320 6237 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13319 vdd 6237 6235 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13318 6236 6232 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13317 vdd 6236 6234 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13316 6234 6235 6233 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13315 6233 6237 6231 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13314 6228 6442 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13313 vdd 6229 6442 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13312 6442 6229 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13311 6231 6230 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13310 6230 6233 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13309 vdd 6976 6230 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13308 6229 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13307 6229 6235 6228 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13306 6230 6237 6229 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13305 vdd 5127 5129 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13304 5129 5132 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13303 5129 5343 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13302 vdd 5342 5129 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13301 5141 5129 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13300 vdd 3449 3302 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13299 3302 3455 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13298 4233 3863 3302 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13297 3301 4071 4233 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13296 3302 3458 3301 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13295 2898 2896 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13294 vdd 2897 2898 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13293 2895 2898 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13292 1577 1578 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13291 1575 1757 1577 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13290 vdd 4241 1575 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13289 vdd 4649 4166 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13288 4855 4163 4121 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13287 4121 4649 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13286 4121 4166 4855 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13285 vdd 4164 4121 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13284 4164 4163 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13283 775 1652 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13282 vdd 1505 775 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13281 774 775 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13280 3196 3591 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13279 vdd 3201 3196 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13278 3195 3196 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13277 1651 1649 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13276 vdd 2086 1651 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13275 5949 1651 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13274 5945 5943 5819 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13273 5819 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13272 vdd 6678 5819 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13271 5942 5945 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13270 5818 6637 5945 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13269 5819 6619 5818 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13268 5376 5423 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13267 5374 5424 5417 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13266 vdd 6665 5374 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13265 5421 5424 5376 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13264 5375 5425 5421 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13263 vdd 5419 5375 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13262 5419 5421 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13261 5417 5425 5419 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13260 vdd 5417 6665 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13259 6665 5417 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13258 vdd 6580 5425 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13257 5424 5425 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13256 vdd 5857 5423 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13255 6744 6902 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13254 6742 6901 6895 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13253 vdd 6893 6742 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13252 6898 6901 6744 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13251 6743 6904 6898 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13250 vdd 6896 6743 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13249 6896 6898 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13248 6895 6904 6896 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13247 vdd 6895 6893 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13246 6893 6895 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13245 vdd 6984 6904 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13244 6901 6904 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13243 vdd 6900 6902 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13242 vdd 6934 6688 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13241 vdd 6694 6689 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13240 6688 6689 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13239 5816 6190 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13238 6144 6191 5816 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13237 vdd 5965 6144 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13236 vdd 6590 1624 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13235 6119 6807 1593 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13234 1593 6590 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13233 1593 1624 6119 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13232 vdd 1622 1593 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13231 1622 6807 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13230 594 603 564 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13229 564 1655 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13228 vdd 596 564 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13227 591 594 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13226 563 592 594 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13225 564 607 563 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13224 2831 2830 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13223 vdd 5069 2831 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13222 3649 2831 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13221 4408 4411 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13220 4404 4412 4405 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13219 vdd 4918 4404 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13218 4409 4412 4408 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13217 4407 4413 4409 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13216 vdd 4406 4407 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13215 4406 4409 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13214 4405 4413 4406 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13213 vdd 4405 4918 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13212 4918 4405 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13211 vdd 6580 4413 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13210 4412 4413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13209 vdd 4410 4411 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13208 273 480 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13207 317 477 273 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13206 272 482 317 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13205 vdd 478 272 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13204 766 317 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13203 1251 4176 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13202 1323 1322 1251 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13201 vdd 2747 1323 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13200 5347 5559 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13199 vdd 5346 5347 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13198 5345 5347 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13197 vdd 2307 2305 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13196 2305 2303 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13195 2304 2479 2305 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13194 2302 2319 2304 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13193 2305 2483 2302 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13192 vdd 5749 5316 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13191 5316 5748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13190 5316 6885 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13189 vdd 6440 5316 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13188 5315 5316 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13187 vdd 6839 6615 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13186 6613 6850 6614 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13185 6614 6839 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13184 6614 6615 6613 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13183 vdd 6612 6614 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13182 6612 6850 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13181 4551 4673 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13180 4672 4671 4551 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13179 vdd 5965 4672 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13178 6288 6420 6423 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13177 6289 6421 6288 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13176 vdd 6422 6289 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13175 4395 4396 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13174 vdd 4394 4395 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13173 vdd 619 614 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13172 611 1513 566 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13171 566 619 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13170 566 614 611 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13169 vdd 610 566 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13168 610 1513 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13167 526 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13166 2157 1190 526 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13165 vdd 525 2157 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13164 vdd 1688 1680 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13163 1680 3593 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13162 1680 2347 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13161 vdd 1679 1680 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13160 1682 1680 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13159 3329 5054 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13158 vdd 3329 3328 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13157 3327 3565 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13156 vdd 3327 3272 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13155 3272 3328 3326 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13154 3326 3329 3271 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13153 3279 3573 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13152 vdd 3385 3573 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13151 3573 3385 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13150 3271 3323 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13149 3323 3326 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13148 vdd 6976 3323 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13147 3385 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13146 3385 3328 3279 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13145 3323 3329 3385 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13144 2045 1669 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13143 vdd 1670 2045 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13142 5736 5735 5737 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13141 5734 5738 5736 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13140 vdd 5733 5734 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13139 vdd 4572 4449 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13138 4450 6186 4452 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13137 4451 6220 4450 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13136 4449 5300 4451 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13135 vdd 5502 3687 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13134 3688 4013 3947 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13133 3686 3797 3688 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13132 3687 4217 3686 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13131 285 2048 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13130 vdd 502 284 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13129 vdd 830 367 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13128 365 830 285 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13127 284 367 365 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13126 364 365 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13125 6291 6903 6425 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13124 6290 6877 6291 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13123 vdd 6876 6290 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13122 6424 6425 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13121 3216 4456 3217 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13120 3215 5987 3216 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13119 vdd 4477 3215 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13118 3715 3547 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13117 3715 3947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13116 vdd 6423 3715 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13115 187 2386 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13114 vdd 527 186 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13113 vdd 830 259 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13112 257 830 187 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13111 186 259 257 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13110 258 257 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13109 831 2793 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13108 vdd 829 833 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13107 vdd 830 834 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13106 832 830 831 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13105 833 834 832 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13104 828 832 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13103 813 2741 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13102 vdd 988 812 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13101 vdd 830 815 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13100 814 830 813 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13099 812 815 814 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13098 810 814 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13097 4502 4501 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13096 4502 5889 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13095 vdd 5773 4502 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13094 vdd 6440 4502 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13093 vdd 4083 2892 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13092 2892 4082 3047 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13091 3046 3047 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13090 3633 3632 3635 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13089 3635 3634 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13088 vdd 3636 3633 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13087 3631 3633 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13086 3951 3709 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13085 3951 3947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13084 vdd 6423 3951 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13083 177 917 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13082 vdd 636 176 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13081 vdd 1004 226 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13080 224 1004 177 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13079 176 226 224 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13078 225 224 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13077 520 1196 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13076 vdd 825 518 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13075 vdd 1004 521 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13074 519 1004 520 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13073 518 521 519 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13072 517 519 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13071 293 1208 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13070 vdd 522 292 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13069 vdd 1004 391 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13068 389 1004 293 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13067 292 391 389 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13066 387 389 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13065 2804 2803 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13064 vdd 4676 2802 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13063 vdd 3046 2806 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13062 2805 3046 2804 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13061 2802 2806 2805 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13060 2801 2805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13059 vdd 4726 3699 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13058 3699 5575 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13057 5115 4053 3699 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13056 3698 5992 5115 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13055 3699 5773 3698 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13054 5413 5999 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13053 5552 6000 5413 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13052 vdd 6440 5552 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13051 6948 6704 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13050 6948 6701 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13049 vdd 6702 6948 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13048 vdd 6700 6948 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13047 vdd 2553 1942 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13046 1942 2356 1943 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13045 2154 1943 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13044 965 1649 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13043 vdd 2086 965 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13042 6700 6963 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13041 6700 6917 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13040 vdd 6921 6700 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13039 4558 4689 4887 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13038 4690 4688 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13037 vdd 4690 4558 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13036 4680 4679 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13035 vdd 4682 4680 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13034 4878 4680 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13033 4073 4086 4074 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13032 vdd 4071 4074 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13031 4074 4281 4073 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13030 4072 4073 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13029 2281 2551 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13028 vdd 2361 2280 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13027 vdd 4673 2362 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13026 2359 4673 2281 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13025 2280 2362 2359 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13024 2360 2359 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13023 6966 6951 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13022 6966 6705 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13021 vdd 6704 6966 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13020 1704 2544 1609 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13019 1609 2142 1704 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13018 vdd 1703 1609 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13017 vdd 488 490 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13016 490 779 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13015 592 489 490 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13014 487 491 592 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13013 490 486 487 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13012 3205 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13011 3204 3414 3205 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13010 vdd 5262 3204 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13009 4065 4071 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_13008 4456 4708 4065 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_13007 4064 4261 4456 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_13006 vdd 6221 4064 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_13005 1367 4748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13004 1367 1732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13003 vdd 1218 1367 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13002 vdd 6843 6846 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13001 6846 6842 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13000 vdd 6849 6846 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12999 6841 6846 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12998 vdd 6591 5917 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12997 5917 6616 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12996 5917 6905 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12995 vdd 6807 5917 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12994 5914 5917 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12993 5814 5967 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12992 6132 5993 5814 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12991 vdd 5927 6132 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12990 5271 5947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12989 5324 5949 5271 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12988 vdd 5964 5324 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12987 2787 1953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12986 2787 857 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12985 vdd 2194 2787 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12984 vdd 3836 2787 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12983 1996 2852 2406 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12982 1995 3460 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12981 vdd 1995 1996 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12980 5844 5986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12979 5985 6214 5844 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12978 vdd 6893 5985 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12977 vdd 2919 2722 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12976 2938 2720 2721 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12975 2721 2919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12974 2721 2722 2938 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12973 vdd 2719 2721 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12972 2719 2720 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12971 5007 5008 4968 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12970 4968 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12969 vdd 6678 4968 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12968 5003 5007 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12967 4967 6637 5007 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12966 4968 5004 4967 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12965 3695 4275 3801 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12964 3696 3800 3695 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12963 3694 4708 3696 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12962 vdd 6224 3694 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12961 4463 3801 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12960 3203 3596 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12959 vdd 3204 3203 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12958 3202 3203 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12957 vdd 3062 3058 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12956 3058 4509 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12955 vdd 3060 3058 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12954 3632 3058 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12953 vdd 6186 5826 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12952 5826 6431 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12951 6629 5959 5826 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12950 5825 6182 6629 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12949 5826 6183 5825 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12948 6933 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12947 vdd 6933 6932 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12946 6931 6930 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12945 vdd 6931 6750 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12944 6750 6932 6928 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12943 6928 6933 6751 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12942 6749 6934 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12941 vdd 6923 6934 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12940 6934 6923 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12939 6751 6926 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12938 6926 6928 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12937 vdd 6976 6926 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12936 6923 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12935 6923 6932 6749 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12934 6926 6933 6923 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12933 6587 6585 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12932 6594 6586 6587 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12931 vdd 6867 6594 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12930 1930 2544 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12929 vdd 2142 1930 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12928 1929 1930 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12927 2759 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12926 vdd 4687 2759 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12925 2758 2759 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12924 796 2122 797 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12923 797 2124 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12922 vdd 2125 797 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12921 793 796 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12920 795 794 796 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12919 797 801 795 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12918 3845 4265 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12917 vdd 5773 3845 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12916 4082 3845 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12915 4516 4523 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12914 vdd 5144 4516 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12913 4517 4516 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12912 894 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12911 1931 987 894 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12910 vdd 988 1931 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12909 3175 3182 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12908 vdd 3174 3175 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12907 3570 3175 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12906 3562 5949 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12905 3561 5947 3562 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12904 vdd 3969 3561 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12903 2859 2906 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12902 2857 2907 2901 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12901 vdd 3376 2857 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12900 2903 2907 2859 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12899 2858 2908 2903 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12898 vdd 2902 2858 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12897 2902 2903 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12896 2901 2908 2902 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12895 vdd 2901 3376 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12894 3376 2901 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12893 vdd 3160 2908 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12892 2907 2908 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12891 vdd 3152 2906 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12890 2376 3006 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12889 vdd 3010 2376 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12888 2375 2376 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12887 5111 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12886 vdd 6917 5111 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12885 5113 5111 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12884 2190 2615 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12883 vdd 3818 2190 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12882 2195 2190 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12881 3690 4213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12880 3789 4212 3690 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12879 vdd 4696 3789 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12878 2492 3741 2425 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12877 2425 2739 2492 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12876 vdd 2733 2425 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12875 vdd 1320 1157 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12874 1157 1501 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12873 vdd 2314 1157 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12872 1156 1157 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12871 vdd 6778 6314 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12870 6585 6310 6266 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12869 6266 6778 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12868 6266 6314 6585 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12867 vdd 6312 6266 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12866 6312 6310 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12865 5793 5791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12864 5903 5792 5793 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12863 vdd 6250 5903 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12862 1250 2755 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12861 1317 3586 1250 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12860 vdd 2111 1317 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12859 3200 3199 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12858 3201 3618 3200 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12857 vdd 5959 3201 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12856 634 1190 543 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12855 543 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12854 vdd 633 634 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12853 918 634 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12852 3444 3632 3297 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12851 3297 3634 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12850 vdd 3442 3444 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12849 4947 3444 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12848 2089 2479 2005 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12847 2005 2303 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12846 vdd 2307 2005 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12845 2088 2089 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12844 2004 2319 2089 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12843 2005 2483 2004 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12842 3256 3258 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12841 3253 3261 3252 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12840 vdd 3460 3253 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12839 3257 3261 3256 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12838 3255 3260 3257 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12837 vdd 3254 3255 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12836 3254 3257 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12835 3252 3260 3254 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12834 vdd 3252 3460 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12833 3460 3252 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12832 vdd 3259 3260 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12831 3261 3260 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12830 vdd 3459 3258 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12829 807 808 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12828 802 809 803 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12827 vdd 988 802 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12826 806 809 807 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12825 805 811 806 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12824 vdd 804 805 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12823 804 806 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12822 803 811 804 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12821 vdd 803 988 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12820 988 803 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12819 vdd 3160 811 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12818 809 811 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12817 vdd 810 808 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12816 vdd 5268 4698 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12815 4698 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12814 4698 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12813 vdd 6440 4698 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12812 4699 4698 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12811 4139 4726 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12810 4507 4265 4139 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12809 vdd 5773 4507 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12808 3754 5054 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12807 vdd 3754 3753 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12806 3752 3750 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12805 vdd 3752 3675 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12804 3675 3753 3748 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12803 3748 3754 3674 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12802 3673 3972 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12801 vdd 3746 3972 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12800 3972 3746 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12799 3674 3747 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12798 3747 3748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12797 vdd 6976 3747 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12796 3746 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12795 3746 3753 3673 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12794 3747 3754 3746 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12793 288 374 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12792 286 377 369 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12791 vdd 663 286 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12790 372 377 288 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12789 287 376 372 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12788 vdd 371 287 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12787 371 372 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12786 369 376 371 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12785 vdd 369 663 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12784 663 369 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12783 vdd 3259 376 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12782 377 376 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12781 vdd 661 374 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12780 970 1649 881 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12779 881 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12778 vdd 1172 970 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12777 968 970 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12776 4476 6224 5112 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12775 4475 4708 4476 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12774 vdd 4524 4475 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12773 2095 2299 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12772 vdd 2492 2095 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12771 3666 5967 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12770 3948 5993 3666 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12769 vdd 3969 3948 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12768 3315 3717 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12767 vdd 3561 3315 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12766 3620 4611 3621 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12765 3619 4066 3620 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12764 vdd 3618 3619 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12763 5442 5670 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12762 5442 6910 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12761 vdd 6806 5442 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12760 1608 1704 2344 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12759 1607 1700 1608 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12758 vdd 1699 1607 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12757 2834 2615 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12756 vdd 3818 2834 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12755 2511 3741 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12754 vdd 2739 2511 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12753 6947 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12752 vdd 6947 6945 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12751 6944 6946 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12750 vdd 6944 6754 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12749 6754 6945 6942 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12748 6942 6947 6753 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12747 6752 6963 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12746 vdd 6939 6963 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12745 6963 6939 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12744 6753 6940 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12743 6940 6942 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12742 vdd 6976 6940 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12741 6939 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12740 6939 6945 6752 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12739 6940 6947 6939 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12738 5252 6877 5253 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12737 5253 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12736 vdd 5524 5252 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12735 5254 5252 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12734 4052 4051 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12733 vdd 4613 4052 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12732 3371 3658 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12731 vdd 4286 3371 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12730 2739 3186 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12729 vdd 5804 2739 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12728 2889 4737 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12727 3039 3042 2889 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12726 vdd 3044 3039 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12725 4651 5014 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12724 vdd 5026 4651 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12723 4649 4651 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12722 5340 5337 5339 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12721 vdd 5336 5339 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12720 5339 5338 5340 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12719 6232 5340 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12718 1196 1925 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12717 vdd 1694 1196 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12716 3585 3738 3587 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12715 3587 3737 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12714 vdd 4308 3585 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12713 3586 3585 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12712 1914 1911 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12711 1914 1687 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12710 vdd 1679 1914 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12709 1151 1727 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12708 1151 2728 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12707 vdd 1169 1151 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12706 4051 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12705 4051 2830 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12704 vdd 5069 4051 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12703 1559 2799 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12702 1559 2830 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12701 vdd 5069 1559 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12700 vdd 6440 1559 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12699 2010 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12698 2306 2512 2010 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12697 vdd 2314 2306 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12696 1594 1888 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12695 1627 2304 1594 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12694 vdd 1884 1627 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12693 5937 6375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12692 5937 6374 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12691 vdd 6423 5937 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12690 vdd 5936 5937 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12689 vdd 3757 3554 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12688 3554 3553 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12687 vdd 3953 3554 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12686 3552 3554 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12685 vdd 6364 6367 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12684 6367 6363 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12683 vdd 6632 6367 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12682 6362 6367 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12681 vdd 4948 4949 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12680 4949 4946 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12679 vdd 4947 4949 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12678 4945 4949 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12677 2530 5725 2434 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12676 2434 3186 2530 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12675 vdd 2758 2434 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12674 1909 2044 1912 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12673 1910 2046 1909 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12672 vdd 2045 1910 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12671 5721 1912 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12670 3198 3199 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12669 3197 3618 3198 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12668 vdd 5958 3197 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12667 1984 1986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12666 vdd 4509 1984 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12665 1985 1984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12664 869 4524 2352 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12663 868 4748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12662 vdd 868 869 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12661 vdd 4153 4154 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12660 4154 4150 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12659 vdd 6118 4154 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12658 4151 4154 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12657 vdd 1372 1373 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12656 1373 2506 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12655 vdd 1985 1373 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12654 3042 1373 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12653 vdd 5524 5012 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12652 5012 5914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12651 5012 5670 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12650 vdd 6665 5012 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12649 5014 5012 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12648 4068 3664 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12647 4068 3866 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12646 vdd 3849 4068 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12645 5979 6434 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12644 vdd 6919 5979 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12643 6186 5979 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12642 2760 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12641 vdd 4441 2760 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12640 2952 2760 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12639 vdd 488 219 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12638 489 784 220 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12637 220 488 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12636 220 219 489 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12635 vdd 218 220 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12634 218 784 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12633 1179 1332 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12632 vdd 1177 1179 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12631 1178 1179 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12630 6492 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12629 vdd 6492 6490 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12628 6489 6726 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12627 vdd 6489 6309 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12626 6309 6490 6487 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12625 6487 6492 6308 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12624 6307 6480 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12623 vdd 6483 6480 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12622 6480 6483 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12621 6308 6484 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12620 6484 6487 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12619 vdd 6976 6484 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12618 6483 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12617 6483 6490 6307 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12616 6484 6492 6483 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12615 3363 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12614 vdd 3363 3364 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12613 3362 3640 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12612 vdd 3362 3278 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12611 3278 3364 3360 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12610 3360 3363 3277 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12609 3298 4239 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12608 vdd 3445 4239 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12607 4239 3445 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12606 3277 3358 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12605 3358 3360 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12604 vdd 6976 3358 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12603 3445 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12602 3445 3364 3298 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12601 3358 3363 3445 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12600 3590 3776 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12599 vdd 3589 3590 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12598 3591 3590 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12597 2509 2508 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12596 vdd 2507 2509 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12595 3566 2509 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12594 vdd 2125 1766 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12593 1766 1991 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12592 1766 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12591 vdd 5363 1766 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12590 2180 1766 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12589 2988 3610 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12588 vdd 2987 2988 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12587 2986 2988 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12586 2008 3167 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12585 2097 2495 2008 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12584 vdd 2111 2097 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12583 6577 6579 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12582 6572 6578 6573 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12581 vdd 6905 6572 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12580 6575 6578 6577 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12579 6576 6582 6575 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12578 vdd 6574 6576 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12577 6574 6575 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12576 6573 6582 6574 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12575 vdd 6573 6905 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12574 6905 6573 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12573 vdd 6580 6582 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12572 6578 6582 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12571 vdd 6589 6579 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12570 vdd 6705 6241 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12569 6241 6690 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12568 6241 6951 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12567 vdd 6703 6241 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12566 6959 6241 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12565 vdd 640 600 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12564 600 1513 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12563 vdd 2314 600 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12562 598 600 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12561 6747 6915 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12560 6745 6916 6908 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12559 vdd 6906 6745 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12558 6912 6916 6747 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12557 6746 6918 6912 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12556 vdd 6909 6746 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12555 6909 6912 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12554 6908 6918 6909 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12553 vdd 6908 6906 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12552 6906 6908 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12551 vdd 6984 6918 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12550 6916 6918 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12549 vdd 6914 6915 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12548 vdd 6590 6318 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12547 6792 6581 6267 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12546 6267 6590 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12545 6267 6318 6792 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12544 vdd 6315 6267 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12543 6315 6581 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12542 6305 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12541 6475 6473 6305 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12540 vdd 6471 6475 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12539 2416 4088 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12538 vdd 3849 2416 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12537 2415 2416 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12536 vdd 3593 1691 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12535 1691 1688 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12534 vdd 2347 1691 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12533 1687 1691 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12532 4389 4391 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12531 4385 4392 4386 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12530 vdd 5026 4385 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12529 4390 4392 4389 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12528 4388 4393 4390 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12527 vdd 4387 4388 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12526 4387 4390 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12525 4386 4393 4387 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12524 vdd 4386 5026 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12523 5026 4386 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12522 vdd 6580 4393 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12521 4392 4393 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12520 vdd 4395 4391 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12519 1202 1205 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12518 1197 1204 1198 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12517 vdd 3790 1197 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12516 1200 1204 1202 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12515 1201 1206 1200 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12514 vdd 1199 1201 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12513 1199 1200 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12512 1198 1206 1199 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12511 vdd 1198 3790 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12510 3790 1198 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12509 vdd 3259 1206 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12508 1204 1206 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12507 vdd 1203 1205 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12506 5257 5723 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12505 5681 5721 5257 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12504 vdd 5927 5681 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12503 vdd 6839 6840 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12502 6847 6835 6764 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12501 6764 6839 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12500 6764 6840 6847 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12499 vdd 6836 6764 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12498 6836 6835 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12497 4983 5062 5490 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12496 5063 5065 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12495 vdd 5063 4983 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12494 5431 5258 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12493 vdd 5444 5431 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12492 5263 5264 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12491 vdd 5262 5263 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12490 584 2086 562 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12489 562 586 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12488 vdd 946 562 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12487 1312 584 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12486 561 588 584 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12485 562 774 561 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12484 5405 5986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12483 5518 6214 5405 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12482 vdd 6874 5518 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12481 vdd 4616 4717 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12480 4717 6951 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12479 4717 4613 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12478 vdd 5772 4717 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12477 4722 4717 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12476 6304 6469 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12475 6470 6713 6304 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12474 6303 6715 6470 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12473 vdd 6962 6303 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12472 6704 6470 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12471 274 319 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12470 323 320 274 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12469 vdd 328 323 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12468 3606 5737 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12467 vdd 3608 3606 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12466 3618 5116 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12465 vdd 3218 3618 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12464 2294 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_12463 2723 2291 2294 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_12462 2293 2304 2723 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_12461 vdd 2292 2293 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_12460 6174 6172 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12459 6398 6173 6174 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12458 vdd 6188 6398 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12457 899 2793 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12456 vdd 1002 898 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12455 vdd 1004 1008 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12454 1006 1004 899 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12453 898 1008 1006 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12452 1001 1006 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12451 896 2741 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12450 vdd 1191 895 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12449 vdd 1004 994 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12448 992 1004 896 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12447 895 994 992 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12446 990 992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12445 280 2048 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12444 vdd 1182 279 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12443 vdd 1004 352 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12442 353 1004 280 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12441 279 352 353 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12440 350 353 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12439 175 914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12438 vdd 633 174 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12437 vdd 1004 223 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12436 221 1004 175 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12435 174 223 221 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12434 222 221 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12433 5965 4453 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12432 vdd 4472 5965 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12431 5948 5116 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12430 vdd 3617 5948 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12429 4665 4862 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12428 vdd 4587 4665 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12427 4273 3866 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12426 4273 4942 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12425 vdd 4089 4273 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12424 vdd 3836 4273 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12423 2086 2161 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12422 vdd 1900 2086 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12421 4153 3946 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12420 4153 3947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12419 vdd 6423 4153 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12418 3284 3401 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12417 vdd 3403 3285 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12416 vdd 3976 3402 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12415 3399 3976 3284 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12414 3285 3402 3399 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12413 3397 3399 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12412 2764 2763 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12411 vdd 3190 2761 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12410 vdd 3976 2765 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12409 2762 3976 2764 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12408 2761 2765 2762 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12407 2961 2762 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12406 2872 2981 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12405 vdd 2979 2871 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12404 vdd 3976 2984 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12403 2983 3976 2872 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12402 2871 2984 2983 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12401 2977 2983 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12400 185 2386 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12399 vdd 525 184 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12398 vdd 1004 256 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12397 253 1004 185 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12396 184 256 253 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12395 255 253 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12394 6713 6974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12393 6713 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12392 vdd 6952 6713 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12391 vdd 6963 6713 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12390 481 480 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_12389 961 477 481 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_12388 479 478 961 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_12387 vdd 482 479 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_12386 vdd 2308 2289 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12385 2291 2298 2290 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12384 2290 2308 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12383 2290 2289 2291 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12382 vdd 2288 2290 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12381 2288 2298 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12380 878 1289 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12379 947 1158 878 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12378 vdd 946 947 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12377 4217 4485 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12376 4217 6600 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12375 vdd 4220 4217 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12374 vdd 5259 5260 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12373 5260 5263 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12372 vdd 5261 5260 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12371 5258 5260 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12370 847 849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12369 vdd 845 846 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12368 vdd 2394 850 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12367 848 2394 847 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12366 846 850 848 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12365 1563 848 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12364 2284 4241 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12363 vdd 4935 2283 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12362 vdd 4094 2395 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12361 2393 4094 2284 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12360 2283 2395 2393 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12359 2394 2393 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12358 vdd 6442 5893 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12357 vdd 6714 5892 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12356 5893 5892 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12355 6703 6963 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12354 6703 6917 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12353 vdd 6974 6703 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12352 vdd 4524 849 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12351 vdd 4748 538 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12350 849 538 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12349 3226 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12348 3226 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12347 vdd 3818 3226 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12346 vdd 6440 3226 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12345 4220 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12344 4220 5068 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12343 vdd 5069 4220 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12342 vdd 6440 4220 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12341 vdd 3391 1604 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12340 1604 2326 1665 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12339 1667 1665 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12338 2717 2727 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12337 2717 1877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12336 vdd 1875 2717 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12335 vdd 1876 2717 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12334 vdd 2919 2920 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12333 6172 2915 2882 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12332 2882 2919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12331 2882 2920 6172 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12330 vdd 2917 2882 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12329 2917 2915 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12328 vdd 5036 5038 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12327 5038 5041 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12326 vdd 5942 5038 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12325 5034 5038 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12324 4844 5017 4846 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12323 4846 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12322 vdd 6678 4846 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12321 4843 4844 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12320 4845 6637 4844 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12319 4846 5250 4845 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12318 vdd 4489 3808 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12317 3808 4042 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12316 3808 3813 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12315 vdd 4051 3808 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12314 4453 3808 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12313 vdd 86 68 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12312 1649 69 22 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12311 22 86 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12310 22 68 1649 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12309 vdd 71 22 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12308 71 69 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12307 1282 1287 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12306 vdd 1484 1282 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12305 1478 1282 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12304 2768 5953 2769 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12303 2769 2773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12302 vdd 4441 2769 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12301 2766 2768 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12300 2767 3199 2768 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12299 2769 3618 2767 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12298 792 793 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12297 vdd 791 792 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12296 973 792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12295 1160 1320 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12294 vdd 2314 1160 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12293 1298 1160 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12292 vdd 6116 5251 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12291 5250 5524 5249 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12290 5249 6116 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12289 5249 5251 5250 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12288 vdd 5248 5249 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12287 5248 5524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12286 1769 3263 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12285 vdd 3460 1769 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12284 2400 1769 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12283 4221 4220 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12282 vdd 4485 4221 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12281 4472 4221 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12280 vdd 4524 1590 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12279 1590 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12278 1590 4299 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12277 vdd 5363 1590 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12276 2412 1590 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12275 4882 4880 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12274 5708 4881 4882 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12273 vdd 5948 5708 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12272 1141 1144 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12271 1137 1143 1138 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12270 vdd 3382 1137 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12269 1142 1143 1141 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12268 1140 1145 1142 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12267 vdd 1139 1140 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12266 1139 1142 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12265 1138 1145 1139 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12264 vdd 1138 3382 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12263 3382 1138 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12262 vdd 3160 1145 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12261 1143 1145 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12260 vdd 3315 1144 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12259 617 3188 568 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12258 568 1904 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12257 vdd 3217 568 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12256 615 617 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12255 567 2746 617 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12254 568 1322 567 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12253 vdd 1521 1520 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12252 1520 1527 1669 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12251 3628 4942 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12250 vdd 4941 3628 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12249 4053 3628 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12248 vdd 4088 1983 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12247 1983 4501 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12246 vdd 3460 1983 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12245 1982 1983 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12244 vdd 2728 2480 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12243 2480 2727 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12242 vdd 2723 2480 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12241 2720 2480 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12240 556 674 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12239 554 675 669 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12238 vdd 829 554 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12237 673 675 556 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12236 555 676 673 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12235 vdd 670 555 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12234 670 673 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12233 669 676 670 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12232 vdd 669 829 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12231 829 669 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12230 vdd 3259 676 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12229 675 676 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12228 vdd 828 674 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12227 vdd 5954 5282 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12226 5282 5502 6374 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12225 4487 4737 4486 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12224 4486 4485 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12223 vdd 4488 4487 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12222 5342 4487 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12221 vdd 3226 2783 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12220 2783 2788 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12219 2783 4220 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12218 vdd 4485 2783 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12217 2782 2783 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12216 vdd 6917 6215 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12215 6215 6974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12214 vdd 6963 6215 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12213 6214 6215 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12212 1272 1580 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12211 1379 1749 1272 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12210 vdd 4748 1379 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12209 vdd 6870 6860 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12208 6858 6874 6767 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12207 6767 6870 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12206 6767 6860 6858 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12205 vdd 6856 6767 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12204 6856 6874 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12203 2776 5993 2779 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12202 2777 2775 2776 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12201 vdd 5967 2777 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12200 3603 3600 3602 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12199 3601 3783 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12198 vdd 3601 3603 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12197 2942 3738 2863 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12196 2863 3737 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12195 vdd 5272 2942 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12194 2950 2942 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12193 4891 5721 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12192 5104 5723 4891 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12191 vdd 5964 5104 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12190 3318 3549 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12189 vdd 3317 3318 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12188 9 112 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12187 7 40 107 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12186 vdd 504 7 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12185 39 40 9 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12184 8 111 39 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12183 vdd 37 8 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12182 37 39 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12181 107 111 37 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12180 vdd 107 504 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12179 504 107 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12178 vdd 3259 111 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12177 40 111 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12176 vdd 239 112 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12175 vdd 6725 6729 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12174 6729 6728 6730 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12173 6726 6730 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12172 2785 2998 2786 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12171 2786 4220 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12170 vdd 5116 2786 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12169 4483 2785 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12168 2784 2999 2785 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12167 2786 2997 2784 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12166 1300 1313 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12165 vdd 961 1300 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12164 6491 5533 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12163 vdd 5531 6491 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12162 3548 3714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12161 vdd 3558 3548 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12160 399 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12159 399 402 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12158 vdd 863 399 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12157 1949 2057 1948 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12156 1950 2155 1949 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12155 1949 2135 1950 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12154 1948 1947 1949 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12153 1948 2360 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12152 vdd 1946 1948 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12151 5925 6665 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12150 5925 6910 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12149 vdd 6806 5925 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12148 5788 5792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12147 vdd 5789 5788 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12146 vdd 6966 6772 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12145 6772 6968 6969 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12144 6967 6969 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12143 6970 6951 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12142 6970 6707 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12141 vdd 6705 6970 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12140 6951 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12139 vdd 6917 6951 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12138 5401 5730 5498 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12137 5497 5508 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12136 vdd 5497 5401 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12135 4446 4447 4679 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12134 4445 4444 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12133 vdd 4445 4446 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12132 6363 6375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12131 6363 6374 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12130 vdd 6423 6363 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12129 vdd 6165 6363 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12128 2346 2344 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12127 vdd 2345 2346 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12126 3617 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12125 3617 5748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12124 vdd 5749 3617 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12123 4616 5341 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12122 vdd 5992 4616 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12121 1554 1749 1555 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12120 1555 1580 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12119 vdd 4275 1554 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12118 2521 1554 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12117 2333 3186 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12116 vdd 6187 2333 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12115 1947 2138 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12114 1947 2139 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12113 vdd 1945 1947 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12112 6634 6855 6635 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12111 6635 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12110 vdd 6678 6635 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12109 6632 6634 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12108 6633 6637 6634 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12107 6635 6858 6633 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12106 4490 4496 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12105 vdd 4489 4490 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12104 4488 4490 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12103 2887 3792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12102 2996 3793 2887 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12101 vdd 3423 2996 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12100 494 629 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12099 494 3195 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12098 vdd 641 494 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12097 vdd 3217 494 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12096 1744 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12095 1744 2352 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12094 vdd 4937 1744 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12093 1562 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12092 1562 2125 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12091 vdd 1576 1562 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12090 2173 2389 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12089 2173 2170 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12088 vdd 2392 2173 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12087 1194 851 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12086 1194 844 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12085 vdd 3813 1194 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12084 vdd 3226 1194 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12083 911 1171 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12082 vdd 1727 911 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12081 vdd 2924 2725 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12080 3174 2723 2726 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12079 2726 2924 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12078 2726 2725 3174 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12077 vdd 2724 2726 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12076 2724 2723 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12075 4884 4886 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12074 vdd 4883 4884 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12073 5702 4884 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12072 5041 6375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12071 5041 6374 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12070 vdd 6423 5041 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12069 vdd 5039 5041 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12068 vdd 6186 4443 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12067 4443 6431 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12066 4444 4441 4443 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12065 4442 6220 4444 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12064 4443 5300 4442 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12063 vdd 6167 6168 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12062 6168 6360 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12061 vdd 6371 6168 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12060 6166 6168 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12059 vdd 5029 4864 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12058 4864 4866 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12057 vdd 4863 4864 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12056 4862 4864 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12055 3304 3453 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12054 3652 3451 3304 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12053 vdd 3452 3652 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12052 2520 2562 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12051 2520 3004 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12050 vdd 2165 2520 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12049 vdd 2157 2520 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12048 vdd 6186 5281 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12047 5281 6431 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12046 5279 6187 5281 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12045 5280 5954 5279 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12044 5281 5502 5280 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12043 1519 1517 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12042 vdd 1518 1519 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12041 3401 1519 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12040 976 980 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12039 vdd 975 976 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12038 1328 976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12037 271 335 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12036 314 310 271 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12035 vdd 607 314 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12034 4133 4275 4225 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12033 4131 4224 4133 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12032 4132 4708 4131 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12031 vdd 6224 4132 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12030 4929 4225 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12029 1916 2535 2046 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12028 1917 2521 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12027 vdd 1917 1916 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12026 vdd 6448 5785 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12025 5785 6917 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12024 vdd 6682 5785 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12023 6014 5785 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12022 460 581 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12021 vdd 1169 460 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12020 569 460 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12019 1915 1913 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12018 vdd 1914 1915 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12017 2044 1915 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12016 134 133 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12015 vdd 2387 134 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12014 987 134 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12013 1894 2495 1895 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12012 1895 3167 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12011 vdd 2111 1894 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12010 1893 1894 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12009 764 941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12008 vdd 947 764 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12007 770 764 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12006 2287 2286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12005 vdd 2895 2287 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12004 2716 2287 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12003 vdd 1945 1941 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12002 1941 2154 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12001 vdd 2122 1941 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12000 2050 1941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11999 2884 2950 2951 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11998 2949 2953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11997 vdd 2949 2884 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11996 vdd 494 337 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11995 337 784 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11994 vdd 2314 337 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11993 335 337 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11992 883 973 1172 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11991 974 1178 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11990 vdd 974 883 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11989 1896 2161 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11988 vdd 1900 1896 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11987 2106 1896 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11986 1739 1967 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11985 vdd 1758 1739 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11984 1737 1739 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11983 2094 2485 2007 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11982 2007 2095 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11981 vdd 2102 2007 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11980 2092 2094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11979 2006 2319 2094 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11978 2007 2320 2006 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11977 3164 5723 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11976 3317 5721 3164 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11975 vdd 3969 3317 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11974 6733 6787 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11973 6731 6789 6781 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11972 vdd 6807 6731 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11971 6784 6789 6733 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11970 6732 6790 6784 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11969 vdd 6783 6732 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11968 6783 6784 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11967 6781 6790 6783 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11966 vdd 6781 6807 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11965 6807 6781 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11964 vdd 6832 6790 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11963 6789 6790 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11962 vdd 6786 6787 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11961 5713 5716 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11960 5710 5717 5709 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11959 vdd 5953 5710 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11958 5714 5717 5713 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11957 5712 5718 5714 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11956 vdd 5711 5712 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11955 5711 5714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11954 5709 5718 5711 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11953 vdd 5709 5953 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11952 5953 5709 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11951 vdd 6832 5718 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11950 5717 5718 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11949 vdd 5715 5716 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11948 vdd 5748 5137 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11947 5137 5749 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11946 vdd 6440 5137 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11945 5133 5137 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11944 vdd 3226 3214 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11943 3214 4220 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11942 vdd 4485 3214 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11941 3424 3214 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11940 vdd 6186 5726 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11939 5726 6431 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11938 6167 5725 5726 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11937 5724 6182 6167 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11936 5726 6183 5724 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11935 854 1035 855 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11934 855 863 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11933 vdd 1038 854 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11932 1004 854 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11931 547 648 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11930 545 650 643 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11929 vdd 3796 545 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11928 646 650 547 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11927 546 651 646 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11926 vdd 645 546 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11925 645 646 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11924 643 651 645 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11923 vdd 643 3796 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11922 3796 643 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11921 vdd 3160 651 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11920 650 651 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11919 vdd 652 648 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11918 4713 5748 4574 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11917 vdd 4715 4574 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11916 4574 5545 4713 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11915 6188 4713 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11914 2998 2553 2025 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11913 2025 2521 2998 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11912 vdd 2520 2025 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11911 2025 2534 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11910 3406 3414 3286 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11909 3286 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11908 vdd 5243 3406 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11907 3404 3406 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11906 vdd 4088 4090 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11905 4090 4091 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11904 4090 4089 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11903 vdd 4087 4090 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11902 5889 4090 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11901 vdd 4491 3053 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11900 3053 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11899 vdd 4524 3053 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11898 3051 3053 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11897 5682 5680 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11896 vdd 5681 5682 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11895 vdd 1309 1311 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11894 4673 1306 1248 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11893 1248 1309 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11892 1248 1311 4673 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11891 vdd 1308 1248 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11890 1308 1306 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11889 2832 3456 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11888 5069 3457 2832 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11887 vdd 3455 5069 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11886 vdd 1737 1496 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11885 1496 2506 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11884 1632 1882 1496 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11883 1495 1885 1632 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11882 1496 1891 1495 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11881 5436 5264 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11880 vdd 5372 5436 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11879 3179 3178 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11878 vdd 3395 3176 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11877 vdd 3976 3180 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11876 3177 3976 3179 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11875 3176 3180 3177 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11874 3337 3177 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11873 6108 6422 6210 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11872 6109 6420 6108 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11871 vdd 6421 6109 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11870 6211 6210 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11869 6795 6877 6734 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11868 6734 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11867 vdd 6807 6795 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11866 6794 6795 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11865 195 470 197 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11864 197 1900 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11863 vdd 2161 197 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11862 302 195 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11861 194 598 195 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11860 197 307 194 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11859 3615 3792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11858 3616 3793 3615 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11857 vdd 3802 3616 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11856 3969 3814 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11855 3969 5115 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11854 vdd 3816 3969 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11853 3679 3761 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11852 vdd 3759 3678 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11851 vdd 3976 3762 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11850 3764 3976 3679 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11849 3678 3762 3764 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11848 3758 3764 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11847 3543 3570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11846 vdd 3972 3542 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11845 vdd 3976 3569 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11844 3568 3976 3543 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11843 3542 3569 3568 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11842 3750 3568 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11841 3978 3975 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11840 vdd 3979 3973 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11839 vdd 3976 3977 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11838 3974 3976 3978 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11837 3973 3977 3974 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11836 3986 3974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11835 3541 3566 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11834 vdd 3573 3540 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11833 vdd 3976 3567 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11832 3564 3976 3541 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11831 3540 3567 3564 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11830 3565 3564 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11829 4410 4414 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11828 vdd 4175 4410 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11827 603 2314 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11826 603 640 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11825 vdd 1317 603 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11824 4920 5756 4922 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11823 4922 5805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11822 vdd 4918 4920 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11821 4919 4920 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11820 2058 3006 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11819 vdd 3010 2058 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11818 4007 4213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11817 4009 4212 4007 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11816 vdd 4897 4009 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11815 vdd 6434 3677 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11814 3677 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11813 3757 5243 3677 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11812 3676 4217 3757 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11811 3677 5502 3676 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11810 vdd 6226 5741 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11809 5741 6426 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11808 6205 5804 5741 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11807 5740 6182 6205 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11806 5741 6183 5740 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11805 1136 1196 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11804 vdd 3790 1135 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11803 vdd 2797 1195 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11802 1193 2797 1136 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11801 1135 1195 1193 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11800 1203 1193 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11799 901 1208 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11798 vdd 3423 900 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11797 vdd 2797 1012 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11796 1011 2797 901 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11795 900 1012 1011 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11794 1007 1011 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11793 4860 6877 4861 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11792 4861 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11791 vdd 4914 4860 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11790 4859 4860 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11789 6611 6839 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11788 vdd 6850 6611 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11787 6814 6611 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11786 476 2314 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11785 476 640 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11784 vdd 1513 476 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11783 640 3217 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11782 640 2544 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11781 vdd 2142 640 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11780 69 772 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11779 vdd 1151 69 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11778 4048 3816 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11777 vdd 3814 4048 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11776 4285 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11775 4285 4287 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11774 vdd 4941 4285 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11773 vdd 4524 4285 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11772 2116 2740 2015 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11771 2015 2520 2116 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11770 vdd 2117 2015 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11769 5829 6191 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11768 6748 6190 5829 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11767 vdd 5964 6748 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11766 vdd 5975 5977 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11765 5977 6209 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11764 vdd 5973 5977 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11763 5972 5977 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11762 1212 1953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11761 1212 845 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11760 vdd 2194 1212 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11759 vdd 3836 1212 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11758 4485 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11757 4485 2807 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11756 vdd 5069 4485 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11755 vdd 6440 4485 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11754 2343 2535 2342 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11753 2341 2349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11752 vdd 2341 2343 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11751 vdd 2744 2743 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11750 2743 2940 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11749 vdd 2938 2743 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11748 2742 2743 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11747 778 776 777 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11746 777 1300 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11745 vdd 870 778 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11744 1163 778 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11743 vdd 5157 2285 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11742 2285 4299 2417 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11741 2418 2417 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11740 vdd 2080 2079 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11739 2919 2895 2000 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11738 2000 2080 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11737 2000 2079 2919 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11736 vdd 2081 2000 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11735 2081 2895 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11734 vdd 6885 6646 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11733 6646 6874 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11732 6646 6893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11731 vdd 6906 6646 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11730 6839 6646 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11729 1701 2553 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11728 vdd 2534 1701 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11727 1700 1701 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11726 1267 1580 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11725 1356 1749 1267 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11724 vdd 4275 1356 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11723 1889 2299 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11722 vdd 2492 1889 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11721 1888 1889 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11720 vdd 6116 6113 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11719 6115 6112 6117 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11718 6117 6116 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11717 6117 6113 6115 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11716 vdd 6114 6117 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11715 6114 6112 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11714 2756 5725 2757 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11713 vdd 2758 2757 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11712 2757 3186 2756 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11711 2755 2756 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11710 2941 2940 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11709 vdd 2938 2941 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11708 3975 2941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11707 5414 5749 5559 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11706 5560 5784 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11705 vdd 5560 5414 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11704 3630 4942 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11703 vdd 3658 3630 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11702 5068 3630 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11701 2334 2349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11700 vdd 2512 2334 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11699 2519 2334 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11698 2709 2711 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11697 2704 2710 2705 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11696 vdd 3546 2704 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11695 2708 2710 2709 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11694 2706 2713 2708 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11693 vdd 2707 2706 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11692 2707 2708 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11691 2705 2713 2707 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11690 vdd 2705 3546 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11689 3546 2705 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11688 vdd 3160 2713 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11687 2710 2713 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11686 vdd 3318 2711 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11685 vdd 4265 4264 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11684 4264 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11683 vdd 6440 4264 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11682 4492 4264 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11681 vdd 4062 3623 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11680 3623 5068 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11679 vdd 5069 3623 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11678 3798 3623 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11677 3643 3658 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11676 vdd 4286 3643 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11675 3818 3643 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11674 vdd 2498 1497 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11673 1497 2161 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11672 vdd 1900 1497 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11671 1640 1497 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11670 1275 2409 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11669 1389 2198 1275 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11668 vdd 1587 1389 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11667 2013 2106 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11666 5993 2107 2013 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11665 vdd 2109 5993 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11664 vdd 5936 5732 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11663 5732 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11662 5732 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11661 vdd 6440 5732 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11660 5735 5732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11659 1499 2736 1502 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11658 1502 2498 1500 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11657 1500 2106 1502 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11656 1499 2535 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11655 vdd 3217 1499 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11654 1502 2111 1499 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11653 1498 1500 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11652 18 132 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11651 16 55 126 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11650 vdd 527 16 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11649 54 55 18 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11648 17 131 54 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11647 vdd 52 17 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11646 52 54 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11645 126 131 52 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11644 vdd 126 527 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11643 527 126 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11642 vdd 3259 131 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11641 55 131 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11640 vdd 258 132 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11639 5399 5954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11638 5727 5502 5399 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11637 vdd 5804 5727 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11636 5318 5986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11635 5320 6214 5318 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11634 vdd 6885 5320 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11633 vdd 3866 1980 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11632 1980 2352 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11631 1980 3849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11630 vdd 3664 1980 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11629 2399 1980 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11628 vdd 4477 3223 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11627 3224 5987 3225 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11626 3222 3221 3224 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11625 3223 4456 3222 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11624 2891 3245 2890 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11623 3044 6727 2891 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11622 2891 3046 3044 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11621 2890 3042 2891 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11620 2890 3248 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11619 vdd 4748 2890 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11618 232 234 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11617 227 233 228 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11616 vdd 500 227 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11615 231 233 232 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11614 230 235 231 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11613 vdd 229 230 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11612 229 231 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11611 228 235 229 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11610 vdd 228 500 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11609 500 228 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11608 vdd 3160 235 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11607 233 235 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11606 vdd 237 234 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11605 vdd 6186 5833 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11604 5834 6420 6806 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11603 5835 6222 5834 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11602 5833 6422 5835 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11601 6697 6935 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11600 6930 6696 6697 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11599 vdd 6706 6930 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11598 3685 4213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11597 3781 4212 3685 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11596 vdd 4438 3781 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11595 4553 5954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11594 4682 5502 4553 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11593 vdd 5953 4682 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11592 3712 3950 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11591 vdd 3725 3712 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11590 6192 6190 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11589 6203 6191 6192 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11588 vdd 6188 6203 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11587 2821 2820 2822 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11586 2822 3040 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11585 vdd 3238 2821 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11584 2824 2821 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11583 5392 5949 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11582 5444 5947 5392 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11581 vdd 5927 5444 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11580 6705 6480 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11579 6705 6448 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11578 vdd 6917 6705 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11577 4990 5986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11576 5097 6214 4990 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11575 vdd 6740 5097 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11574 1561 1989 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11573 3793 1745 1561 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11572 vdd 1560 3793 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11571 2886 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11570 2987 3414 2886 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11569 vdd 6265 2987 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11568 1620 2921 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11567 1620 2896 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11566 vdd 2897 1620 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11565 3949 4151 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11564 vdd 3948 3949 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11563 5729 5728 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11562 vdd 5727 5729 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11561 6170 5729 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11560 6798 6905 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11559 6798 6910 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11558 vdd 6806 6798 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11557 6808 6807 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11556 6808 6910 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11555 vdd 6806 6808 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11554 5791 5907 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11553 vdd 6440 5791 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11552 6701 6917 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11551 6701 6449 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11550 vdd 6448 6701 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11549 6702 6682 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11548 6702 6448 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11547 vdd 6917 6702 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11546 586 591 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11545 vdd 589 586 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11544 4613 5341 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11543 vdd 5575 4613 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11542 1171 1209 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11541 vdd 1876 1171 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11540 1883 2095 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11539 1883 1882 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11538 vdd 2088 1883 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11537 1976 1975 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11536 vdd 2400 1976 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11535 3221 1976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11534 vdd 4675 4415 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11533 4415 4865 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11532 vdd 4668 4415 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11531 4414 4415 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11530 1509 2946 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11529 1508 2950 1509 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11528 vdd 2111 1508 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11527 vdd 2924 2925 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11526 6190 2921 2883 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11525 2883 2924 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11524 2883 2925 6190 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11523 vdd 2922 2883 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11522 2922 2921 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11521 vdd 5953 5822 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11520 5822 5954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11519 5867 6867 5822 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11518 5821 5951 5867 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11517 5822 5952 5821 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11516 vdd 6616 6320 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11515 6320 6591 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11514 vdd 6807 6320 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11513 6778 6320 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11512 202 607 203 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11511 203 1900 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11510 vdd 2161 203 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11509 200 202 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11508 201 335 202 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11507 203 310 201 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11506 3035 3259 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11505 vdd 3035 3036 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11504 3034 3039 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11503 vdd 3034 2877 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11502 2877 3036 3032 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11501 3032 3035 2876 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11500 2875 4937 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11499 vdd 3029 4937 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11498 4937 3029 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11497 2876 3030 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11496 3030 3032 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11495 vdd 6976 3030 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11494 3029 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11493 3029 3036 2875 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11492 3030 3035 3029 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11491 4559 6220 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11490 4903 5300 4559 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11489 vdd 4696 4903 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11488 5812 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11487 5915 6877 5812 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11486 vdd 6905 5915 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11485 vdd 1662 1516 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11484 1516 1517 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11483 vdd 1518 1516 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11482 1695 1516 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11481 6002 6440 5846 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11480 5846 6691 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11479 vdd 6921 5846 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11478 6182 6002 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11477 5845 5999 6002 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11476 5846 6000 5845 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11475 3597 4213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11474 3598 4212 3597 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11473 vdd 4205 3598 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11472 1905 2375 1906 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11471 1906 1904 1905 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11470 vdd 2382 1906 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11469 3684 3775 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11468 3682 3774 3769 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11467 vdd 5963 3682 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11466 3772 3774 3684 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11465 3683 3777 3772 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11464 vdd 3770 3683 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11463 3770 3772 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11462 3769 3777 3770 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11461 vdd 3769 5963 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11460 5963 3769 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11459 vdd 5054 3777 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11458 3774 3777 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11457 vdd 4200 3775 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11456 vdd 3598 3599 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11455 3599 5737 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11454 vdd 3608 3599 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11453 3596 3599 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11452 1386 2400 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11451 vdd 1395 1386 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11450 1385 1386 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11449 5546 5545 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11448 vdd 5748 5546 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11447 5544 5546 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11446 vdd 2407 1981 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11445 1981 2125 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11444 1981 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11443 vdd 3664 1981 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11442 1979 1981 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11441 2207 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11440 2207 1991 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11439 vdd 2125 2207 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11438 vdd 5363 2207 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11437 1994 2418 1993 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11436 1993 2629 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11435 vdd 2208 1994 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11434 1992 1994 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11433 1887 2299 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11432 vdd 2489 1887 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11431 1885 1887 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11430 952 1171 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11429 vdd 1727 952 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11428 2727 952 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11427 2496 3186 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11426 vdd 5963 2496 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11425 2495 2496 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11424 2443 2999 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11423 5125 2997 2443 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11422 vdd 2998 5125 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11421 4565 5753 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11420 4703 5767 4565 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11419 vdd 4914 4703 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11418 vdd 3602 2547 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11417 2547 2545 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11416 vdd 2546 2547 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11415 2544 2547 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11414 2953 5953 2885 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11413 2885 3186 2953 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11412 vdd 2952 2885 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11411 5554 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11410 vdd 5575 5554 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11409 5999 5554 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11408 vdd 3263 2613 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11407 2613 5157 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11406 vdd 5363 2613 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11405 2807 2613 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11404 2198 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11403 2198 2125 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11402 vdd 2407 2198 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11401 vdd 3664 2198 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11400 5760 5766 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11399 vdd 5758 5760 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11398 5759 5760 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11397 2014 2116 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11396 2109 2514 2014 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11395 vdd 2323 2109 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11394 vdd 1877 1878 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11393 1878 2727 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11392 vdd 1876 1878 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11391 2080 1878 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11390 1036 1039 909 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11389 909 6469 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11388 vdd 1578 1036 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11387 1035 1036 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11386 3999 3998 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11385 3994 4000 3993 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11384 vdd 5725 3994 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11383 3997 4000 3999 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11382 3996 4001 3997 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11381 vdd 3995 3996 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11380 3995 3997 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11379 3993 4001 3995 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11378 vdd 3993 5725 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11377 5725 3993 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11376 vdd 5054 4001 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11375 4000 4001 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11374 vdd 4002 3998 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11373 193 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11372 576 191 193 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11371 192 322 576 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11370 vdd 200 192 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11369 vdd 5501 5298 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11368 5298 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11367 5298 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11366 vdd 6440 5298 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11365 5297 5298 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11364 3188 5958 3189 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11363 3189 3186 3188 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11362 vdd 3187 3189 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11361 vdd 3227 3011 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11360 3011 5116 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11359 vdd 3218 3011 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11358 3006 3011 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11357 vdd 3831 3437 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11356 3437 3629 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11355 3437 4253 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11354 vdd 3827 3437 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11353 3438 3437 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11352 3392 5372 3282 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11351 3282 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11350 vdd 4897 3282 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11349 3391 3392 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11348 3281 3737 3392 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11347 3282 3738 3281 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11346 512 515 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11345 508 514 509 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11344 vdd 3607 508 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11343 513 514 512 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11342 511 516 513 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11341 vdd 510 511 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11340 510 513 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11339 509 516 510 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11338 vdd 509 3607 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11337 3607 509 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11336 vdd 3259 516 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11335 514 516 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11334 vdd 657 515 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11333 4991 5112 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11332 5319 5113 4991 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11331 vdd 5134 5319 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11330 vdd 4941 4943 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11329 4943 4942 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11328 4943 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11327 vdd 6440 4943 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11326 5545 4943 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11325 vdd 4094 3704 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11324 3704 4748 4287 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11323 5857 5918 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11322 vdd 5856 5857 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11321 5919 5264 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11320 vdd 5902 5919 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11319 vdd 6225 5415 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11318 5415 5567 5566 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11317 5573 5566 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11316 vdd 1309 1161 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11315 2138 1163 1164 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11314 1164 1309 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11313 1164 1161 2138 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11312 vdd 1162 1164 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11311 1162 1163 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11310 4913 5756 4912 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11309 4912 5805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11308 vdd 5026 4913 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11307 4911 4913 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11306 1673 2122 1606 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11305 1606 2124 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11304 vdd 2125 1606 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11303 1913 1673 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11302 1605 1682 1673 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11301 1606 1911 1605 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11300 vdd 3458 3306 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11299 3306 3863 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11298 3453 3455 3306 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11297 3305 3456 3453 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11296 3306 3457 3305 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11295 4138 5112 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11294 4462 5113 4138 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11293 vdd 4241 4462 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11292 1233 3263 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11291 vdd 3460 1233 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11290 1237 1239 1238 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11289 1238 1588 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11288 vdd 1576 1237 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11287 1236 1237 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11286 2441 3199 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11285 2550 3618 2441 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11284 vdd 5804 2550 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11283 2433 2749 2940 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11282 2432 2750 2433 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11281 vdd 2752 2432 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11280 2445 2741 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11279 vdd 3421 2444 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11278 vdd 2797 2565 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11277 2564 2797 2445 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11276 2444 2565 2564 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11275 2560 2564 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11274 1538 2048 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11273 vdd 3604 1537 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11272 vdd 2797 1540 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11271 1539 2797 1538 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11270 1537 1540 1539 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11269 1549 1539 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11268 551 914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11267 vdd 3607 550 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11266 vdd 2797 662 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11265 660 2797 551 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11264 550 662 660 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11263 657 660 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11262 549 917 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11261 vdd 3796 548 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11260 vdd 2797 656 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11259 654 2797 549 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11258 548 656 654 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11257 652 654 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11256 5585 5528 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11255 vdd 5978 5585 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11254 986 3021 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11253 986 395 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11252 vdd 686 986 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11251 558 2386 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11250 vdd 3434 557 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11249 vdd 2797 681 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11248 679 2797 558 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11247 557 681 679 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11246 677 679 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11245 2795 2793 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11244 vdd 3802 2796 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11243 vdd 2797 2798 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11242 2794 2797 2795 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11241 2796 2798 2794 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11240 2792 2794 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11239 3661 3663 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11238 vdd 3660 3661 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11237 3662 3661 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11236 6677 6877 6679 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11235 6679 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11234 vdd 6893 6677 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11233 6676 6677 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11232 4479 4572 4481 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11231 4480 4709 4479 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11230 4478 5548 4480 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11229 vdd 4477 4478 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11228 4612 4481 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11227 vdd 3606 3211 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11226 3211 3212 3213 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11225 3210 3213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11224 3636 4726 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11223 vdd 5575 3636 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11222 2040 4941 2039 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11221 2039 4089 2204 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11220 2204 2412 2039 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11219 2040 2411 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11218 vdd 2615 2040 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11217 2039 2415 2040 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11216 2202 2204 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11215 2329 2740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11214 2329 2331 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11213 vdd 2520 2329 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11212 vdd 2336 2278 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11211 2278 2342 2335 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11210 2750 2335 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11209 vdd 6184 6181 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11208 6181 6390 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11207 vdd 6869 6181 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11206 6180 6181 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11205 2450 5125 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11204 vdd 2583 2449 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11203 vdd 2587 2588 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11202 2586 2587 2450 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11201 2449 2588 2586 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11200 2582 2586 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11199 vdd 6919 6131 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11198 6131 6434 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11197 6129 6867 6131 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11196 6130 6128 6129 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11195 6131 6127 6130 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11194 2454 2823 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11193 2601 2600 2454 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11192 vdd 2817 2601 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11191 179 914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11190 vdd 500 178 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11189 vdd 830 238 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11188 236 830 179 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11187 178 238 236 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11186 237 236 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11185 181 917 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11184 vdd 504 180 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11183 vdd 830 241 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11182 240 830 181 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11181 180 241 240 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11180 239 240 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11179 553 1196 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11178 vdd 663 552 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11177 vdd 830 667 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11176 666 830 553 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11175 552 667 666 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11174 661 666 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11173 183 1208 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11172 vdd 392 182 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11171 vdd 830 244 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11170 242 830 183 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11169 182 244 242 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11168 243 242 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11167 6260 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11166 vdd 6260 6259 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11165 6257 6256 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11164 vdd 6257 6258 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11163 6258 6259 6254 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11162 6254 6260 6255 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11161 6251 6263 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11160 vdd 6252 6263 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11159 6263 6252 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11158 6255 6253 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11157 6253 6254 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11156 vdd 6976 6253 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11155 6252 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11154 6252 6259 6251 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11153 6253 6260 6252 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11152 vdd 4732 4736 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11151 4736 4618 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11150 4736 5115 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11149 vdd 5552 4736 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11148 4948 4736 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11147 1572 3836 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11146 1572 2194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11145 vdd 1953 1572 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11144 vdd 6440 1572 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11143 575 573 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11142 vdd 571 575 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11141 776 575 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11140 4086 4089 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11139 4086 4091 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11138 vdd 4088 4086 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11137 vdd 4087 4086 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11136 2888 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11135 3003 3414 2888 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11134 vdd 6727 3003 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11133 4134 4524 4232 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11132 4135 6224 4134 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11131 vdd 4708 4135 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11130 4470 4232 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11129 vdd 5068 4208 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11128 4208 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11127 4208 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11126 vdd 4308 4208 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11125 4689 4208 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11124 vdd 3849 3665 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11123 3665 3866 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11122 3665 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11121 vdd 3664 3665 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11120 3663 3665 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11119 4029 4275 4031 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11118 4030 4028 4029 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11117 4027 4708 4030 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11116 vdd 6224 4027 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11115 5321 4031 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11114 1269 4748 1553 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11113 1359 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11112 vdd 1359 1269 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11111 2189 3229 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11110 vdd 4501 2189 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11109 2188 2189 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11108 4871 4874 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11107 4867 4875 4868 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11106 vdd 5039 4867 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11105 4872 4875 4871 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11104 4870 4877 4872 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11103 vdd 4869 4870 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11102 4869 4872 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11101 4868 4877 4869 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11100 vdd 4868 5039 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11099 5039 4868 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11098 vdd 5054 4877 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11097 4875 4877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11096 vdd 4873 4874 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11095 vdd 1558 1557 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11094 1557 1968 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11093 vdd 1559 1557 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11092 1724 1557 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11091 vdd 2553 2147 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11090 2147 2356 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11089 vdd 2331 2147 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11088 2146 2147 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11087 vdd 3781 3780 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11086 3780 4909 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11085 vdd 3788 3780 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11084 3776 3780 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11083 623 1737 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11082 vdd 2506 623 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11081 2498 623 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11080 4136 5112 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11079 4238 5113 4136 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11078 vdd 4235 4238 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11077 3235 3233 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11076 vdd 3234 3235 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11075 3231 3235 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11074 vdd 3866 1384 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11073 1384 3849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11072 vdd 3664 1384 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11071 1965 1384 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11070 vdd 5745 3611 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11069 3611 3616 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11068 vdd 4018 3611 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11067 3610 3611 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11066 vdd 1972 1974 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11065 1974 1973 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11064 vdd 3442 1974 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11063 1971 1974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11062 3270 3375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11061 3268 3313 3373 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11060 vdd 3547 3268 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11059 3312 3313 3270 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11058 3269 3314 3312 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11057 vdd 3310 3269 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11056 3310 3312 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11055 3373 3314 3310 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11054 vdd 3373 3547 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11053 3547 3373 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11052 vdd 6580 3314 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11051 3313 3314 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11050 vdd 3548 3375 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11049 vdd 1988 1987 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11048 1987 1989 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11047 vdd 1990 1987 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11046 2623 1987 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11045 2734 2944 2735 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11044 2735 3572 2734 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11043 vdd 2733 2735 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11042 vdd 5069 2800 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11041 2800 2830 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11040 2800 2799 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11039 vdd 6440 2800 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11038 3414 2800 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11037 3955 4157 3956 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11036 3956 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11035 vdd 6678 3956 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11034 3953 3955 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11033 3954 6637 3955 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11032 3956 4643 3954 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11031 250 252 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11030 245 251 246 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11029 vdd 522 245 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11028 249 251 250 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11027 247 254 249 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11026 vdd 248 247 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11025 248 249 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11024 246 254 248 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11023 vdd 246 522 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11022 522 246 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11021 vdd 3259 254 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11020 251 254 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11019 vdd 387 252 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11018 1532 3210 1531 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11017 1531 1534 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11016 vdd 2349 1532 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11015 1530 1532 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11014 vdd 6974 5847 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11013 5847 6963 6448 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11012 4678 6600 4552 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11011 4552 4676 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11010 vdd 6601 4678 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11009 4675 4678 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11008 5023 6877 4974 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11007 4974 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11006 vdd 5670 5023 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11005 5022 5023 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11004 5416 5791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11003 5800 5792 5416 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11002 vdd 5573 5800 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11001 4129 4213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11000 4215 4212 4129 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10999 vdd 4687 4215 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10998 vdd 6242 4077 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10997 4078 4083 4520 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10996 4076 4075 4078 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10995 4077 4082 4076 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10994 283 361 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10993 281 362 355 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10992 vdd 502 281 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10991 358 362 283 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10990 282 363 358 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10989 vdd 357 282 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10988 357 358 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10987 355 363 357 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10986 vdd 355 502 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10985 502 355 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10984 vdd 3160 363 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10983 362 363 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10982 vdd 364 361 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10981 6683 6682 6684 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10980 6681 6934 6683 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10979 vdd 6694 6681 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10978 6680 6684 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10977 2349 1968 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10976 vdd 1559 2349 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10975 2002 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10974 2085 2291 2002 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10973 2001 2292 2085 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10972 vdd 2304 2001 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10971 2921 2085 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10970 1886 2303 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10969 1886 1884 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10968 vdd 2092 1886 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10967 4013 4452 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10966 vdd 4051 4013 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10965 5264 5116 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10964 5264 5329 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10963 vdd 5552 5264 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10962 589 1652 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10961 vdd 1508 589 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10960 vdd 6974 6962 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10959 vdd 6963 6965 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10958 6962 6965 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10957 1973 2399 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10956 vdd 1757 1973 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10955 1972 1975 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10954 vdd 1234 1972 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10953 3605 3792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10952 4010 3793 3605 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10951 vdd 3604 4010 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10950 1491 1498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10949 1491 1490 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10948 vdd 1635 1491 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10947 1484 1482 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10946 1484 1627 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10945 vdd 1483 1484 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10944 vdd 2518 2430 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10943 2431 2519 3184 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10942 2429 2536 2431 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10941 2430 2522 2429 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10940 1278 1989 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_10939 1565 1745 1278 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_10938 1279 6469 1565 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_10937 vdd 2787 1279 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_10936 6177 6375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10935 6177 6374 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10934 vdd 6423 6177 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10933 vdd 6522 6177 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10932 2820 2604 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10931 2820 3242 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10930 vdd 2603 2820 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10929 3186 4485 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10928 3186 3226 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10927 vdd 4220 3186 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10926 5772 6917 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10925 vdd 6963 5772 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10924 1357 1749 1268 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10923 1268 1580 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10922 vdd 4524 1357 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10921 2534 1357 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10920 933 1169 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10919 933 941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10918 vdd 947 933 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10917 2286 1876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10916 2286 1877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10915 vdd 2727 2286 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10914 vdd 5932 5934 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10913 5934 6347 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10912 vdd 5937 5934 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10911 5931 5934 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10910 vdd 6176 6179 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10909 6179 6177 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10908 vdd 6393 6179 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10907 6175 6179 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10906 vdd 6226 5302 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10905 5302 6426 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10904 5493 5299 5302 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10903 5301 6220 5493 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10902 5302 5300 5301 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10901 3021 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10900 3021 3023 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10899 vdd 5068 3021 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10898 1587 3849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10897 1587 2125 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10896 vdd 3866 1587 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10895 vdd 3664 1587 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10894 vdd 6434 3681 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10893 3681 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10892 3766 4308 3681 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10891 3680 4217 3766 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10890 3681 5502 3680 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10889 vdd 3856 3857 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10888 3857 3853 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10887 vdd 4524 3857 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10886 4075 3857 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10885 vdd 5877 5751 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10884 5751 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10883 vdd 6440 5751 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10882 6183 5751 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10881 6006 6238 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10880 vdd 6440 6006 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10879 6004 6006 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10878 1613 2058 1729 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10877 1611 1740 1613 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10876 1612 1728 1611 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10875 vdd 1727 1612 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10874 2156 1729 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10873 791 624 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10872 791 794 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10871 vdd 3193 791 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10870 vdd 625 791 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10869 1578 3849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10868 1578 2352 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10867 vdd 3866 1578 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10866 vdd 3664 1578 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10865 1951 2381 1952 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10864 1952 2379 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10863 vdd 4748 1951 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10862 2350 1951 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10861 939 1156 875 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10860 875 1146 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10859 vdd 2086 939 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10858 938 939 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10857 5460 5699 5395 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10856 5395 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10855 vdd 6678 5395 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10854 5456 5460 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10853 5394 6637 5460 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10852 5395 5695 5394 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10851 2398 2603 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10850 vdd 2604 2398 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10849 2823 2398 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10848 2554 2553 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10847 vdd 2951 2554 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10846 2551 2554 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10845 2133 2344 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10844 vdd 2345 2133 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10843 2129 2133 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10842 4578 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10841 4744 5992 4578 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10840 vdd 5889 4744 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10839 4060 4275 4061 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10838 4057 4059 4060 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10837 4058 4708 4057 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10836 vdd 6224 4058 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10835 5538 4061 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10834 1600 2111 1599 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10833 1645 2106 1600 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10832 1600 2498 1645 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10831 1599 2736 1600 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10830 1599 2535 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10829 vdd 3217 1599 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10828 3804 5068 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10827 vdd 5069 3804 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10826 3805 3804 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10825 2330 2353 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10824 vdd 2329 2330 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10823 2517 2330 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10822 5289 5288 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10821 5284 5290 5283 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10820 vdd 5804 5284 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10819 5286 5290 5289 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10818 5287 5291 5286 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10817 vdd 5285 5287 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10816 5285 5286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10815 5283 5291 5285 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10814 vdd 5283 5804 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10813 5804 5283 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10812 vdd 6832 5291 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10811 5290 5291 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10810 vdd 5292 5288 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10809 vdd 5914 4384 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10808 4839 6665 4383 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10807 4383 5914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10806 4383 4384 4839 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10805 vdd 4382 4383 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10804 4382 6665 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10803 vdd 6702 6240 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10802 6240 6701 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10801 6240 6704 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10800 vdd 6700 6240 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10799 6957 6240 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10798 vdd 2396 2179 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10797 2179 2074 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10796 2179 2070 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10795 vdd 2506 2179 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10794 2603 2179 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10793 vdd 4703 4227 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10792 4227 4228 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10791 4227 4925 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10790 vdd 4238 4227 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10789 4226 4227 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10788 4573 4708 4709 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10787 4710 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10786 vdd 4710 4573 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10785 3013 3816 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10784 vdd 3814 3013 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10783 3010 3013 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10782 vdd 4726 4729 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10781 4729 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10780 vdd 6440 4729 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10779 4725 4729 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10778 1986 5359 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10777 1986 2407 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10776 vdd 2406 1986 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10775 vdd 3836 1986 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10774 vdd 3263 1757 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10773 vdd 3460 1759 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10772 1757 1759 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10771 1481 1480 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10770 1479 1478 1481 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10769 vdd 1620 1479 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10768 4433 4436 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10767 4428 4435 4429 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10766 vdd 5959 4428 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10765 4432 4435 4433 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10764 4431 4437 4432 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10763 vdd 4430 4431 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10762 4430 4432 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10761 4429 4437 4430 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10760 vdd 4429 5959 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10759 5959 4429 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10758 vdd 5054 4437 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10757 4435 4437 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10756 vdd 4434 4436 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10755 vdd 4658 4657 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10754 4857 4853 4549 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10753 4549 4658 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10752 4549 4657 4857 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10751 vdd 4659 4549 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10750 4659 4853 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10749 6223 6224 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10748 6222 6221 6223 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10747 vdd 6702 6222 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10746 vdd 493 492 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10745 492 615 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10744 vdd 2314 492 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10743 491 492 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10742 vdd 4726 4718 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10741 4718 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10740 vdd 6440 4718 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10739 4715 4718 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10738 vdd 3369 3251 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10737 3251 3371 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10736 3451 3455 3251 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10735 3250 3456 3451 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10734 3251 3457 3250 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10733 5108 5341 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10732 vdd 5575 5108 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10731 5986 5108 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10730 vdd 5993 3584 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10729 3584 5967 3761 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10728 4012 4213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10727 4016 4212 4012 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10726 vdd 5064 4016 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10725 5393 5949 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10724 5859 5947 5393 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10723 vdd 5965 5859 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10722 1547 1550 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10721 1543 1551 1544 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10720 vdd 3604 1543 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10719 1548 1551 1547 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10718 1546 1552 1548 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10717 vdd 1545 1546 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10716 1545 1548 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10715 1544 1552 1545 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10714 vdd 1544 3604 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10713 3604 1544 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10712 vdd 3259 1552 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10711 1551 1552 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10710 vdd 1549 1550 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10709 1253 1328 1517 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10708 1327 1326 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10707 vdd 1327 1253 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10706 vdd 1313 960 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10705 1518 961 880 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10704 880 1313 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10703 880 960 1518 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10702 vdd 962 880 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10701 962 961 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10700 vdd 5345 4508 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10699 4508 4507 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10698 vdd 4505 4508 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10697 4506 4508 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10696 vdd 4276 2616 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10695 2616 4089 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10694 2616 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10693 vdd 3866 2616 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10692 4491 2616 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10691 5907 5893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10690 6471 6728 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10689 6226 6480 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10688 6025 6261 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10687 vdd 6571 5997 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10686 5997 5889 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10685 5997 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10684 vdd 6440 5997 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10683 5998 5997 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10682 vdd 6434 4125 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10681 4125 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10680 4171 6265 4125 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10679 4124 4217 4171 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10678 4125 5502 4124 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10677 vdd 2999 955 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10676 1309 953 879 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10675 879 2999 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10674 879 955 1309 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10673 vdd 956 879 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10672 956 953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10671 3689 3792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10670 3788 3793 3689 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10669 vdd 3796 3788 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10668 6023 6263 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10667 vdd 5157 3657 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10666 3657 4299 3658 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10665 2338 2737 2749 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10664 2337 2535 2338 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10663 vdd 2355 2337 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10662 6610 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10661 6609 6877 6610 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10660 vdd 6820 6609 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10659 261 3229 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10658 vdd 845 261 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10657 839 841 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10656 835 842 836 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10655 vdd 3423 835 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10654 840 842 839 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10653 838 843 840 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10652 vdd 837 838 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10651 837 840 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10650 836 843 837 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10649 vdd 836 3423 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10648 3423 836 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10647 vdd 3259 843 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10646 842 843 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10645 vdd 1007 841 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10644 5485 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10643 5485 6431 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10642 vdd 6434 5485 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10641 6589 6593 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10640 vdd 6588 6589 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10639 6597 6600 6599 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10638 6599 6598 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10637 vdd 6601 6597 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10636 6596 6597 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10635 6690 6691 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10634 vdd 6921 6690 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10633 507 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10632 2545 987 507 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10631 vdd 663 2545 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10630 972 1322 882 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10629 882 4176 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10628 vdd 2747 972 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10627 981 972 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10626 1596 1885 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10625 1635 1891 1596 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10624 vdd 1882 1635 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10623 5278 5279 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10622 vdd 5277 5278 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10621 6364 5278 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10620 6647 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10619 6648 6877 6647 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10618 vdd 6885 6648 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10617 269 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10616 303 305 269 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10615 268 302 303 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10614 vdd 312 268 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10613 301 303 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10612 332 2314 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10611 332 494 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10610 vdd 784 332 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10609 2741 2940 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10608 vdd 2938 2741 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10607 3199 3814 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10606 3199 3631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10605 vdd 3816 3199 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10604 263 4501 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10603 263 1732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10602 vdd 1231 263 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10601 503 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10600 1688 987 503 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10599 vdd 502 1688 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10598 vdd 6814 6608 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10597 6607 6820 6606 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10596 6606 6814 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10595 6606 6608 6607 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10594 vdd 6605 6606 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10593 6605 6820 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10592 3990 4217 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10591 3991 5502 3990 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10590 vdd 6727 3991 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10589 3220 3225 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10588 vdd 3438 3220 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10587 3976 3220 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10586 4898 5300 4900 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10585 4900 6220 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10584 vdd 4897 4898 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10583 4896 4898 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10582 5246 5914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10581 vdd 6665 5246 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10580 5245 5246 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10579 2408 3062 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10578 2408 2207 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10577 vdd 2198 2408 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10576 vdd 3060 2408 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10575 2840 4094 4087 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10574 2841 5363 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10573 vdd 2841 2840 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10572 vdd 5299 3672 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10571 3672 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10570 3741 6265 3672 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10569 3671 3737 3741 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10568 3672 3738 3671 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10567 vdd 1298 1153 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10566 1490 1647 1155 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10565 1155 1298 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10564 1155 1153 1490 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10563 vdd 1154 1155 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10562 1154 1647 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10561 5373 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10560 vdd 5373 5371 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10559 5370 5369 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10558 vdd 5370 5368 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10557 5368 5371 5367 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10556 5367 5373 5366 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10555 5362 5363 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10554 vdd 5364 5363 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10553 5363 5364 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10552 5366 5365 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10551 5365 5367 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10550 vdd 6976 5365 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10549 5364 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10548 5364 5371 5362 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10547 5365 5373 5364 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10546 4123 5044 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10545 4394 5045 4123 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10544 vdd 5927 4394 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10543 vdd 6691 6227 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10542 6227 6226 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10541 vdd 6921 6227 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10540 6225 6227 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10539 1266 1580 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10538 1353 1749 1266 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10537 vdd 4524 1353 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10536 vdd 2520 2276 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10535 2276 2740 2322 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10534 2323 2322 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10533 vdd 4878 4879 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10532 4879 5269 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10531 vdd 5456 4879 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10530 4876 4879 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10529 2825 2823 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10528 2826 5792 2825 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10527 vdd 2824 2826 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10526 908 1033 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10525 2607 1223 908 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10524 vdd 1732 2607 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10523 vdd 1572 1220 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10522 1220 1381 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10521 1220 1367 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10520 vdd 2070 1220 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10519 2797 1220 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10518 vdd 4453 4454 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10517 4454 4460 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10516 4454 4455 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10515 vdd 4472 4454 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10514 6375 4454 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10513 966 968 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10512 vdd 965 966 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10511 3178 966 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10510 vdd 3217 788 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10509 788 1904 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10508 787 3188 788 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10507 786 2746 787 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10506 788 1322 786 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10505 5817 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10504 5943 6877 5817 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10503 vdd 6740 5943 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10502 4970 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10501 5011 6877 4970 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10500 vdd 6665 5011 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10499 vdd 579 462 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10498 462 2727 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10497 vdd 1876 462 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10496 466 462 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10495 3232 5773 3230 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10494 3233 5575 3232 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10493 3232 4726 3233 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10492 3230 4053 3232 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10491 3230 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10490 vdd 3229 3230 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10489 3296 3634 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10488 5964 3632 3296 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10487 vdd 3442 5964 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10486 1228 2194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10485 1745 2195 1228 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10484 vdd 6440 1745 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10483 5382 5455 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10482 5380 5454 5448 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10481 vdd 5501 5380 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10480 5452 5454 5382 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10479 5381 5457 5452 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10478 vdd 5449 5381 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10477 5449 5452 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10476 5448 5457 5449 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10475 vdd 5448 5501 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10474 5501 5448 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10473 vdd 6832 5457 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10472 5454 5457 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10471 vdd 5453 5455 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10470 4126 4880 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10469 4175 4881 4126 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10468 vdd 5927 4175 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10467 vdd 6714 6438 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10466 6438 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10465 6438 6952 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10464 vdd 6963 6438 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10463 6691 6438 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10462 2177 2399 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10461 vdd 2799 2177 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10460 2174 2177 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10459 3007 3429 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10458 vdd 3003 3007 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10457 3004 3007 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10456 vdd 6186 4440 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10455 4440 6431 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10454 4685 4438 4440 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10453 4439 6220 4685 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10452 4440 5300 4439 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10451 3148 3149 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10450 3143 3150 3144 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10449 vdd 3709 3143 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10448 3147 3150 3148 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10447 3146 3151 3147 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10446 vdd 3145 3146 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10445 3145 3147 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10444 3144 3151 3145 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10443 vdd 3144 3709 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10442 3709 3144 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10441 vdd 3160 3151 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10440 3150 3151 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10439 vdd 3712 3149 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10438 vdd 3217 2164 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10437 2164 3006 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10436 vdd 3010 2164 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10435 2161 2164 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10434 3959 3962 3960 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10433 3960 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10432 vdd 6678 3960 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10431 3957 3959 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10430 3958 6637 3959 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10429 3960 4160 3958 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10428 vdd 4942 4934 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10427 4934 4941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10426 vdd 5773 4934 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10425 5756 4934 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10424 vdd 4286 3835 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10423 3835 4941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10422 3835 3836 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10421 vdd 4524 3835 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10420 4250 3835 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10419 vdd 1953 1954 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10418 1954 2194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10417 1954 2125 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10416 vdd 3836 1954 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10415 2514 1954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10414 5861 5931 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10413 vdd 5859 5861 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10412 5744 5967 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10411 6417 5993 5744 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10410 vdd 5948 6417 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10409 4427 4673 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10408 5270 4671 4427 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10407 vdd 5948 5270 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10406 291 385 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10405 289 384 379 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10404 vdd 825 289 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10403 382 384 291 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10402 290 386 382 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10401 vdd 380 290 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10400 380 382 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10399 379 386 380 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10398 vdd 379 825 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10397 825 379 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10396 vdd 3259 386 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10395 384 386 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10394 vdd 517 385 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10393 6479 6477 6306 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10392 6306 6974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10391 vdd 6480 6479 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10390 6725 6479 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10389 4561 4695 4604 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10388 4560 5089 4561 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10387 vdd 4919 4560 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10386 1334 3408 1256 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10385 1256 1340 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10384 vdd 2534 1334 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10383 1333 1334 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10382 4969 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10381 5008 6877 4969 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10380 vdd 5670 5008 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10379 vdd 2188 2032 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10378 2033 4213 2074 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10377 2031 2174 2033 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10376 2032 3051 2031 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10375 vdd 3263 1616 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10374 1616 3460 1778 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10373 4589 4876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10372 vdd 4672 4589 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10371 3970 4673 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10370 3971 4671 3970 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10369 vdd 3969 3971 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10368 5815 6172 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10367 6143 6173 5815 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10366 vdd 5965 6143 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10365 1336 3408 1257 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10364 1257 1340 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10363 vdd 2349 1336 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10362 1338 1336 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10361 3659 3660 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10360 vdd 4087 3659 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10359 3856 3659 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10358 1728 1559 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10357 1728 1558 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10356 vdd 1968 1728 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10355 2136 2544 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10354 vdd 2142 2136 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10353 3655 3652 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10352 3655 3654 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10351 vdd 3653 3655 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10350 1758 5359 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10349 1758 2412 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10348 vdd 2406 1758 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10347 vdd 4501 1758 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10346 6988 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10345 vdd 6988 6986 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10344 6985 6981 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10343 vdd 6985 6758 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10342 6758 6986 6982 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10341 6982 6988 6757 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10340 6756 6974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10339 vdd 6978 6974 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10338 6974 6978 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10337 6757 6979 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10336 6979 6982 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10335 vdd 6976 6979 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10334 6978 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10333 6978 6986 6756 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10332 6979 6988 6978 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10331 vdd 5014 4647 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10330 4647 4918 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10329 vdd 5026 4647 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10328 4658 4647 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10327 4236 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10326 vdd 4233 4236 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10325 6422 4236 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10324 1661 2375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10323 1661 1737 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10322 vdd 1904 1661 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10321 vdd 2755 2019 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10320 2019 3586 2121 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10319 2135 2121 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10318 2587 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10317 2587 2807 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10316 vdd 5069 2587 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10315 vdd 5363 2629 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10314 vdd 3263 2078 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10313 2629 2078 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10312 2111 2501 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10311 2111 2506 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10310 vdd 3217 2111 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10309 vdd 2782 2111 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10308 2099 2512 2009 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10307 2009 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10306 vdd 2314 2099 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10305 2299 2099 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10304 3239 4083 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10303 3238 4082 3239 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10302 vdd 6265 3238 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10301 vdd 6596 6595 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10300 6595 6594 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10299 vdd 6798 6595 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10298 6593 6595 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10297 2403 5157 2404 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10296 2402 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10295 vdd 2402 2403 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10294 3559 6172 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10293 3558 6173 3559 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10292 vdd 3969 3558 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10291 vdd 5068 4902 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10290 4902 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10289 4902 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10288 vdd 5902 4902 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10287 5062 4902 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10286 6468 6694 6302 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10285 6302 6466 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10284 vdd 6476 6302 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10283 6463 6468 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10282 6301 6464 6468 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10281 6302 6690 6301 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10280 958 1313 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10279 vdd 961 958 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10278 1165 958 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10277 2414 2415 2413 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10276 2622 2412 2414 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10275 2414 4089 2622 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10274 2413 4941 2414 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10273 2413 2411 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10272 vdd 2615 2413 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10271 1148 1485 1147 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10270 1147 1488 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10269 vdd 1490 1148 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10268 1146 1148 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10267 4426 4880 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10266 4591 4881 4426 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10265 vdd 5965 4591 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10264 1614 1735 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10263 1959 1950 1614 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10262 vdd 2801 1959 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10261 vdd 6959 6961 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10260 6961 6957 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10259 vdd 6974 6961 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10258 6972 6961 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10257 vdd 1229 1042 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10256 1042 1039 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10255 vdd 1038 1042 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10254 2604 1042 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10253 1343 2544 1261 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10252 1261 2142 1343 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10251 vdd 1353 1261 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10250 1017 1214 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10249 vdd 1215 1017 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10248 1210 1017 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10247 683 859 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10246 vdd 682 683 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10245 844 683 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10244 1283 1292 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10243 vdd 1491 1283 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10242 1480 1283 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10241 6626 6877 6625 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10240 6625 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10239 vdd 6740 6626 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10238 6624 6626 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10237 4959 4962 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10236 4956 4964 4955 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10235 vdd 5359 4956 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10234 4960 4964 4959 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10233 4958 4963 4960 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10232 vdd 4957 4958 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10231 4957 4960 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10230 4955 4963 4957 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10229 vdd 4955 5359 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10228 5359 4955 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10227 vdd 6984 4963 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10226 4964 4963 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10225 vdd 4961 4962 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10224 4988 5080 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10223 4986 5082 5075 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10222 vdd 5742 4986 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10221 5077 5082 4988 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10220 4987 5081 5077 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10219 vdd 5076 4987 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10218 5076 5077 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10217 5075 5081 5076 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10216 vdd 5075 5742 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10215 5742 5075 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10214 vdd 6984 5081 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10213 5082 5081 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10212 vdd 5306 5080 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10211 6284 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10210 6640 6877 6284 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10209 vdd 6893 6640 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10208 vdd 5914 5909 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10207 6128 5910 5811 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10206 5811 5914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10205 5811 5909 6128 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10204 vdd 5912 5811 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10203 5912 5910 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10202 4509 2406 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10201 4509 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10200 vdd 3866 4509 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10199 vdd 3836 4509 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10198 1222 1221 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10197 vdd 1224 1222 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10196 1365 1222 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10195 1902 2375 1903 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10194 vdd 2382 1903 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10193 1903 1904 1902 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10192 2319 1902 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10191 vdd 5064 3173 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10190 3173 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10189 3172 5902 3173 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10188 3171 3737 3172 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10187 3173 3738 3171 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10186 vdd 6893 6645 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10185 6644 6906 6643 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10184 6643 6893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10183 6643 6645 6644 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10182 vdd 6642 6643 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10181 6642 6906 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10180 vdd 5749 5090 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10179 5090 5748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10178 5090 6740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10177 vdd 6440 5090 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10176 5089 5090 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10175 2405 2404 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10174 vdd 2407 2405 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10173 2830 2405 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10172 vdd 936 763 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10171 763 1479 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10170 vdd 933 763 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10169 769 763 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10168 4980 5053 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10167 4978 5055 5048 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10166 vdd 5958 4978 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10165 5050 5055 4980 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10164 4979 5056 5050 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10163 vdd 5049 4979 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10162 5049 5050 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10161 5048 5056 5049 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10160 vdd 5048 5958 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10159 5958 5048 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10158 vdd 5054 5056 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10157 5055 5056 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10156 vdd 5057 5053 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10155 vdd 4658 4652 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10154 4653 4914 4548 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10153 4548 4658 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10152 4548 4652 4653 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10151 vdd 4655 4548 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10150 4655 4914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10149 4734 4733 4577 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10148 4577 6469 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10147 vdd 4731 4734 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10146 4732 4734 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10145 vdd 1313 768 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10144 5044 766 767 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10143 767 1313 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10142 767 768 5044 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10141 vdd 765 767 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10140 765 766 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10139 4514 4517 4515 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10138 4513 4622 4514 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10137 vdd 6000 4513 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10136 6447 5272 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10135 4676 4308 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10134 4176 5243 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10133 2746 5262 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10132 6598 6265 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10131 6603 6727 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10130 vdd 2852 2459 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10129 2459 3460 4089 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10128 3244 4083 3245 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10127 3243 3246 3244 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10126 vdd 4082 3243 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10125 2368 2370 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10124 2363 2369 2364 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10123 vdd 3421 2363 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10122 2367 2369 2368 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10121 2366 2372 2367 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10120 vdd 2365 2366 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10119 2365 2367 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10118 2364 2372 2365 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10117 vdd 2364 3421 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10116 3421 2364 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10115 vdd 3259 2372 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10114 2369 2372 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10113 vdd 2560 2370 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10112 2966 3160 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10111 vdd 2966 2965 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10110 2964 2961 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10109 vdd 2964 2867 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10108 2867 2965 2962 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10107 2962 2966 2866 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10106 2865 3190 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10105 vdd 2958 3190 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10104 3190 2958 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10103 2866 2959 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10102 2959 2962 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10101 vdd 6976 2959 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10100 2958 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10099 2958 2965 2865 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10098 2959 2966 2958 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10097 506 987 505 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10096 505 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10095 vdd 504 506 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10094 1189 506 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10093 4032 3423 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10092 5705 6591 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10091 4853 4914 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10090 3800 3790 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10089 2442 3199 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10088 2562 3618 2442 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10087 vdd 5742 2562 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10086 5410 5986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10085 5540 6214 5410 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10084 vdd 6906 5540 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10083 4522 4520 4630 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10082 4519 4521 4522 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10081 vdd 4518 4519 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10080 6786 6800 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10079 vdd 6132 6786 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10078 6220 6701 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10077 vdd 6702 6220 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10076 2896 1880 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10075 vdd 1883 2896 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10074 1875 2896 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10073 vdd 2897 1875 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10072 4851 6877 4852 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10071 4852 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10070 vdd 5026 4851 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10069 4850 4851 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10068 vdd 6970 6773 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10067 6773 6972 6971 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10066 6981 6971 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10065 vdd 1641 1639 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10064 1884 2097 1597 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10063 1597 1641 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10062 1597 1639 1884 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10061 vdd 1636 1597 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10060 1636 2097 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10059 2897 1632 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10058 vdd 1886 2897 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10057 vdd 6814 6816 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10056 6817 6811 6762 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10055 6762 6814 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10054 6762 6816 6817 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10053 vdd 6813 6762 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10052 6813 6811 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10051 vdd 6186 4557 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10050 4557 6431 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10049 4688 4687 4557 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10048 4556 6220 4688 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10047 4557 5300 4556 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10046 870 2727 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10045 870 579 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10044 vdd 576 870 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10043 vdd 1876 870 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10042 3411 3414 3290 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10041 3290 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10040 vdd 4308 3411 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10039 3600 3411 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10038 845 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10037 vdd 4748 845 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10036 3703 4094 4276 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10035 3858 4748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10034 vdd 3858 3703 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10033 2314 1900 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10032 2314 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10031 vdd 2161 2314 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10030 405 3460 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10029 405 2411 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10028 vdd 2615 405 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10027 682 4748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10026 682 1732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10025 vdd 1231 682 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10024 vdd 1298 1299 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10023 1483 1501 1246 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10022 1246 1298 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10021 1246 1299 1483 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10020 vdd 1295 1246 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10019 1295 1501 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10018 2525 2535 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10017 vdd 2737 2525 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10016 3992 4452 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10015 vdd 3991 3992 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10014 4150 3992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10013 vdd 6186 4985 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10012 4985 6685 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10011 5065 5064 4985 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10010 4984 6220 5065 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10009 4985 5300 4984 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10008 4484 4483 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10007 vdd 4482 4484 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10006 5154 4484 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10005 vdd 2852 1588 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10004 vdd 3460 1589 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10003 1588 1589 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10002 1990 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10001 1990 2352 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10000 vdd 1991 1990 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09999 vdd 5363 1990 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09998 1989 4087 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09997 1989 2352 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09996 vdd 4089 1989 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09995 vdd 4299 1989 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09994 5758 6906 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09993 5758 5545 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09992 vdd 5748 5758 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09991 vdd 5993 2282 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09990 2282 5967 2385 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09989 2386 2385 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09988 vdd 6405 6404 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09987 6404 6401 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09986 vdd 6660 6404 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09985 6400 6404 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09984 vdd m_clock 3419 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09983 5334 3419 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09982 vdd 3419 5334 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09981 vdd 3419 5334 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09980 5334 3419 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09979 vdd 5334 5335 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09978 6984 5335 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09977 vdd 5335 6984 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09976 vdd 5335 6984 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09975 6984 5335 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09974 vdd 5334 5333 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09973 5332 5333 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09972 vdd 5333 5332 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09971 vdd 5333 5332 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09970 5332 5333 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09969 vdd 5334 5122 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09968 5121 5122 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09967 vdd 5122 5121 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09966 vdd 5122 5121 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09965 5121 5122 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09964 vdd 5334 5267 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09963 6832 5267 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09962 vdd 5267 6832 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09961 vdd 5267 6832 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09960 6832 5267 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09959 vdd 5334 5266 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09958 6580 5266 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09957 vdd 5266 6580 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09956 vdd 5266 6580 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09955 6580 5266 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09954 886 918 978 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09953 884 3210 886 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09952 885 2537 884 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09951 vdd 919 885 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09950 1176 978 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09949 vdd 6974 6111 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09948 6111 6963 6218 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09947 6219 6218 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09946 vdd 4708 4576 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09945 4576 6224 4730 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09944 4731 4730 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09943 2731 2944 2732 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09942 vdd 2733 2732 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09941 2732 3572 2731 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09940 2730 2731 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09939 1184 1190 1183 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09938 1183 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09937 vdd 1182 1184 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09936 1919 1184 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09935 2513 2512 2016 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09934 2016 2511 2513 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09933 vdd 2117 2016 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09932 vdd 5068 4691 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09931 4691 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09930 4691 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09929 vdd 5243 4691 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09928 4692 4691 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09927 4977 5044 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09926 5864 5045 4977 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09925 vdd 6188 5864 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09924 vdd 1900 1242 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09923 1242 2161 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09922 1287 1490 1242 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09921 1241 1488 1287 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09920 1242 1485 1241 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09919 4046 4275 4047 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09918 4044 4043 4046 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09917 4045 4708 4044 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09916 vdd 6224 4045 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09915 5327 4047 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09914 vdd 6434 4128 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09913 4128 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09912 4181 5272 4128 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09911 4127 4217 4181 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09910 4128 5502 4127 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09909 5688 5690 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09908 5685 5691 5684 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09907 vdd 5936 5685 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09906 5689 5691 5688 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09905 5687 5692 5689 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09904 vdd 5686 5687 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09903 5686 5689 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09902 5684 5692 5686 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09901 vdd 5684 5936 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09900 5936 5684 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09899 vdd 6580 5692 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09898 5691 5692 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09897 vdd 5861 5690 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09896 4933 6422 6678 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09895 4932 4939 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09894 vdd 4932 4933 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09893 vdd 1953 692 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09892 692 2194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09891 692 3836 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09890 vdd 6440 692 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09889 690 692 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09888 1047 1991 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09887 vdd 1779 1047 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09886 1218 1047 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09885 139 405 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09884 vdd 4299 139 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09883 138 139 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09882 1615 1746 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09881 3792 1745 1615 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09880 vdd 2184 3792 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09879 6121 6123 6122 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09878 6122 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09877 vdd 6678 6122 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09876 6118 6121 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09875 6120 6637 6121 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09874 6122 6119 6120 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09873 vdd 6186 5828 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09872 5828 6685 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09871 6401 5963 5828 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09870 5827 6182 6401 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09869 5828 6183 5827 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09868 6639 6640 6641 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09867 6641 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09866 vdd 6678 6641 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09865 6636 6639 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09864 6638 6637 6639 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09863 6641 6644 6638 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09862 4055 4053 4056 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09861 4056 5575 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09860 vdd 4726 4056 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09859 5927 4055 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09858 4054 5992 4055 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09857 4056 5773 4054 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09856 vdd 5097 4464 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09855 4464 4463 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09854 4464 4701 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09853 vdd 4462 4464 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09852 4461 4464 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09851 vdd 1652 475 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09850 473 1505 474 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09849 474 1652 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09848 474 475 473 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09847 vdd 472 474 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09846 472 1505 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09845 vdd 1320 1159 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09844 1159 1647 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09843 vdd 2314 1159 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09842 1158 1159 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09841 2421 2467 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09840 2419 2468 2461 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09839 vdd 3946 2419 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09838 2465 2468 2421 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09837 2420 2469 2465 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09836 vdd 2463 2420 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09835 2463 2465 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09834 2461 2469 2463 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09833 vdd 2461 3946 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09832 3946 2461 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09831 vdd 3160 2469 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09830 2468 2469 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09829 vdd 3949 2467 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09828 vdd 4942 4067 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09827 4067 4941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09826 vdd 5349 4067 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09825 5749 4067 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09824 vdd 4276 3840 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09823 3840 4941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09822 3840 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09821 vdd 4524 3840 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09820 4726 3840 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09819 6 106 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09818 4 35 101 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09817 vdd 636 4 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09816 34 35 6 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09815 5 105 34 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09814 vdd 32 5 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09813 32 34 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09812 101 105 32 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09811 vdd 101 636 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09810 636 101 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09809 vdd 3160 105 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09808 35 105 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09807 vdd 225 106 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09806 771 911 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09805 772 769 771 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09804 vdd 770 772 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09803 1392 1394 1276 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09802 1276 1992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09801 vdd 2198 1392 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09800 1390 1392 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09799 1969 1982 1966 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09798 1967 5992 1969 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09797 1969 4053 1967 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09796 1966 1965 1969 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09795 1966 3229 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09794 vdd 2125 1966 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09793 2070 1732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09792 vdd 1223 2070 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09791 vdd 2299 2295 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09790 2298 2489 2297 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09789 2297 2299 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09788 2297 2295 2298 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09787 vdd 2296 2297 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09786 2296 2489 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09785 3340 5054 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09784 vdd 3340 3339 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09783 3338 3337 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09782 vdd 3338 3274 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09781 3274 3339 3335 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09780 3335 3340 3273 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09779 3280 3395 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09778 vdd 3388 3395 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09777 3395 3388 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09776 3273 3332 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09775 3332 3335 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09774 vdd 6976 3332 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09773 3388 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09772 3388 3339 3280 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09771 3332 3340 3388 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09770 6139 6362 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09769 vdd 5862 6139 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09768 3693 3798 3799 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09767 3692 4611 3693 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09766 vdd 3969 3692 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09765 3797 3799 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09764 vdd 6434 3968 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09763 3968 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09762 3967 5902 3968 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09761 3966 4217 3967 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09760 3968 5502 3966 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09759 vdd 6919 4973 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09758 4973 6434 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09757 5440 6867 4973 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09756 4972 5019 5440 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09755 4973 5022 4972 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09754 6706 6242 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09753 6706 6243 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09752 vdd 6476 6706 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09751 1536 3210 1535 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09750 1535 1534 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09749 vdd 2521 1536 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09748 1533 1536 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09747 2718 2915 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09746 2909 2716 2718 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09745 vdd 2717 2909 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09744 3458 5363 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09743 3458 3263 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09742 vdd 5157 3458 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09741 4873 5034 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09740 vdd 4591 4873 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09739 5955 6591 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09738 5955 6631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09737 vdd 6806 5955 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09736 5361 5359 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09735 5361 5570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09734 vdd 5788 5361 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09733 1277 1992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09732 1395 1394 1277 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09731 vdd 2198 1395 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09730 3448 3863 3300 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09729 3300 3455 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09728 vdd 3449 3300 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09727 3639 3448 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09726 3299 4071 3448 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09725 3300 3458 3299 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09724 1977 2180 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09723 3442 1979 1977 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09722 vdd 2193 3442 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09721 2355 3793 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09720 vdd 2352 2355 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09719 6371 6740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09718 6371 6631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09717 vdd 6806 6371 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09716 6372 6375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09715 6372 6374 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09714 vdd 6423 6372 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09713 vdd 6376 6372 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09712 6659 6893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09711 vdd 6906 6659 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09710 6890 6659 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09709 6420 4947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09708 6420 5549 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09707 vdd 4946 6420 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09706 1235 1233 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09705 1235 1975 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09704 vdd 1234 1235 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09703 773 1300 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09702 1306 776 773 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09701 vdd 870 1306 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09700 vdd 2346 2279 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09699 2279 2340 2339 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09698 4881 2339 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09697 66 310 21 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09696 21 335 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09695 vdd 607 66 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09694 307 66 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09693 3609 3792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09692 3608 3793 3609 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09691 vdd 3607 3608 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09690 1560 3836 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09689 1560 2194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09688 vdd 1953 1560 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09687 6687 6963 6919 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09686 6686 6974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09685 vdd 6686 6687 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09684 876 1146 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09683 941 1156 876 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09682 vdd 2086 941 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09681 vdd 6261 6021 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09680 6021 6023 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09679 vdd 6476 6021 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09678 6247 6021 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09677 1755 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09676 vdd 3866 1755 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09675 2183 1755 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09674 3065 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09673 vdd 5363 3065 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09672 3849 3065 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09671 2728 933 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09670 2728 936 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09669 vdd 1479 2728 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09668 2915 2723 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09667 2915 2728 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09666 vdd 2727 2915 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09665 vdd 5702 5703 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09664 5703 6342 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09663 vdd 5700 5703 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09662 5701 5703 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09661 vdd 4258 4249 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09660 4249 4253 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09659 vdd 4616 4249 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09658 4482 4249 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09657 vdd 1724 1725 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09656 1725 1722 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09655 vdd 1730 1725 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09654 2775 1725 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09653 2819 2820 2818 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09652 2818 3037 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09651 vdd 3236 2819 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09650 2817 2819 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09649 3192 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09648 vdd 4438 3192 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09647 3191 3192 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09646 1131 1188 1185 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09645 1132 3408 1131 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09644 1130 2770 1132 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09643 vdd 1189 1130 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09642 1186 1185 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09641 5752 5753 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09640 5761 5767 5752 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09639 vdd 6905 5761 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09638 5820 5949 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09637 6357 5947 5820 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09636 vdd 5948 6357 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09635 6462 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09634 vdd 6462 6461 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09633 6460 6463 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09632 vdd 6460 6300 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09631 6300 6461 6457 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09630 6457 6462 6299 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09629 6298 6694 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09628 vdd 6455 6694 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09627 6694 6455 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09626 6299 6456 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09625 6456 6457 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09624 vdd 6976 6456 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09623 6455 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09622 6455 6461 6298 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09621 6456 6462 6455 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09620 1170 1313 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09619 vdd 1169 1170 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09618 2999 1170 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09617 217 493 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09616 vdd 2314 217 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09615 216 217 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09614 3651 3649 3654 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09613 3650 4080 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09612 vdd 3650 3651 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09611 vdd 2406 1581 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09610 1581 2407 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09609 1581 5359 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09608 vdd 3836 1581 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09607 1580 1581 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09606 4995 5152 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09605 4993 5153 5146 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09604 vdd 5144 4993 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09603 5149 5153 4995 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09602 4994 5155 5149 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09601 vdd 5147 4994 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09600 5147 5149 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09599 5146 5155 5147 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09598 vdd 5146 5144 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09597 5144 5146 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09596 vdd 6984 5155 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09595 5153 5155 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09594 vdd 5151 5152 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09593 vdd 5014 4641 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09592 4643 5026 4547 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09591 4547 5014 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09590 4547 4641 4643 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09589 vdd 4642 4547 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09588 4642 5026 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09587 vdd 473 316 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09586 316 314 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09585 vdd 476 316 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09584 312 316 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09583 5105 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09582 vdd 6440 5105 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09581 5102 5105 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09580 2789 3617 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09579 vdd 2787 2789 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09578 2788 2789 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09577 696 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09576 vdd 4748 696 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09575 857 696 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09574 3025 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09573 vdd 6440 3025 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09572 3023 3025 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09571 3822 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09570 vdd 3818 3822 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09569 3819 3822 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09568 2439 3199 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09567 2542 3618 2439 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09566 vdd 5963 2542 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09565 vdd 4892 4893 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09564 4893 4899 5478 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09563 3708 3874 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09562 3706 3873 3868 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09561 vdd 4094 3706 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09560 3870 3873 3708 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09559 3707 3875 3870 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09558 vdd 3869 3707 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09557 3869 3870 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09556 3868 3875 3869 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09555 vdd 3868 4094 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09554 4094 3868 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09553 vdd 6984 3875 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09552 3873 3875 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09551 vdd 4093 3874 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09550 985 2122 890 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09549 890 2124 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09548 vdd 2125 890 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09547 980 985 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09546 889 981 985 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09545 890 982 889 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09544 5786 5787 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09543 vdd 5893 5786 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09542 5784 5786 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09541 4711 5341 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09540 vdd 5992 4711 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09539 5753 4711 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09538 541 2411 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09537 vdd 2615 541 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09536 1033 541 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09535 1617 1779 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09534 1988 4087 1617 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09533 vdd 1991 1988 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09532 4102 4188 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09531 4100 4189 4183 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09530 vdd 6187 4100 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09529 4186 4189 4102 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09528 4101 4190 4186 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09527 vdd 4184 4101 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09526 4184 4186 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09525 4183 4190 4184 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09524 vdd 4183 6187 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09523 6187 4183 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09522 vdd 5054 4190 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09521 4189 4190 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09520 vdd 4191 4188 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09519 vdd 6921 5771 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09518 5771 6691 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09517 5770 6440 5771 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09516 5769 5999 5770 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09515 5771 6000 5769 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09514 826 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09513 2142 1190 826 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09512 vdd 825 2142 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09511 2373 4051 2374 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09510 2374 2799 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09509 vdd 2790 2373 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09508 2371 2373 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09507 6352 6740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09506 4163 4918 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09505 4024 3796 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09504 2894 3460 3660 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09503 3067 3263 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09502 vdd 3067 2894 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09501 1273 3051 1381 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09500 1274 1380 1273 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09499 vdd 1749 1274 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09498 2448 2572 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09497 2446 2573 2567 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09496 vdd 3802 2446 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09495 2570 2573 2448 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09494 2447 2574 2570 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09493 vdd 2568 2447 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09492 2568 2570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09491 2567 2574 2568 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09490 vdd 2567 3802 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09489 3802 2567 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09488 vdd 3259 2574 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09487 2573 2574 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09486 vdd 2792 2572 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09485 3241 4083 3242 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09484 3240 3637 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09483 vdd 3240 3241 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09482 781 2747 782 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09481 782 1904 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09480 vdd 3217 782 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09479 779 781 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09478 780 4176 781 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09477 782 1322 780 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09476 3637 4265 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09475 vdd 5773 3637 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09474 6811 6820 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09473 4836 5026 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09472 6835 6850 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09471 6112 5524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09470 6695 6694 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09469 6935 6934 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09468 3989 5054 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09467 vdd 3989 3987 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09466 3988 3986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09465 vdd 3988 3983 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09464 3983 3987 3985 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09463 3985 3989 3984 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09462 3980 3979 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09461 vdd 3981 3979 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09460 3979 3981 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09459 3984 3982 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09458 3982 3985 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09457 vdd 6976 3982 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09456 3981 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09455 3981 3987 3980 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09454 3982 3989 3981 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09453 4122 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09452 4401 6877 4122 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09451 vdd 4914 4401 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09450 6583 6877 6584 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09449 6584 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09448 vdd 6905 6583 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09447 6586 6583 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09446 5954 5329 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09445 vdd 5552 5954 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09444 5551 6238 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09443 vdd 6440 5551 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09442 1706 2544 1265 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09441 1265 2142 1706 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09440 vdd 1356 1265 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09439 4733 4491 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09438 vdd 5773 4733 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09437 4224 3604 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09436 5409 5993 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09435 5531 5967 5409 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09434 vdd 5964 5531 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09433 1181 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09432 1679 1190 1181 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09431 vdd 1182 1679 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09430 3670 4880 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09429 3736 4881 3670 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09428 vdd 3969 3736 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09427 4832 5372 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09426 vdd 5157 4831 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09425 vdd 5893 4833 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09424 4965 5893 4832 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09423 4831 4833 4965 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09422 5164 4965 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09421 3265 5262 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09420 vdd 3263 3264 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09419 vdd 5893 3267 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09418 3266 5893 3265 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09417 3264 3267 3266 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09416 3262 3266 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09415 4536 5243 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09414 vdd 4748 4535 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09413 vdd 5893 4538 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09412 4537 5893 4536 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09411 4535 4538 4537 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09410 4751 4537 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09409 4117 4308 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09408 vdd 4524 4116 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09407 vdd 5893 4309 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09406 4307 5893 4117 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09405 4116 4309 4307 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09404 4531 4307 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09403 6601 6434 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09402 vdd 6919 6601 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09401 1514 3586 1515 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09400 1515 2755 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09399 vdd 2111 1514 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09398 1513 1514 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09397 vdd 1188 893 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09396 891 3408 982 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09395 892 2770 891 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09394 893 1189 892 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09393 4622 4744 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09392 vdd 4745 4622 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09391 vdd 1641 1630 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09390 1882 1893 1595 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09389 1595 1641 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09388 1595 1630 1882 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09387 vdd 1628 1595 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09386 1628 1893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09385 2855 6727 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09384 vdd 2852 2854 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09383 vdd 5893 2856 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09382 2853 5893 2855 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09381 2854 2856 2853 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09380 2851 2853 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09379 3308 6265 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09378 vdd 3460 3307 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09377 vdd 5893 3464 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09376 3462 5893 3308 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09375 3307 3464 3462 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09374 3459 3462 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09373 4115 5902 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09372 vdd 4299 4114 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09371 vdd 5893 4304 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09370 4302 5893 4115 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09369 4114 4304 4302 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09368 4300 4302 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09367 1372 690 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09366 vdd 857 1372 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09365 4069 4273 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09364 vdd 4068 4069 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09363 4503 4069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09362 3821 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09361 vdd 6440 3821 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09360 3625 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09359 vdd 6440 3625 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09358 6024 5762 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09357 vdd 6748 6024 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09356 4521 4512 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09355 vdd 6690 4521 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09354 4971 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09353 5017 6877 4971 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09352 vdd 5524 5017 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09351 1664 2325 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09350 vdd 3178 1664 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09349 1662 1664 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09348 vdd 5773 4141 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09347 4141 4491 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09346 4505 5992 4141 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09345 4140 4726 4505 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09344 4141 4265 4140 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09343 5406 5805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09342 5746 5756 5406 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09341 vdd 6905 5746 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09340 vdd 3967 3719 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09339 3719 3715 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09338 vdd 4838 3719 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09337 3714 3719 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09336 vdd 4181 3730 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09335 3730 3728 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09334 vdd 4399 3730 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09333 3727 3730 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09332 vdd 5440 5439 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09331 5439 5436 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09330 vdd 5442 5439 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09329 5680 5439 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09328 vdd 6839 6623 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09327 6623 6820 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09326 vdd 6850 6623 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09325 6622 6623 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09324 887 918 979 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09323 888 919 887 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09322 vdd 2537 888 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09321 1534 979 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09320 1787 4299 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09319 vdd 5363 1787 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09318 2407 1787 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09317 1676 2347 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09316 1676 3593 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09315 vdd 1688 1676 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09314 vdd 1679 1676 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09313 3667 6190 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09312 3725 6191 3667 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09311 vdd 3969 3725 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09310 vdd 5068 4693 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09309 4693 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09308 4693 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09307 vdd 5372 4693 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09306 4895 4693 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09305 298 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09304 953 305 298 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09303 299 312 953 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09302 vdd 302 299 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09301 2753 2752 2754 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09300 2751 2749 2753 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09299 vdd 2750 2751 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09298 6173 2754 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09297 2791 2799 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09296 3738 4051 2791 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09295 vdd 2790 3738 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09294 4936 5112 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09293 5326 5113 4936 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09292 vdd 4935 5326 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09291 5719 6877 5720 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09290 5720 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09289 vdd 6591 5719 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09288 5952 5719 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09287 1271 1565 1735 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09286 1368 1367 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09285 vdd 1368 1271 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09284 5803 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09283 vdd 5803 5802 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09282 5801 5800 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09281 vdd 5801 5798 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09280 5798 5802 5797 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09279 5797 5803 5799 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09278 5795 6682 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09277 vdd 5794 6682 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09276 6682 5794 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09275 5799 5796 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09274 5796 5797 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09273 vdd 6976 5796 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09272 5794 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09271 5794 5802 5795 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09270 5796 5803 5794 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09269 vdd 4491 3638 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09268 3638 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09267 vdd 4275 3638 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09266 4083 3638 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09265 1264 1346 1347 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09264 1263 2778 1264 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09263 1262 2766 1263 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09262 vdd 1345 1262 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09261 2553 1347 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09260 vdd 216 91 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09259 212 787 24 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09258 24 216 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09257 24 91 212 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09256 vdd 92 24 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09255 92 787 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09254 1579 5359 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09253 1579 2412 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09252 vdd 2406 1579 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09251 1964 3259 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09250 vdd 1964 1963 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09249 1962 1959 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09248 vdd 1962 1961 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09247 1961 1963 1960 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09246 1960 1964 1958 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09245 1955 4241 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09244 vdd 1956 4241 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09243 4241 1956 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09242 1958 1957 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09241 1957 1960 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09240 vdd 6976 1957 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09239 1956 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09238 1956 1963 1955 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09237 1957 1964 1956 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09236 3185 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09235 vdd 4205 3185 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09234 3187 3185 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09233 3062 3836 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09232 3062 2407 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09231 vdd 2406 3062 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09230 4523 3060 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09229 4523 3062 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09228 vdd 4509 4523 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09227 1192 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09226 1933 1190 1192 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09225 vdd 1191 1933 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09224 6415 6675 6287 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09223 6287 6637 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09222 vdd 6413 6415 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09221 6414 6415 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09220 6138 6140 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09219 6134 6141 6133 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09218 vdd 6165 6134 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09217 6137 6141 6138 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09216 6136 6142 6137 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09215 vdd 6135 6136 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09214 6135 6137 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09213 6133 6142 6135 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09212 vdd 6133 6165 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09211 6165 6133 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09210 vdd 6832 6142 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09209 6141 6142 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09208 vdd 6139 6140 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09207 vdd 1652 471 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09206 470 1508 469 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09205 469 1652 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09204 469 471 470 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09203 vdd 468 469 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09202 468 1508 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09201 499 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09200 641 987 499 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09199 vdd 504 641 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09198 4422 4423 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09197 4417 4424 4418 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09196 vdd 5268 4417 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09195 4421 4424 4422 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09194 4420 4425 4421 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09193 vdd 4419 4420 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09192 4419 4421 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09191 4418 4425 4419 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09190 vdd 4418 5268 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09189 5268 4418 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09188 vdd 5054 4425 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09187 4424 4425 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09186 vdd 4589 4423 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09185 15 123 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09184 13 50 121 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09183 vdd 525 13 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09182 48 50 15 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09181 14 124 48 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09180 vdd 47 14 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09179 47 48 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09178 121 124 47 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09177 vdd 121 525 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09176 525 121 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09175 vdd 3259 124 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09174 50 124 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09173 vdd 255 123 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09172 vdd 4094 2030 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09171 2030 4524 2170 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09170 vdd 6165 5731 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09169 5731 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09168 5731 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09167 vdd 6440 5731 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09166 5730 5731 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09165 vdd 6522 5970 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09164 5970 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09163 5970 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09162 vdd 6440 5970 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09161 5971 5970 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09160 5408 5525 5523 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09159 5407 5983 5408 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09158 vdd 5521 5407 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09157 4468 4708 5880 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09156 4467 4466 4468 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09155 vdd 6224 4467 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09154 vdd 2194 852 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09153 852 857 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09152 852 1953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09151 vdd 3836 852 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09150 1029 852 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09149 vdd 1218 1013 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09148 1013 1732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09147 1013 4239 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09146 vdd 4748 1013 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09145 1169 1013 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09144 3583 5054 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09143 vdd 3583 3582 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09142 3581 3758 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09141 vdd 3581 3580 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09140 3580 3582 3579 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09139 3579 3583 3577 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09138 3575 3759 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09137 vdd 3576 3759 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09136 3759 3576 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09135 3577 3578 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09134 3578 3579 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09133 vdd 6976 3578 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09132 3576 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09131 3576 3582 3575 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09130 3578 3583 3576 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09129 3 96 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09128 1 30 95 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09127 vdd 633 1 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09126 29 30 3 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09125 2 99 29 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09124 vdd 27 2 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09123 27 29 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09122 95 99 27 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09121 vdd 95 633 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09120 633 95 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09119 vdd 3160 99 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09118 30 99 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09117 vdd 222 96 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09116 4416 4673 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09115 4587 4671 4416 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09114 vdd 5927 4587 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09113 6124 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09112 6123 6877 6124 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09111 vdd 6807 6123 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09110 vdd 6876 6110 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09109 6110 6877 6213 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09108 6421 6213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09107 vdd 5748 2828 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09106 2828 3049 2829 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09105 2827 2829 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09104 204 320 205 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09103 205 319 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09102 vdd 328 204 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09101 310 204 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09100 4569 5753 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09099 4927 5767 4569 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09098 vdd 5670 4927 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09097 264 3229 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09096 vdd 4501 264 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09095 1601 3391 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09094 1647 2326 1601 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09093 vdd 2111 1647 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09092 4954 5144 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09091 4954 5570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09090 vdd 5788 4954 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09089 5569 5575 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09088 5569 5570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09087 vdd 5788 5569 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09086 5556 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09085 5556 5570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09084 vdd 5788 5556 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09083 vdd 2050 2022 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09082 2023 2146 2139 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09081 2024 2052 2023 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09080 2022 2051 2024 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09079 4563 4699 4608 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09078 4562 4921 4563 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09077 vdd 4916 4562 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09076 2747 5959 2748 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09075 2748 3186 2747 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09074 vdd 3191 2748 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09073 528 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09072 2165 987 528 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09071 vdd 527 2165 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09070 vdd 6622 6620 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09069 6619 6740 6621 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09068 6621 6622 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09067 6621 6620 6619 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09066 vdd 6618 6621 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09065 6618 6740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09064 6662 6889 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09063 6660 6661 6662 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09062 vdd 6867 6660 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09061 6627 6820 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09060 6627 6631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09059 vdd 6806 6627 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09058 2598 3259 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09057 vdd 2598 2599 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09056 2597 2601 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09055 vdd 2597 2453 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09054 2453 2599 2594 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09053 2594 2598 2452 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09052 2451 4235 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09051 vdd 2591 4235 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09050 4235 2591 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09049 2452 2593 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09048 2593 2594 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09047 vdd 6976 2593 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09046 2591 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09045 2591 2599 2451 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09044 2593 2598 2591 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09043 5564 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09042 5564 5570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09041 vdd 5788 5564 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09040 5348 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09039 5348 5141 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09038 vdd 5140 5348 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09037 3234 5359 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09036 3234 2412 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09035 vdd 2406 3234 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09034 vdd 4748 3234 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09033 2479 2487 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09032 vdd 2734 2479 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09031 2485 2487 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09030 vdd 2730 2485 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09029 4402 4401 4403 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09028 4403 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09027 vdd 6678 4403 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09026 4399 4402 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09025 4400 6637 4402 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09024 4403 4653 4400 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09023 6842 6850 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09022 6842 6631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09021 vdd 6806 6842 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09020 596 1652 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09019 vdd 1505 596 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09018 4212 4253 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09017 4212 3629 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09016 vdd 3831 4212 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09015 vdd 3827 4212 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09014 5787 6963 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09013 5787 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09012 vdd 6952 5787 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09011 2196 1990 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09010 2196 1988 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09009 vdd 1989 2196 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09008 vdd 6170 6171 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09007 6171 6636 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09006 vdd 6372 6171 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09005 6169 6171 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09004 5973 6375 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09003 5973 6374 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09002 vdd 6423 5973 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09001 vdd 6571 5973 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09000 5790 5907 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08999 vdd 6440 5790 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08998 5789 5790 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08997 297 461 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_08996 579 301 297 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_08995 296 1169 579 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_08994 vdd 581 296 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_08993 1173 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08992 5947 1649 1173 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08991 vdd 1172 5947 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08990 501 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08989 624 987 501 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08988 vdd 500 624 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08987 3049 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08986 3049 4942 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08985 vdd 4941 3049 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08984 vdd 5157 2632 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08983 vdd 4299 2634 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08982 2632 2634 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08981 6351 6348 6278 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08980 6278 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08979 vdd 6678 6278 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08978 6347 6351 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08977 6277 6637 6351 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08976 6278 6613 6277 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08975 4207 5300 4109 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08974 4109 6220 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08973 vdd 4205 4207 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08972 4892 4207 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08971 4944 5116 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08970 5336 5125 4944 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08969 vdd 4945 5336 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08968 vdd 2396 2397 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08967 2397 2827 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08966 2397 2607 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08965 vdd 2506 2397 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08964 4946 2397 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08963 1939 2050 1940 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08962 1938 2146 1939 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08961 1937 2052 1938 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08960 vdd 2051 1937 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08959 4671 1940 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08958 1935 2356 1936 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08957 1936 2553 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08956 vdd 2514 1935 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08955 2051 1935 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08954 1134 1188 1187 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08953 1133 1189 1134 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08952 vdd 2770 1133 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08951 1340 1187 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08950 vdd 3263 867 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08949 867 3460 866 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08948 1234 866 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08947 2893 3263 4286 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08946 3064 5363 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08945 vdd 3064 2893 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08944 2436 2535 2536 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08943 2533 2534 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08942 vdd 2533 2436 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08941 4848 4847 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08940 4849 4850 4848 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08939 vdd 6867 4849 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08938 vdd 5773 4500 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08937 4500 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08936 4500 4748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08935 vdd 6440 4500 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08934 4499 4500 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08933 3194 3202 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08932 vdd 3197 3194 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08931 3193 3194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08930 1487 2304 1486 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08929 1486 1888 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08928 vdd 1884 1487 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08927 1485 1487 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08926 vdd 5014 4834 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08925 4847 4836 4837 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08924 4837 5014 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08923 4837 4834 4847 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08922 vdd 4835 4837 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08921 4835 4836 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08920 3627 3639 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_08919 5502 3821 3627 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_08918 3626 3624 5502 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_08917 vdd 3625 3626 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_08916 4092 5157 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08915 vdd 4299 4092 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08914 4091 4092 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08913 1734 1732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08912 vdd 1760 1734 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08911 2155 1734 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08910 136 138 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08909 vdd 2387 136 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08908 1190 136 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08907 5391 5584 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08906 5389 5583 5577 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08905 vdd 5575 5389 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08904 5581 5583 5391 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08903 5390 5586 5581 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08902 vdd 5578 5390 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08901 5578 5581 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08900 5577 5586 5578 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08899 vdd 5577 5575 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08898 5575 5577 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08897 vdd 6984 5586 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08896 5583 5586 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08895 vdd 5580 5584 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08894 4529 4532 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08893 4526 4534 4525 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08892 vdd 4524 4526 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08891 4530 4534 4529 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08890 4528 4533 4530 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08889 vdd 4527 4528 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08888 4527 4530 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08887 4525 4533 4527 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08886 vdd 4525 4524 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08885 4524 4525 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08884 vdd 6984 4533 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08883 4534 4533 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08882 vdd 4531 4532 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08881 6249 6247 6250 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08880 6248 6475 6249 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08879 vdd 6245 6248 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08878 vdd 1304 1166 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08877 1694 1165 1168 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08876 1168 1304 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08875 1168 1166 1694 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08874 vdd 1167 1168 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08873 1167 1165 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08872 496 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08871 629 1190 496 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08870 vdd 636 629 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08869 vdd 86 73 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08868 73 772 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08867 vdd 1151 73 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08866 320 73 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08865 vdd 4927 4930 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08864 4930 4929 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08863 4930 5518 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08862 vdd 4928 4930 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08861 5106 4930 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08860 3207 3414 3206 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08859 3206 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08858 vdd 5262 3207 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08857 3212 3207 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08856 vdd 5877 4037 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08855 4037 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08854 vdd 6440 4037 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08853 4038 4037 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08852 vdd 5749 4923 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08851 4923 5748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08850 4923 6591 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08849 vdd 6440 4923 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08848 4921 4923 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08847 vdd 2194 1207 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08846 1207 1953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08845 vdd 3836 1207 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08844 2124 1207 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08843 vdd 5759 3433 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08842 3433 3430 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08841 vdd 3789 3433 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08840 3429 3433 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08839 vdd 2320 2317 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08838 2499 2319 2321 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08837 2321 2320 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08836 2321 2317 2499 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08835 vdd 2318 2321 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08834 2318 2319 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08833 vdd 2356 2029 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08832 2029 2155 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08831 2600 2156 2029 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08830 2028 4673 2600 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08829 2029 4671 2028 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08828 2992 3414 2873 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08827 2873 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08826 vdd 5272 2992 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08825 2990 2992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08824 5520 6214 5387 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08823 5387 5986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08822 vdd 6850 5520 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08821 5521 5520 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08820 5910 6665 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08819 6886 6885 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08818 4028 3421 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08817 3641 4239 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08816 5244 5670 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08815 6861 6874 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08814 vdd 5069 2166 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08813 2166 2807 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08812 2166 2583 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08811 vdd 5992 2166 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08810 2381 2166 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08809 vdd 3866 1397 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08808 1397 2125 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08807 1397 3849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08806 vdd 3664 1397 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08805 1975 1397 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08804 vdd 6186 6189 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08803 6189 6431 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08802 6184 6187 6189 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08801 6185 6182 6184 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08800 6189 6183 6185 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08799 533 535 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08798 529 536 530 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08797 vdd 3434 529 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08796 534 536 533 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08795 532 537 534 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08794 vdd 531 532 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08793 531 534 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08792 530 537 531 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08791 vdd 530 3434 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08790 3434 530 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08789 vdd 3259 537 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08788 536 537 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08787 vdd 677 535 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08786 5837 6420 6637 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08785 5836 6222 5837 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08784 vdd 6422 5836 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08783 5412 5789 5549 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08782 5411 5548 5412 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08781 vdd 6004 5411 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08780 637 1190 544 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08779 544 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08778 vdd 636 637 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08777 1188 637 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08776 4137 5112 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08775 4928 5113 4137 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08774 vdd 4239 4928 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08773 vdd 3866 1774 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08772 1774 1778 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08771 1774 3849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08770 vdd 3664 1774 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08769 3229 1774 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08768 6903 6906 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08767 4059 3434 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08766 6310 6905 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08765 4043 3802 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08764 3653 3451 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08763 vdd 5992 3653 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08762 3863 4091 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08761 vdd 4286 3863 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08760 4555 4692 4883 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08759 4686 4685 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08758 vdd 4686 4555 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08757 5468 5270 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08756 vdd 5474 5468 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08755 6015 5907 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08754 vdd 6025 6015 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08753 3247 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08752 3246 4273 3247 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08751 vdd 4937 3246 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08750 6879 6877 6741 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08749 6741 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08748 vdd 6874 6879 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08747 6875 6879 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08746 6191 3184 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08745 vdd 3183 6191 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08744 2793 3182 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08743 vdd 3174 2793 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08742 6412 6414 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08741 vdd 6410 6412 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08740 6418 6412 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08739 5830 5967 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08738 5969 5993 5830 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08737 vdd 5965 5969 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08736 5330 5331 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08735 vdd 6690 5330 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08734 5329 5330 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08733 4489 3658 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08732 4489 4062 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08731 vdd 5069 4489 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08730 vdd 5363 4489 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08729 975 641 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08728 975 981 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08727 vdd 3195 975 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08726 vdd 629 975 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08725 495 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08724 625 1190 495 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08723 vdd 633 625 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08722 vdd 2913 2473 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08721 2507 2712 2422 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08720 2422 2913 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08719 2422 2473 2507 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08718 vdd 2470 2422 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08717 2470 2712 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08716 2315 2520 2316 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08715 2316 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08714 vdd 2314 2315 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08713 2487 2315 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08712 4885 5954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08711 4886 5502 4885 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08710 vdd 5959 4886 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08709 vdd 3856 3249 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08708 3249 3853 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08707 vdd 4275 3249 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08706 3248 3249 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08705 vdd 4953 4951 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08704 4951 4952 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08703 vdd 5154 4951 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08702 5140 4951 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08701 vdd 2779 2745 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08700 2745 3182 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08699 vdd 3174 2745 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08698 2744 2745 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08697 1618 3460 1991 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08696 1789 2852 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08695 vdd 1789 1618 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08694 1574 1745 1573 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08693 1573 1989 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08692 vdd 1572 1574 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08691 2396 1574 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08690 1718 2350 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08689 vdd 2534 1718 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08688 1716 1718 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08687 2947 5953 2864 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08686 vdd 2952 2864 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08685 2864 3186 2947 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08684 2946 2947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08683 1503 2326 1504 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08682 1504 3391 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08681 vdd 2111 1503 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08680 1501 1503 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08679 3295 3607 4466 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08678 3422 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08677 vdd 3422 3295 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08676 vdd 216 84 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08675 86 615 23 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08674 23 216 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08673 23 84 86 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08672 vdd 85 23 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08671 85 615 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08670 vdd 3866 1751 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08669 1751 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08668 1751 2406 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08667 vdd 3836 1751 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08666 1749 1751 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08665 1556 1968 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08664 vdd 1559 1556 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08663 1703 1556 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08662 2524 2521 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08661 vdd 2520 2524 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08660 2522 2524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08659 6270 6328 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08658 6268 6330 6322 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08657 vdd 6522 6268 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08656 6327 6330 6270 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08655 6269 6331 6327 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08654 vdd 6324 6269 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08653 6324 6327 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08652 6322 6331 6324 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08651 vdd 6322 6522 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08650 6522 6322 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08649 vdd 6832 6331 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08648 6330 6331 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08647 vdd 6326 6328 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08646 3056 3263 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08645 vdd 5363 3056 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08644 4942 3056 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08643 vdd 1478 1240 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08642 1240 1480 1280 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08641 4474 5125 4473 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08640 4473 4472 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08639 vdd 4471 4474 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08638 4952 4474 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08637 2540 5958 2438 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08636 2438 2773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08635 vdd 4205 2438 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08634 2537 2540 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08633 2437 3199 2540 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08632 2438 3618 2437 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08631 2715 2716 2714 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08630 2714 2915 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08629 vdd 2717 2715 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08628 2712 2715 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08627 vdd 3231 3228 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08626 3228 4258 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08625 vdd 3438 3228 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08624 3227 3228 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08623 3656 3866 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08622 vdd 3664 3656 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08621 3853 3656 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08620 vdd 1732 1219 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08619 1219 1218 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08618 vdd 4748 1219 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08617 1564 1219 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08616 1709 2349 1592 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08615 vdd 1716 1592 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08614 1592 2553 1709 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08613 1708 1709 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08612 278 347 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08611 276 348 342 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08610 vdd 1182 276 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08609 345 348 278 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08608 277 349 345 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08607 vdd 343 277 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08606 343 345 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08605 342 349 343 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08604 vdd 342 1182 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08603 1182 342 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08602 vdd 3160 349 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08601 348 349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08600 vdd 350 347 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08599 6326 6175 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08598 vdd 6143 6326 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08597 vdd 4492 4494 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08596 4495 4497 4496 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08595 4493 4499 4495 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08594 4494 4725 4493 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08593 5325 5523 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08592 vdd 5324 5325 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08591 vdd 5144 2036 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08590 2036 5359 2192 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08589 2193 2192 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08588 133 405 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08587 vdd 4299 133 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08586 5453 5701 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08585 vdd 5265 5453 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08584 vdd 6622 6356 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08583 6359 6352 6279 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08582 6279 6622 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08581 6279 6356 6359 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08580 vdd 6354 6279 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08579 6354 6352 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08578 6666 6668 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08577 6667 6676 6666 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08576 vdd 6867 6667 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08575 5030 6600 4975 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08574 4975 6447 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08573 vdd 6601 5030 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08572 5029 5030 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08571 5839 6422 5981 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08570 5838 6420 5839 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08569 vdd 6222 5838 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08568 6867 5981 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08567 5132 6447 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08566 5132 5125 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08565 vdd 5133 5132 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08564 573 1876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08563 573 579 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08562 vdd 2727 573 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08561 6390 6874 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08560 6390 6631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08559 vdd 6806 6390 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08558 5842 6906 5982 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08557 5841 6420 5842 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08556 5840 6222 5841 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08555 vdd 6422 5840 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08554 6208 5982 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08553 vdd 4397 4398 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08552 4398 4849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08551 vdd 5025 4398 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08550 4396 4398 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08549 4609 6951 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08548 4609 4469 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08547 vdd 4470 4609 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08546 2993 4608 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08545 vdd 2996 2993 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08544 4915 5756 4917 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08543 4917 5805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08542 vdd 4914 4915 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08541 4916 4915 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08540 267 1583 266 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08539 266 3460 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08538 vdd 264 267 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08537 265 267 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08536 2773 2578 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08535 vdd 3438 2773 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08534 vdd 3734 3723 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08533 3723 3720 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08532 vdd 4843 3723 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08531 3717 3723 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08530 6405 6885 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08529 6405 6631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08528 vdd 6806 6405 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08527 6663 6877 6664 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08526 6664 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08525 vdd 6885 6663 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08524 6661 6663 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08523 vdd 5329 4926 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08522 4926 5552 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08521 vdd 5116 4926 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08520 6600 4926 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08519 484 489 485 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08518 485 2506 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08517 vdd 1737 485 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08516 482 484 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08515 483 491 484 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08514 485 486 483 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08513 vdd 3592 3287 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08512 3287 3404 3407 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08511 3408 3407 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08510 vdd 5068 5070 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08509 5070 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08508 5070 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08507 vdd 6265 5070 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08506 5496 5070 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08505 4025 4275 4026 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08504 4023 4024 4025 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08503 4022 4708 4023 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08502 vdd 6224 4022 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08501 4469 4026 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08500 1978 2406 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08499 vdd 3836 1978 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08498 2182 1978 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08497 6345 6609 6275 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08496 6275 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08495 vdd 6678 6275 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08494 6342 6345 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08493 6274 6637 6345 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08492 6275 6607 6274 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08491 4119 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08490 4157 6877 4119 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08489 vdd 5026 4157 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08488 6264 6263 6466 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08487 6262 6261 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08486 vdd 6262 6264 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08485 vdd 6959 6954 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08484 6954 6957 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08483 vdd 6952 6954 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08482 6968 6954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08481 vdd 4896 4894 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08480 4894 4895 5277 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08479 vdd 1737 1721 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08478 1721 1904 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08477 vdd 2375 1721 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08476 1722 1721 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08475 vdd 3217 785 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08474 785 1904 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08473 784 2747 785 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08472 783 4176 784 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08471 785 1322 783 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08470 3700 4250 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08469 3827 4491 3700 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08468 vdd 5349 3827 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08467 3209 4014 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08466 vdd 3416 3209 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08465 3208 3209 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08464 5808 5996 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08463 5806 5885 5991 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08462 vdd 5992 5806 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08461 5884 5885 5808 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08460 5807 5886 5884 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08459 vdd 5882 5807 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08458 5882 5884 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08457 5991 5886 5882 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08456 vdd 5991 5992 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08455 5992 5991 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08454 vdd 6984 5886 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08453 5885 5886 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08452 vdd 5994 5996 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08451 vdd 1304 1305 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08450 4880 1300 1247 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08449 1247 1304 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08448 1247 1305 4880 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08447 vdd 1302 1247 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08446 1302 1300 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08445 vdd 611 326 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08444 326 323 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08443 vdd 332 326 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08442 322 326 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08441 4063 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08440 vdd 6440 4063 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08439 4062 4063 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08438 2631 2632 2460 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08437 2460 2629 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08436 vdd 4280 2631 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08435 2628 2631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08434 6280 6359 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08433 6360 6624 6280 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08432 vdd 6867 6360 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08431 4546 4752 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08430 4544 4639 4749 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08429 vdd 4748 4544 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08428 4638 4639 4546 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08427 4545 4640 4638 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08426 vdd 4636 4545 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08425 4636 4638 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08424 4749 4640 4636 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08423 vdd 4749 4748 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08422 4748 4749 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08421 vdd 6984 4640 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08420 4639 4640 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08419 vdd 4751 4752 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08418 vdd 2352 1056 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08417 1056 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08416 vdd 3664 1056 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08415 2615 1056 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08414 vdd 2506 1713 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08413 1713 2371 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08412 vdd 2782 1713 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08411 1904 1713 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08410 vdd 4942 4931 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08409 4931 4941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08408 vdd 5992 4931 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08407 5805 4931 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08406 5396 5954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08405 5483 5502 5396 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08404 vdd 5958 5483 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08403 vdd 6919 5256 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08402 5256 6434 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08401 5259 6867 5256 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08400 5255 6115 5259 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08399 5256 5254 5255 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08398 6950 6963 6755 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08397 vdd 6948 6755 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08396 6755 6959 6950 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08395 6946 6950 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08394 5516 5756 5386 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08393 5386 5805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08392 vdd 5524 5516 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08391 5733 5516 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08390 2377 4051 2378 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08389 2378 2799 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08388 vdd 2384 2377 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08387 2501 2377 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08386 6224 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08385 4282 5575 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08384 6581 6807 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08383 vdd 2487 2486 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08382 2483 2734 2423 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08381 2423 2487 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08380 2423 2486 2483 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08379 vdd 2482 2423 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08378 2482 2734 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08377 vdd 5749 5511 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08376 5511 5748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08375 5511 6874 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08374 vdd 6440 5511 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08373 5510 5511 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08372 5385 5472 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08371 5383 5471 5465 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08370 vdd 6591 5383 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08369 5469 5471 5385 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08368 5384 5473 5469 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08367 vdd 5466 5384 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08366 5466 5469 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08365 5465 5473 5466 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08364 vdd 5465 6591 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08363 6591 5465 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08362 vdd 6832 5473 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08361 5471 5473 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08360 vdd 5468 5472 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08359 6473 6243 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08358 vdd 6242 6473 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08357 2357 2553 2361 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08356 2358 2356 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08355 vdd 2358 2357 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08354 393 987 294 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08353 294 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08352 vdd 392 393 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08351 1345 393 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08350 1526 1919 1525 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08349 1525 1918 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08348 vdd 2521 1526 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08347 1524 1526 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08346 vdd 4088 3859 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08345 3859 4091 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08344 3859 4089 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08343 vdd 4087 3859 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08342 5877 3859 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08341 5567 6682 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08340 3634 5359 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08339 4280 5144 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08338 3037 4235 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08337 1576 4937 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08336 3040 4935 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08335 5303 5315 5305 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08334 5304 5971 5303 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08333 vdd 5312 5304 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08332 vdd 6616 5697 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08331 5695 6591 5696 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08330 5696 6616 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08329 5696 5697 5695 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08328 vdd 5694 5696 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08327 5694 6591 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08326 6160 5708 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08325 vdd 6166 6160 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08324 6672 6893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08323 vdd 6893 6670 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08322 6669 6906 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08321 vdd 6669 6672 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08320 6672 6670 6671 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08319 6671 6906 6672 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08318 6668 6671 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08317 vdd 6671 6668 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08316 4668 4918 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08315 4668 6910 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08314 vdd 6806 4668 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08313 4961 5361 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08312 vdd 4953 4961 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08311 vdd 918 800 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08310 798 3210 801 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08309 799 2537 798 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08308 800 919 799 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08307 3369 4942 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08306 vdd 3658 3369 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08305 4261 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08304 539 2195 540 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08303 540 2194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08302 vdd 6440 539 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08301 1732 539 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08300 6150 6628 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08299 vdd 5864 6150 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08298 3624 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08297 vdd 3818 3624 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08296 4019 4213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08295 4018 4212 4019 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08294 vdd 5299 4018 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08293 1482 1641 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08292 vdd 1893 1482 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08291 2127 2122 2021 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08290 2021 2124 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08289 vdd 2125 2021 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08288 2526 2127 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08287 2020 2535 2127 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08286 2021 2737 2020 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08285 6761 6792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08284 6802 6794 6761 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08283 vdd 6867 6802 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08282 vdd 1330 1252 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08281 1252 1328 1325 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08280 5045 1325 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08279 vdd 6714 6711 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08278 vdd 6952 6712 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08277 6711 6712 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08276 2309 2320 2310 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08275 2310 2319 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08274 vdd 2485 2309 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08273 2308 2309 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08272 6765 6847 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08271 6849 6851 6765 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08270 vdd 6867 6849 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08269 5906 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08268 vdd 5906 5905 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08267 5904 5903 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08266 vdd 5904 5810 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08265 5810 5905 5900 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08264 5900 5906 5809 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08263 5852 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08262 vdd 6019 6714 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08261 6714 6019 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08260 5809 5897 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08259 5897 5900 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08258 vdd 6976 5897 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08257 6019 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08256 6019 5905 5852 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08255 5897 5906 6019 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08254 vdd 5914 5247 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08253 5247 5670 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08252 vdd 6665 5247 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08251 6116 5247 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08250 4554 5045 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08249 5088 5044 4554 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08248 vdd 5964 5088 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08247 190 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08246 189 191 190 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08245 188 200 189 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08244 vdd 322 188 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08243 571 189 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08242 vdd 2913 2914 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08241 5723 2909 2881 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08240 2881 2913 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08239 2881 2914 5723 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08238 vdd 2910 2881 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08237 2910 2909 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08236 1877 936 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08235 vdd 1479 1877 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08234 4982 5958 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08233 vdd 5262 4981 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08232 vdd 5309 5061 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08231 5059 5309 4982 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08230 4981 5061 5059 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08229 5057 5059 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08228 4106 5959 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08227 vdd 5243 4105 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08226 vdd 5309 4199 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08225 4198 5309 4106 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08224 4105 4199 4198 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08223 4434 4198 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08222 4006 5725 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08221 vdd 4308 4003 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08220 vdd 5309 4005 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08219 4004 5309 4006 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08218 4003 4005 4004 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08217 4002 4004 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08216 5274 5953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08215 vdd 5272 5275 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08214 vdd 5309 5276 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08213 5273 5309 5274 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08212 5275 5276 5273 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08211 5715 5273 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08210 vdd 6667 6206 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08209 6206 6205 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08208 vdd 6207 6206 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08207 6204 6206 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08206 2816 3259 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08205 vdd 2816 2815 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08204 2813 2826 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08203 vdd 2813 2814 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08202 2814 2815 2812 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08201 2812 2816 2811 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08200 2808 4935 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08199 vdd 2809 4935 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08198 4935 2809 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08197 2811 2810 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08196 2810 2812 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08195 vdd 6976 2810 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08194 2809 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08193 2809 2815 2808 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08192 2810 2816 2809 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08191 vdd 5549 4940 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08190 4940 4946 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08189 vdd 4947 4940 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08188 4939 4940 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08187 5848 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08186 6011 6469 5848 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08185 vdd 6442 6011 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08184 4708 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08183 4708 4287 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08182 vdd 4089 4708 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08181 vdd 3866 4708 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08180 2003 2298 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08179 2292 2301 2003 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08178 vdd 2086 2292 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08177 463 571 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08176 vdd 766 463 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08175 461 463 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08174 6710 6715 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08173 6708 6962 6710 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08172 6709 6711 6708 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08171 vdd 6956 6709 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08170 6707 6708 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08169 vdd 1212 1213 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08168 1213 3217 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08167 vdd 1985 1213 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08166 1558 1213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08165 vdd 1975 1050 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08164 1050 1234 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08163 vdd 1233 1050 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08162 1380 1050 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08161 620 640 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08160 vdd 2314 620 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08159 619 620 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08158 1239 5363 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08157 1239 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08156 vdd 4524 1239 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08155 6738 6831 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08154 6736 6833 6825 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08153 vdd 6850 6736 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08152 6827 6833 6738 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08151 6737 6834 6827 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08150 vdd 6826 6737 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08149 6826 6827 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08148 6825 6834 6826 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08147 vdd 6825 6850 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08146 6850 6825 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08145 vdd 6832 6834 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08144 6833 6834 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08143 vdd 6830 6831 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08142 4856 4855 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08141 4865 4854 4856 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08140 vdd 6867 4865 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08139 vdd 5245 4149 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08138 5004 5670 4118 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08137 4118 5245 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08136 4118 4149 5004 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08135 vdd 4146 4118 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08134 4146 5670 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08133 vdd 6480 6296 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08132 6296 6682 6692 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08131 vdd 946 560 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08130 560 586 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08129 581 2086 560 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08128 559 588 581 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08127 560 774 559 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08126 vdd 619 608 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08125 607 1317 565 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08124 565 619 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08123 565 608 607 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08122 vdd 605 565 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08121 605 1317 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08120 vdd 212 213 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08119 213 772 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08118 vdd 1151 213 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08117 486 213 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08116 2328 3186 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08115 vdd 6187 2328 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08114 2326 2328 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08113 3594 4008 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08112 vdd 3595 3594 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08111 3593 3594 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08110 6273 6337 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08109 6271 6340 6332 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08108 vdd 6376 6271 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08107 6338 6340 6273 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08106 6272 6341 6338 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08105 vdd 6334 6272 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08104 6334 6338 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08103 6332 6341 6334 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08102 vdd 6332 6376 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08101 6376 6332 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08100 vdd 6832 6341 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08099 6340 6341 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08098 vdd 6336 6337 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08097 5124 5125 4992 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08096 4992 6447 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08095 vdd 5544 5124 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08094 5338 5124 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08093 2435 3586 2532 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08092 2531 2530 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08091 vdd 2531 2435 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08090 1523 1919 1522 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08089 1522 1918 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08088 vdd 2349 1523 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08087 1521 1523 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08086 vdd 5320 5323 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08085 5323 5321 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08084 5323 5322 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08083 vdd 5319 5323 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08082 5528 5323 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08081 vdd 4506 4081 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08080 4081 4515 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08079 vdd 4079 4081 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08078 4080 4081 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08077 vdd 5750 5747 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08076 5747 6212 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08075 vdd 5746 5747 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08074 5745 5747 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08073 2426 2498 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08072 5967 2499 2426 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08071 vdd 2517 5967 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08070 6244 6477 6246 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08069 6246 6974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08068 vdd 6714 6244 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08067 6245 6244 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08066 5317 5753 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08065 5322 5767 5317 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08064 vdd 6665 5322 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08063 vdd 3217 2503 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08062 2503 2506 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08061 2503 2501 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08060 vdd 2782 2503 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08059 2733 2503 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08058 5765 5998 5766 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08057 5764 5763 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08056 vdd 5764 5765 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08055 4085 4082 4084 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08054 4084 4083 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08053 vdd 5902 4085 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08052 4518 4085 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08051 6685 6688 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08050 vdd 6692 6685 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08049 1255 1333 1332 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08048 1254 1530 1255 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08047 vdd 1524 1254 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08046 3728 3560 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08045 3728 3947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08044 vdd 6423 3728 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08043 820 822 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08042 816 823 817 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08041 vdd 1191 816 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08040 821 823 820 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08039 819 824 821 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08038 vdd 818 819 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08037 818 821 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08036 817 824 818 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08035 vdd 817 1191 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08034 1191 817 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08033 vdd 3259 824 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08032 823 824 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08031 vdd 990 822 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08030 4564 5753 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08029 4701 5767 4564 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08028 vdd 4918 4701 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08027 914 968 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08026 vdd 965 914 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08025 790 1322 789 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08024 789 2746 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08023 vdd 3188 790 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08022 794 790 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08021 1217 1745 1216 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08020 1216 1989 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08019 vdd 1560 1217 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08018 1215 1217 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08017 1740 1967 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08016 vdd 1758 1740 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08015 946 1737 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08014 vdd 2506 946 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08013 5668 5915 5669 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08012 5669 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08011 vdd 6678 5669 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08010 5666 5668 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08009 5667 6637 5668 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08008 5669 6777 5667 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08007 3556 3379 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08006 3556 3947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08005 vdd 6423 3556 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08004 vdd 6186 5824 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08003 5824 6431 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08002 6843 5958 5824 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08001 5823 6182 6843 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08000 5824 6183 5823 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07999 3545 4082 3647 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07998 3544 4083 3545 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07997 vdd 3662 3544 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07996 3648 3647 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07995 1566 1564 1568 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07994 1567 1565 1566 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07993 vdd 1575 1567 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07992 2803 1568 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07991 5398 5954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07990 5489 5502 5398 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07989 vdd 5963 5489 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07988 4455 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07987 4455 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07986 vdd 5068 4455 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07985 5343 5272 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07984 5343 4737 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07983 vdd 5133 5343 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07982 2578 2399 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07981 vdd 2400 2578 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07980 827 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07979 1541 987 827 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07978 vdd 829 1541 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07977 5331 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07976 5331 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07975 vdd 5773 5331 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07974 3413 2610 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07973 vdd 2607 3413 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07972 1320 3217 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07971 1320 1687 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07970 vdd 1679 1320 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07969 6207 6893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07968 6207 6631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07967 vdd 6806 6207 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07966 5722 5723 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07965 6178 5721 5722 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07964 vdd 5948 6178 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07963 2790 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07962 2790 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07961 vdd 3818 2790 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07960 vdd 6440 2790 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07959 2384 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07958 2384 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07957 vdd 3818 2384 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07956 vdd 6440 2384 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07955 2625 3849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07954 2625 4088 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07953 vdd 4941 2625 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07952 858 1965 856 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07951 859 857 858 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07950 858 3229 859 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07949 856 1982 858 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07948 856 1389 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07947 vdd 3460 856 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07946 1918 2347 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07945 1918 3593 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07944 vdd 1688 1918 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07943 vdd 5478 5481 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07942 5481 5483 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07941 vdd 5485 5481 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07940 5932 5481 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07939 4888 4887 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07938 vdd 4889 4888 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07937 5036 4888 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07936 3642 3641 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07935 3640 3648 3642 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07934 vdd 3645 3640 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07933 4634 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07932 vdd 4634 4633 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07931 4632 4630 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07930 vdd 4632 4543 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07929 4543 4633 4629 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07928 4629 4634 4542 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07927 4580 6242 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_07926 vdd 4747 6242 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07925 6242 4747 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07924 4542 4627 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07923 4627 4629 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07922 vdd 6976 4627 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07921 4747 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07920 4747 4633 4580 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_07919 4627 4634 4747 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_07918 vdd 6680 6427 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07917 6427 6434 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07916 vdd 6919 6427 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07915 6426 6427 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07914 vdd 2742 2327 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07913 2327 2508 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07912 vdd 2507 2327 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07911 2325 2327 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07910 493 625 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07909 493 3193 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07908 vdd 624 493 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07907 vdd 3217 493 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07906 1226 1379 1227 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07905 1227 4748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07904 vdd 1576 1227 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07903 1224 1226 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07902 1225 1746 1226 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07901 1227 1745 1225 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07900 5403 5954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07899 5505 5502 5403 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07898 vdd 5742 5505 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07897 3705 4299 3866 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07896 3865 5157 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07895 vdd 3865 3705 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07894 vdd 5773 3303 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07893 3303 5349 3450 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07892 3452 3450 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07891 2035 2180 2034 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07890 2184 2182 2035 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07889 2035 2183 2184 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07888 2034 2193 2035 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07887 2034 2399 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07886 vdd 2799 2034 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07885 vdd 6434 3965 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07884 3965 6919 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07883 3964 5372 3965 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07882 3963 4217 3964 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07881 3965 5502 3963 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07880 2208 4299 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07879 vdd 5363 2208 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07878 944 1158 877 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07877 877 1289 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07876 vdd 946 944 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07875 943 944 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07874 4890 5954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07873 4889 5502 4890 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07872 vdd 5725 4889 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07871 2847 2848 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07870 2843 2850 2842 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07869 vdd 2852 2843 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07868 2846 2850 2847 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07867 2845 2849 2846 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07866 vdd 2844 2845 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07865 2844 2846 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07864 2842 2849 2844 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07863 vdd 2842 2852 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07862 2852 2842 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07861 vdd 3259 2849 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07860 2850 2849 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07859 vdd 2851 2848 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07858 vdd 6952 6239 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07857 6239 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07856 6239 6974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07855 vdd 6963 6239 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07854 6238 6239 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07853 vdd 4604 3786 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07852 3786 3795 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07851 vdd 4215 3786 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07850 3783 3786 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07849 vdd 328 77 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07848 77 81 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07847 vdd 214 77 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07846 478 77 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07845 2620 2622 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07844 vdd 2623 2620 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07843 3457 2620 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07842 2627 2628 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07841 vdd 2625 2627 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07840 2833 2627 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07839 2401 2399 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07838 vdd 2400 2401 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07837 4213 2401 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07836 2729 2728 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07835 vdd 2727 2729 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07834 2924 2729 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07833 5780 5781 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07832 5774 5782 5775 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07831 vdd 5773 5774 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07830 5779 5782 5780 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07829 5776 5783 5779 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07828 vdd 5777 5776 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07827 5777 5779 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07826 5775 5783 5777 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07825 vdd 5775 5773 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07824 5773 5775 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07823 vdd 6984 5783 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07822 5782 5783 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07821 vdd 5778 5781 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07820 2880 3074 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07819 2878 3075 3069 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07818 vdd 3263 2878 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07817 3073 3075 2880 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07816 2879 3076 3073 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07815 vdd 3070 2879 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07814 3070 3073 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07813 3069 3076 3070 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07812 vdd 3069 3263 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07811 3263 3069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07810 vdd 3259 3076 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07809 3075 3076 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07808 vdd 3262 3074 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07807 4924 5986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07806 4925 6214 4924 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07805 vdd 6591 4925 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07804 vdd 466 467 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07803 1304 571 465 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07802 465 466 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07801 465 467 1304 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07800 vdd 464 465 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07799 464 571 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07798 vdd 5749 5739 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07797 5739 5748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07796 5739 6850 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07795 vdd 6440 5739 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07794 5738 5739 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07793 vdd 5755 5535 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07792 5535 5538 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07791 5535 5540 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07790 vdd 5534 5535 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07789 5533 5535 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07788 6276 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07787 6348 6877 6276 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07786 vdd 6850 6348 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07785 5400 5496 5728 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07784 5495 5493 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07783 vdd 5495 5400 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07782 4571 4611 5127 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07781 4570 4612 4571 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07780 vdd 6422 4570 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07779 vdd 592 58 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07778 191 607 19 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07777 19 592 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07776 19 58 191 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07775 vdd 60 19 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07774 60 607 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07773 vdd 6694 6292 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07772 6292 6934 6430 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07771 5397 6173 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07770 5978 6172 5397 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07769 vdd 5964 5978 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07768 vdd 4696 3574 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07767 3574 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07766 3572 6727 3574 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07765 3571 3737 3572 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07764 3574 3738 3571 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07763 vdd 2487 2312 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07762 2320 2730 2313 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07761 2313 2487 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07760 2313 2312 2320 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07759 vdd 2311 2313 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07758 2311 2730 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07757 3166 5044 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07756 3165 5045 3166 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07755 vdd 3969 3165 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07754 5151 4954 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07753 vdd 4952 5151 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07752 5580 5569 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07751 vdd 5154 5580 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07750 4567 4704 4610 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07749 4566 4609 4567 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07748 vdd 5094 4566 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07747 523 1190 524 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07746 524 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07745 vdd 522 523 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07744 1346 523 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07743 4071 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07742 3836 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07741 4275 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07740 4501 4748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07739 2799 3263 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07738 3664 2852 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07737 vdd 4276 4269 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07736 4269 4941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07735 4269 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07734 vdd 4275 4269 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07733 5341 4269 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07732 vdd 1991 1043 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07731 1043 2352 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07730 1043 4094 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07729 vdd 5363 1043 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07728 1223 1043 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07727 907 1029 906 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07726 1221 5749 907 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07725 907 1031 1221 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07724 906 1232 907 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07723 906 1732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07722 vdd 1231 906 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07721 vdd 2782 2027 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07720 2027 2371 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07719 2057 2154 2027 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07718 2026 4673 2057 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07717 2027 4671 2026 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07716 6162 6161 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07715 6155 6163 6156 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07714 vdd 6740 6155 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07713 6158 6163 6162 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07712 6159 6164 6158 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07711 vdd 6157 6159 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07710 6157 6158 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07709 6156 6164 6157 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07708 vdd 6156 6740 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07707 6740 6156 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07706 vdd 6832 6164 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07705 6163 6164 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07704 vdd 6160 6161 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07703 vdd 4477 4459 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07702 4457 6186 4460 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07701 4458 6220 4457 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07700 4459 4456 4458 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07699 vdd 4212 4039 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07698 4040 5987 4042 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07697 4041 6188 4040 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07696 4039 4038 4041 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07695 5994 5556 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07694 vdd 5557 5994 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07693 5778 5564 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07692 vdd 5561 5778 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07691 5354 5348 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07690 vdd 5788 5354 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07689 3691 3792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07688 3795 3793 3691 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07687 vdd 3790 3795 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07686 3455 2408 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07685 vdd 2409 3455 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07684 3449 2836 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07683 vdd 2837 3449 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07682 863 3460 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07681 6469 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07680 6476 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07679 6921 6974 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07678 2455 3051 2610 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07677 2609 5893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07676 vdd 2609 2455 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07675 vdd 6616 5707 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07674 5951 5705 5706 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07673 5706 6616 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07672 5706 5707 5951 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07671 vdd 5704 5706 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07670 5704 5705 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07669 6830 6357 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07668 vdd 6841 6830 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07667 6017 6694 5851 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07666 5851 6015 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07665 vdd 6263 5851 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07664 6256 6017 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07663 5850 6013 6017 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07662 5851 6014 5850 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07661 6295 6682 6432 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07660 6293 6694 6295 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07659 6294 6480 6293 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07658 vdd 6934 6294 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07657 6431 6432 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07656 5025 5026 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07655 5025 6910 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07654 vdd 6806 5025 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07653 3614 4226 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07652 vdd 3613 3614 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07651 3588 4881 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07650 4020 4880 3588 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07649 vdd 5964 4020 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07648 4705 5767 4568 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07647 4568 5753 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07646 vdd 5026 4705 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07645 4704 4705 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07644 199 607 198 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07643 198 592 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07642 vdd 603 199 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07641 196 199 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07640 4258 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07639 4258 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07638 vdd 5992 4258 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07637 3629 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07636 3629 4726 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07635 vdd 5773 3629 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07634 2836 2622 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07633 vdd 2623 2836 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07632 897 1194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07631 1542 1190 897 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07630 vdd 1002 1542 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07629 6209 6211 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07628 6209 6424 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07627 vdd 6208 6209 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07626 1208 2139 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07625 vdd 2138 1208 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07624 vdd 2946 2277 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07623 2277 2950 2324 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07622 2356 2324 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07621 3831 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07620 3831 4265 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07619 vdd 5773 3831 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07618 6715 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07617 vdd 6952 6715 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07616 vdd 4524 865 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07615 865 4748 2125 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07614 1022 1218 902 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07613 902 1231 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07612 vdd 1732 1022 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07611 1946 1022 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07610 1232 2625 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07609 1232 1236 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07608 vdd 1582 1232 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07607 5404 5805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07606 5508 5756 5404 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07605 vdd 5670 5508 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07604 5295 5804 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07603 vdd 6265 5294 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07602 vdd 5309 5296 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07601 5293 5309 5295 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07600 5294 5296 5293 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07599 5292 5293 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07598 4108 5963 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07597 vdd 5902 4107 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07596 vdd 5309 4204 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07595 4203 5309 4108 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07594 4107 4204 4203 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07593 4200 4203 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07592 4104 6187 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07591 vdd 5372 4103 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07590 vdd 5309 4195 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07589 4192 5309 4104 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07588 4103 4195 4192 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07587 4191 4192 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07586 vdd 6011 4511 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07585 4511 6690 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07584 vdd 4509 4511 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07583 4510 4511 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07582 207 328 208 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07581 208 1900 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07580 vdd 2161 208 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07579 480 207 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07578 206 319 207 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07577 208 320 206 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07576 1177 2331 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07575 1177 1175 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07574 vdd 1176 1177 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07573 1174 2746 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07572 1175 1322 1174 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07571 vdd 3188 1175 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07570 5346 5341 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07569 vdd 5349 5346 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07568 4254 4726 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07567 vdd 5773 4254 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07566 1727 2782 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07565 1727 2506 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07564 vdd 2371 1727 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07563 2117 1953 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07562 2117 1553 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07561 vdd 2194 2117 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07560 vdd 3836 2117 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07559 vdd 4171 3952 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07558 3952 3951 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07557 vdd 5666 3952 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07556 3950 3952 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07555 vdd 3766 3557 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07554 3557 3556 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07553 vdd 3957 3557 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07552 3555 3557 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07551 5311 5742 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07550 vdd 6727 5307 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07549 vdd 5309 5310 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07548 5308 5309 5311 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07547 5307 5310 5308 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07546 5306 5308 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07545 5813 6190 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07544 6588 6191 5813 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07543 vdd 5927 6588 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07542 vdd 5877 4742 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07541 4742 5349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07540 vdd 6440 4742 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07539 5548 4742 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07538 vdd 1151 1150 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07537 2913 1280 1152 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07536 1152 1151 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07535 1152 1150 2913 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07534 vdd 1149 1152 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07533 1149 1280 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07532 6221 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07531 6221 4941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07530 vdd 4276 6221 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07529 vdd 4275 6221 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07528 4281 4286 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07527 4281 4941 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07526 vdd 4276 4281 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07525 vdd 4275 4281 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07524 2354 2350 2351 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07523 2353 2512 2354 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07522 2354 2534 2353 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07521 2351 2521 2354 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07520 2351 2349 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07519 vdd 2520 2351 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07518 1876 4239 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07517 1876 1732 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07516 vdd 1218 1876 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07515 vdd 4748 1876 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07514 1209 4239 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07513 1209 2194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07512 vdd 1953 1209 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07511 vdd 3836 1209 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07510 4096 5272 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07509 vdd 4094 4095 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07508 vdd 5893 4098 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07507 4097 5893 4096 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07506 4095 4098 4097 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07505 4093 4097 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07504 vdd 1695 1697 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07503 1697 1925 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07502 vdd 1694 1697 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07501 1944 1697 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07500 340 494 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07499 vdd 2314 340 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07498 488 340 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07497 vdd 4258 4255 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07496 4255 5551 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07495 4255 4253 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07494 vdd 4254 4255 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07493 4257 4255 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07492 2140 2139 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07491 vdd 2138 2140 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07490 2981 2140 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07489 5314 5756 5313 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07488 5313 5805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07487 vdd 6665 5314 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07486 5312 5314 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07485 5379 5433 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07484 5377 5434 5426 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07483 vdd 5524 5377 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07482 5430 5434 5379 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07481 5378 5435 5430 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07480 vdd 5428 5378 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07479 5428 5430 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07478 5426 5435 5428 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07477 vdd 5426 5524 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07476 5524 5426 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07475 vdd 6580 5435 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07474 5434 5435 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07473 vdd 5431 5433 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07472 6283 6388 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07471 6281 6387 6381 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07470 vdd 6874 6281 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07469 6385 6387 6283 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07468 6282 6389 6385 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07467 vdd 6382 6282 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07466 6382 6385 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07465 6381 6389 6382 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07464 vdd 6381 6874 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07463 6874 6381 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07462 vdd 6832 6389 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07461 6387 6389 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07460 vdd 6384 6388 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07459 vdd 5245 5001 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07458 5019 5244 4966 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07457 4966 5245 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07456 4966 5001 5019 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07455 vdd 4999 4966 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07454 4999 5244 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07453 1249 1312 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07452 2997 1313 1249 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07451 vdd 1661 2997 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07450 1025 5748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07449 vdd 6440 1025 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07448 1031 1025 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07447 4897 3573 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07446 5064 3979 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07445 5299 3972 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07444 4696 3759 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07443 6956 6963 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07442 1934 3793 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07441 vdd 2352 1934 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07440 2331 1934 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07439 vdd 2161 1881 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07438 1881 1900 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07437 1880 1884 1881 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07436 1879 1888 1880 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07435 1881 2304 1879 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07434 874 938 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07433 936 943 874 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07432 vdd 1876 936 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07431 6199 6198 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07430 6193 6201 6194 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07429 vdd 6571 6193 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07428 6200 6201 6199 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07427 6195 6202 6200 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07426 vdd 6196 6195 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07425 6196 6200 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07424 6194 6202 6196 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07423 vdd 6194 6571 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07422 6571 6194 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07421 vdd 6984 6202 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07420 6201 6202 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07419 vdd 6197 6198 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07418 3961 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07417 3962 6877 3961 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07416 vdd 4918 3962 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07415 vdd 6876 6760 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07414 6760 6877 6791 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07413 3612 4671 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07412 3613 4673 3612 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07411 vdd 5964 3613 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07410 1529 3210 1528 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07409 1528 1534 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07408 vdd 2534 1529 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07407 1527 1529 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07406 6436 6714 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07405 vdd 6952 6436 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07404 6434 6436 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07403 4145 4282 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_07402 6000 4285 4145 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_07401 4144 4280 6000 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_07400 vdd 4281 4144 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_07399 5134 6242 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07398 4441 2979 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07397 4687 3190 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07396 4438 3403 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07395 4205 3395 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07394 vdd 2542 1932 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07393 1932 3208 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07392 1932 1931 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07391 vdd 1933 1932 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07390 2535 1932 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07389 vdd 6890 6884 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07388 6883 6885 6770 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07387 6770 6890 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07386 6770 6884 6883 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07385 vdd 6880 6770 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07384 6880 6885 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07383 vdd 5749 5083 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07382 5083 5748 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07381 5083 6820 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07380 vdd 6440 5083 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07379 5084 5083 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07378 2038 2202 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_07377 4079 2196 2038 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_07376 2037 2195 4079 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_07375 vdd 2194 2037 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_07374 vdd 6917 5768 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07373 5768 6921 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07372 vdd 6963 5768 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07371 5767 5768 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07370 3292 3792 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07369 4015 3793 3292 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07368 vdd 3421 4015 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07367 vdd 1737 1245 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07366 1245 2506 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07365 1292 1483 1245 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07364 1244 1645 1292 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07363 1245 1492 1244 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07362 6336 6169 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07361 vdd 6144 6336 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07360 873 1000 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07359 871 924 998 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07358 vdd 1002 871 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07357 923 924 873 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07356 872 925 923 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07355 vdd 921 872 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07354 921 923 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07353 998 925 921 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07352 vdd 998 1002 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07351 1002 998 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07350 vdd 3259 925 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07349 924 925 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07348 vdd 1001 1000 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07347 4904 4906 5504 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07346 4905 4903 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07345 vdd 4905 4904 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07344 4910 5297 4909 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07343 4908 5084 4910 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07342 vdd 4911 4908 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07341 2383 2381 2382 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07340 2380 2379 2383 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07339 vdd 3015 2380 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07338 1038 1965 853 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07337 853 1982 1038 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07336 vdd 857 853 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07335 853 3229 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07334 2300 2319 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07333 2301 2483 2300 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07332 vdd 2479 2301 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07331 3553 3376 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07330 3553 3947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07329 vdd 6423 3553 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07328 4662 6877 4550 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07327 4550 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07326 vdd 4918 4662 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07325 4854 4662 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07324 1924 2340 1925 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07323 1923 2129 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07322 vdd 1923 1924 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07321 2740 3572 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07320 vdd 2944 2740 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07319 1921 2534 1922 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07318 1922 2521 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07317 vdd 2512 1922 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07316 2336 1921 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07315 1920 1918 1921 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07314 1922 1919 1920 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07313 3720 3382 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07312 3720 3947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07311 vdd 6423 3720 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07310 4953 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07309 4953 4523 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07308 vdd 5144 4953 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07307 1329 2331 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07306 1329 1323 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07305 vdd 1186 1329 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07304 1394 3664 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07303 1394 2352 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07302 vdd 4094 1394 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07301 3737 1214 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07300 vdd 1215 3737 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07299 2944 3186 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07298 vdd 5742 2944 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07297 1908 3391 1911 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07296 1907 2333 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07295 vdd 1907 1908 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07294 3289 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07293 3595 3414 3289 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07292 vdd 5372 3595 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07291 6410 6906 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07290 6410 6631 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07289 vdd 6806 6410 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07288 5507 5504 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07287 vdd 5505 5507 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07286 5975 5507 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07285 4950 5132 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07284 vdd 5127 4950 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07283 5561 4950 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07282 5344 5343 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07281 vdd 5342 5344 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07280 5557 5344 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07279 vdd 2993 2781 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07278 2781 2990 2780 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_07277 2778 2780 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07276 851 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07275 851 860 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07274 vdd 2830 851 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07273 vdd 6440 851 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07272 686 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07271 686 1385 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07270 vdd 2830 686 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07269 vdd 6440 686 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07268 4720 4947 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07267 4720 4722 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07266 vdd 4731 4720 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07265 6852 6877 6739 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07264 6739 6876 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07263 vdd 6850 6852 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07262 6851 6852 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07261 6769 6866 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07260 6869 6875 6769 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07259 vdd 6867 6869 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07258 6396 6648 6286 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07257 6286 6791 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07256 vdd 6678 6286 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07255 6393 6396 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07254 6285 6637 6396 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07253 6286 6883 6285 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07252 vdd 6801 6805 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07251 6805 6808 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07250 vdd 6802 6805 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07249 6800 6805 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07248 3237 4083 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07247 3236 4082 3237 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07246 vdd 5272 3236 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07245 3015 5116 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07244 3015 3227 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07243 vdd 3816 3015 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07242 vdd 3218 3015 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07241 vdd 4748 2392 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07240 vdd 4235 2391 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07239 2392 2391 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07238 vdd 5068 4901 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07237 4901 5102 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07236 4901 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07235 vdd 5262 4901 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07234 4899 4901 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07233 vdd 6885 6872 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07232 6872 6893 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07231 vdd 6906 6872 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07230 6870 6872 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07229 3852 3853 3702 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07228 3702 5341 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07227 vdd 5575 3702 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07226 6876 3852 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07225 3701 3849 3852 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07224 3702 3856 3701 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07223 2772 5959 2774 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07222 2774 2773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07221 vdd 4438 2774 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07220 2770 2772 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07219 2771 3199 2772 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07218 2774 3618 2771 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07217 vdd 4094 1053 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07216 1053 4524 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07215 vdd 5363 1053 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07214 1779 1053 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07213 2041 2629 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07212 2411 2418 2041 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07211 vdd 2208 2411 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07210 vdd 2102 1892 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07209 1892 2095 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07208 1891 2485 1892 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07207 1890 2319 1891 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07206 1892 2320 1890 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07205 vdd 6449 6009 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07204 6009 6448 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07203 vdd 6917 6009 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07202 6013 6009 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07201 4579 5773 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07200 4745 5575 4579 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07199 vdd 5889 4745 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07198 3060 2412 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07197 vdd 2406 3060 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07196 vdd 1031 904 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07195 904 5749 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07194 1214 1732 904 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07193 903 1231 1214 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07192 904 1218 903 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07191 1585 2799 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07190 1586 1587 1585 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07189 1584 2198 1586 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07188 vdd 2409 1584 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07187 1583 1586 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07186 1489 1641 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07185 vdd 1893 1489 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07184 1488 1489 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07183 1290 1492 1243 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07182 1243 1645 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07181 vdd 1483 1290 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07180 1289 1290 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07179 2862 2934 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07178 2860 2933 2928 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07177 vdd 3560 2860 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07176 2931 2933 2862 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07175 2861 2935 2931 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07174 vdd 2929 2861 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07173 2929 2931 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07172 2928 2935 2929 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07171 vdd 2928 3560 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07170 3560 2928 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07169 vdd 3160 2935 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07168 2933 2935 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07167 vdd 3563 2934 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07166 vdd 1235 1230 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07165 1230 1985 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07164 vdd 1579 1230 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07163 1229 1230 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07162 905 1231 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07161 2506 1218 905 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07160 vdd 1732 2506 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07159 2738 3172 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07158 vdd 2936 2738 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07157 2737 2738 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07156 5356 5358 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07155 5350 5357 5351 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07154 vdd 5349 5350 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07153 5355 5357 5356 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07152 5353 5360 5355 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07151 vdd 5352 5353 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07150 5352 5355 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07149 5351 5360 5352 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07148 vdd 5351 5349 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07147 5349 5351 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07146 vdd 6984 5360 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07145 5357 5360 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07144 vdd 5354 5358 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07143 vdd 6870 6865 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07142 6866 6861 6768 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07141 6768 6870 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07140 6768 6865 6866 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07139 vdd 6863 6768 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07138 6863 6861 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07137 vdd 196 62 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07136 305 470 20 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07135 20 196 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07134 20 62 305 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07133 vdd 64 20 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07132 64 470 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07131 vdd 5039 4694 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07130 4694 5877 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07129 4694 5992 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07128 vdd 6440 4694 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07127 4695 4694 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07126 vdd 493 215 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07125 215 787 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07124 vdd 2314 215 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07123 319 215 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07122 497 987 498 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07121 498 986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07120 vdd 500 497 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07119 919 497 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07118 vdd 1971 1970 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07117 1970 2610 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07116 vdd 2607 1970 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07115 1968 1970 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07114 3169 5902 3170 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07113 3170 3740 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07112 vdd 5064 3170 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07111 3167 3169 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07110 3168 3737 3169 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07109 3170 3738 3168 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07108 vdd 2511 2332 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07107 2332 2512 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07106 vdd 2331 2332 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07105 2518 2332 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07104 vdd 4748 3646 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07103 3646 3662 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07102 3645 5372 3646 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07101 3644 4083 3645 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07100 3646 4082 3644 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07099 4998 5165 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07098 4996 5166 5159 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07097 vdd 5157 4996 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07096 5162 5166 4998 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07095 4997 5167 5162 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07094 vdd 5160 4997 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07093 5160 5162 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07092 5159 5167 5160 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07091 vdd 5159 5157 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07090 5157 5159 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07089 vdd 6984 5167 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07088 5166 5167 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07087 vdd 5164 5165 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07086 3291 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07085 3416 3414 3291 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07084 vdd 5902 3416 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07083 1999 2169 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07082 1997 2067 2167 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07081 vdd 2583 1997 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07080 2065 2067 1999 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07079 1998 2068 2065 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07078 vdd 2064 1998 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07077 2064 2065 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07076 2167 2068 2064 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07075 vdd 2167 2583 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07074 2583 2167 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07073 vdd 3259 2068 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07072 2067 2068 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07071 vdd 2582 2169 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07070 5369 5570 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07069 vdd 5788 5369 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07068 3288 3413 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07067 3589 3414 3288 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07066 vdd 5243 3589 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07065 3563 3727 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07064 vdd 3971 3563 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07063 6152 6151 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07062 6146 6153 6145 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07061 vdd 6820 6146 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07060 6148 6153 6152 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07059 6147 6154 6148 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07058 vdd 6149 6147 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07057 6149 6148 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07056 6145 6154 6149 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07055 vdd 6145 6820 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07054 6820 6145 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07053 vdd 6832 6154 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07052 6153 6154 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07051 vdd 6150 6151 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07050 5337 5125 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07049 vdd 6447 5337 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07048 1657 2314 1603 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07047 1603 2356 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07046 vdd 2111 1603 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07045 1655 1657 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07044 1602 3740 1657 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07043 1603 2553 1602 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07042 2440 3199 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07041 2546 3618 2440 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07040 vdd 5725 2546 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07039 403 2194 295 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07038 295 2195 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07037 vdd 1033 403 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07036 402 403 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07035 vdd 2320 1898 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07034 2107 1905 1899 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07033 1899 2320 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07032 1899 1898 2107 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07031 vdd 1897 1899 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07030 1897 1905 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07029 6384 6178 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07028 vdd 6180 6384 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07027 4465 4610 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07026 vdd 5088 4465 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07025 5095 6214 4989 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07024 4989 5986 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07023 vdd 6820 5095 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07022 5094 5095 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07021 5527 5767 5388 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07020 5388 5753 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07019 vdd 5524 5527 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07018 5525 5527 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_07017 4253 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07016 4253 4265 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07015 vdd 5992 4253 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07014 vdd 5144 2410 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07013 2410 5359 2409 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_07012 1746 1991 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07011 vdd 1779 1746 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07010 6652 6400 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07009 vdd 6398 6652 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07008 3816 5575 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07007 3816 5068 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07006 vdd 5069 3816 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07005 5116 6440 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07004 5116 4726 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07003 vdd 5992 5116 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07002 3218 5069 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07001 3218 4062 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07000 vdd 5068 3218 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06999 1582 4089 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06998 vdd 2412 1582 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06997 1231 1582 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06996 vdd 2625 1231 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06995 2348 3199 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_06994 2347 3618 2348 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_06993 vdd 6187 2347 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_06992 2936 3186 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06991 vdd 5963 2936 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06990 2736 3172 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06989 vdd 2936 2736 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06988 6592 6616 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06987 vdd 6591 6592 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06986 6590 6592 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_06985 vdd 1708 1610 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_06984 1610 1706 1707 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_06983 2052 1707 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_06982 1945 2553 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06981 vdd 2356 1945 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06980 81 1151 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06979 81 212 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06978 vdd 772 81 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06977 209 1151 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06976 209 86 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06975 vdd 772 209 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06974 6724 6984 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06973 vdd 6724 6723 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06972 6721 6967 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06971 vdd 6721 6722 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06970 6722 6723 6720 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06969 6720 6724 6719 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06968 6716 6952 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_06967 vdd 6717 6952 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_06966 6952 6717 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_06965 6719 6718 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06964 6718 6720 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06963 vdd 6976 6718 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06962 6717 6976 vdd vdd  sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06961 6717 6723 6716 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_06960 6718 6724 6717 vdd sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_06959 6855 6876 6854 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06958 6854 6877 6855 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06957 vss 6874 6854 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06956 155 615 156 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06955 156 493 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06954 214 2314 155 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06953 90 787 89 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06952 89 493 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06951 210 2314 90 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06950 vss 6698 6917 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06949 6698 6714 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06948 6917 6952 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06947 6443 6694 6444 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06946 6444 6934 6443 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06945 vss 6442 6444 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06944 6449 6443 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06943 4035 4275 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06942 vss 4032 4035 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06941 4035 4708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06940 vss 6224 4035 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06939 4228 4035 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06938 1039 2195 745 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06937 745 2194 1039 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06936 vss 1033 745 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06935 4361 5068 4362 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06934 4362 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06933 4360 5069 4361 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06932 4447 4448 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06931 4448 5272 4360 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06930 6819 6817 6818 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06929 6818 6821 6819 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06928 vss 6867 6818 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06927 6511 6740 6512 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06926 6512 6839 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06925 6510 6820 6511 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06924 6616 6617 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06923 6617 6850 6510 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06922 vss 1329 1083 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06921 1083 1339 1180 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06920 1326 1180 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06919 5587 5679 5671 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06918 vss 5670 5587 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06917 5673 5674 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06916 vss 5673 5588 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06915 5671 5678 5673 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06914 5670 5671 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06913 vss 5671 5670 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06912 5588 5678 5674 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06911 5674 5679 5589 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06910 vss 6580 5679 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06909 5678 5679 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06908 vss 5682 5676 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06907 5589 5676 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06906 4161 4162 4160 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06905 vss 4918 4161 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06904 4159 4649 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06903 4160 4158 4159 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06902 vss 4649 4162 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06901 4158 4918 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06900 151 209 152 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06899 152 489 211 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06898 vss 210 151 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06897 477 211 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06896 6076 6919 6075 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06895 6075 6430 6217 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06894 vss 6917 6076 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06893 6216 6217 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06892 vss 1360 1097 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06891 1097 1210 1211 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06890 1322 1211 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06889 vss 263 170 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06888 170 265 262 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06887 395 262 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06886 vss 3183 3088 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06885 3088 3184 3181 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06884 3182 3181 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06883 vss 2525 2527 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06882 2527 2526 2528 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06881 2752 2528 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06880 6533 6658 6650 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06879 vss 6885 6533 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06878 6651 6655 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06877 vss 6651 6534 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06876 6650 6657 6651 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06875 6885 6650 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06874 vss 6650 6885 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06873 6534 6657 6655 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06872 6655 6658 6535 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06871 vss 6984 6658 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06870 6657 6658 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06869 vss 6652 6656 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06868 6535 6656 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06867 3000 2999 3001 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06866 3001 2997 3000 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06865 vss 2998 3001 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06864 4737 3000 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06863 vss 2834 2697 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06862 2697 2833 2835 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06861 2837 2835 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06860 vss 6917 5990 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06859 5990 6219 5989 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06858 5987 5989 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06857 5763 5805 5619 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06856 5619 5756 5763 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06855 vss 6807 5619 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06854 3911 4015 3910 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06853 3910 5305 4017 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06852 vss 4016 3911 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06851 4014 4017 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06850 3733 6434 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06849 3734 6919 3733 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06848 3732 5262 3734 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06847 vss 4217 3732 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06846 3732 5502 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06845 4581 4586 4664 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06844 vss 4914 4581 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06843 4582 4584 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06842 vss 4582 4583 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06841 4664 4585 4582 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06840 4914 4664 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06839 vss 4664 4914 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06838 4583 4585 4584 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06837 4584 4586 4667 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06836 vss 6580 4586 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06835 4585 4586 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06834 vss 4665 4666 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06833 4667 4666 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06832 vss 2046 2508 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06831 2508 2045 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06830 vss 2044 2508 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06829 4251 4250 4252 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06828 4252 4491 4251 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06827 vss 5349 4252 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06826 4572 4251 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06825 3931 4941 3932 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06824 3932 4287 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06823 3930 4286 3931 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06822 4265 4070 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06821 4070 4524 3930 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06820 2491 3741 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06819 2490 2739 2491 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06818 vss 2733 2490 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06817 2489 2490 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06816 5220 5761 5221 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06815 5221 5327 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06814 5219 5985 5220 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06813 5762 5328 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06812 5328 5326 5219 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06811 vss 5334 5033 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06810 5054 5033 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06809 vss 5033 5054 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06808 vss 5033 5054 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06807 5054 5033 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06806 vss 5334 1571 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06805 3259 1571 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06804 vss 1571 3259 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06803 vss 1571 3259 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06802 3259 1571 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06801 vss 5334 1570 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06800 1569 1570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06799 vss 1570 1569 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06798 vss 1570 1569 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06797 1569 1570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06796 vss 5334 1371 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06795 1370 1371 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06794 vss 1371 1370 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06793 vss 1371 1370 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06792 1370 1371 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06791 vss 5334 1512 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06790 3160 1512 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06789 vss 1512 3160 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06788 vss 1512 3160 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06787 3160 1512 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06786 vss 5334 1511 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06785 1510 1511 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06784 vss 1511 1510 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06783 vss 1511 1510 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06782 1510 1511 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06781 vss 5334 1316 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06780 1315 1316 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06779 vss 1316 1315 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06778 vss 1316 1315 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06777 1315 1316 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06776 6888 6891 6889 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06775 vss 6886 6888 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06774 6892 6890 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06773 6889 6887 6892 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06772 vss 6890 6891 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06771 6887 6886 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06770 vss 6877 6675 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06769 6675 6876 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06768 vss 6903 6675 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06767 1763 4089 1764 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06766 1764 2352 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06765 1761 4087 1763 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06764 1760 1762 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06763 1762 4299 1761 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06762 2970 2976 2971 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06761 2967 2978 2970 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06760 2979 2970 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06759 vss 2970 2979 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06758 2974 2975 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06757 vss 2977 2975 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06756 2976 2978 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06755 vss 3160 2978 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06754 2969 2973 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06753 2971 6976 2969 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06752 2973 2978 2974 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06751 2972 2976 2973 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06750 vss 2971 2972 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06749 vss 2979 2968 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06748 2968 6976 2967 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06747 4177 4176 4178 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06746 4178 6600 4177 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06745 vss 6601 4178 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06744 4397 4177 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06743 6126 6876 6031 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06742 6031 6877 6126 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06741 vss 6665 6031 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06740 6127 6126 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06739 5107 5106 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06738 5168 5104 5107 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06737 5755 5753 5618 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06736 5618 5767 5755 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06735 vss 6807 5618 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06734 5265 5044 5032 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06733 5032 5045 5265 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06732 vss 5965 5032 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06731 5879 5972 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06730 6197 5969 5879 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06729 2047 2508 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06728 2048 2507 2047 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06727 3466 6423 3465 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06726 3465 3947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06725 3550 3546 3466 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06724 vss 399 168 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06723 168 261 260 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06722 830 260 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06721 vss 4501 4274 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06720 vss 4273 4274 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06719 4274 4275 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06718 4512 4274 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06717 6877 6469 4721 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06716 4721 4733 6877 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06715 vss 4731 4721 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06714 570 579 572 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06713 572 569 570 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06712 vss 2727 572 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06711 1313 570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06710 3491 4909 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06709 3592 3788 3491 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06708 4941 4299 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06707 vss 5157 4941 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06706 4941 2852 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06705 vss 3460 4941 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06704 1366 1365 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06703 2379 3226 1366 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06702 1731 1732 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06701 1730 1760 1731 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06700 1812 2139 1813 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06699 1813 1944 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06698 5792 2138 1812 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06697 6100 6714 6101 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06696 6101 6440 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06695 6099 6952 6100 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06694 6477 6963 6099 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06693 vss 5880 5984 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06692 5984 6216 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06691 5983 5984 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06690 3471 3550 3470 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06689 3470 3964 3551 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06688 vss 5003 3471 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06687 3549 3551 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06686 3922 4072 3923 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06685 3923 4257 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06684 4066 4953 3922 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06683 3425 3622 3426 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06682 3426 3621 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06681 5309 3424 3425 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06680 5862 5723 5594 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06679 5594 5721 5862 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06678 vss 5965 5594 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06677 4375 4510 4376 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06676 4376 4502 4504 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06675 vss 4503 4375 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06674 4618 4504 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06673 2134 2135 2137 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06672 2137 2136 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06671 2345 2331 2134 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06670 1454 1562 1455 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06669 1455 1744 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06668 1453 2173 1454 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06667 5748 1563 1453 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06666 2389 4235 2252 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06665 vss 4748 2390 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06664 2252 2390 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06663 vss 5363 1045 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06662 1045 1991 1044 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06661 1953 1044 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06660 4789 5068 4790 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06659 4790 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06658 4788 5069 4789 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06657 4906 4907 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06656 4907 6727 4788 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06655 2145 2142 2143 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06654 2143 2544 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06653 2144 2532 2145 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06652 1494 1885 1409 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06651 1409 1891 1494 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06650 vss 1882 1409 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06649 1492 1494 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06648 4841 6791 4758 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06647 4757 5011 4841 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06646 4758 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06645 4838 4841 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06644 vss 6637 4757 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06643 4757 4839 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06642 5119 5115 5120 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06641 5120 5770 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06640 5117 5331 5119 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06639 6910 5118 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06638 5118 5116 5117 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06637 vss 4477 3420 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06636 vss 5987 3420 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06635 3420 4456 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06634 3740 3420 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06633 1642 3217 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06632 1641 2535 1642 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06631 vss 1640 1641 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06630 5856 6172 5590 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06629 5590 6173 5856 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06628 vss 5927 5590 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06627 vss 1694 1693 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06626 1693 1925 1692 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06625 2763 1692 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06624 vss 2144 2131 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06623 2131 2128 2130 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06622 2340 2130 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06621 vss 2782 1805 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06620 1805 2501 1901 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06619 1900 1901 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06618 3080 3162 3153 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06617 vss 3379 3080 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06616 3156 3158 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06615 vss 3156 3081 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06614 3153 3161 3156 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06613 3379 3153 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06612 vss 3153 3379 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06611 3081 3161 3158 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06610 3158 3162 3082 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06609 vss 3160 3162 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06608 3161 3162 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06607 vss 3163 3159 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06606 3082 3159 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06605 6776 6779 6777 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06604 vss 6905 6776 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06603 6780 6778 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06602 6777 6775 6780 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06601 vss 6778 6779 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06600 6775 6905 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06599 1927 2124 1851 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06598 1850 2122 1927 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06597 1851 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06596 2128 1927 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06595 vss 1929 1850 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06594 1850 2532 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06593 3430 3792 3105 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06592 3105 3793 3430 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06591 vss 3434 3105 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06590 4291 4298 4290 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06589 vss 4299 4291 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06588 4292 4293 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06587 vss 4292 4294 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06586 4290 4297 4292 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06585 4299 4290 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06584 vss 4290 4299 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06583 4294 4297 4293 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06582 4293 4298 4295 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06581 vss 6984 4298 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06580 4297 4298 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06579 vss 4300 4296 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06578 4295 4296 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06577 vss 1338 1339 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06576 1339 1343 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06575 vss 1533 1339 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06574 4243 5349 4245 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06573 4245 5341 4244 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06572 vss 6440 4243 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06571 4477 4244 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06570 862 863 746 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06569 746 1390 862 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06568 vss 3263 746 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06567 860 862 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06566 1352 2194 1351 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06565 1351 1553 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06564 1350 1953 1352 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06563 2122 1349 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06562 1349 3836 1350 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06561 2103 2511 2105 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06560 2104 2314 2103 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06559 2105 2111 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06558 2102 2103 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06557 vss 3740 2104 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06556 2104 2512 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06555 3907 5500 3906 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06554 3906 4009 4011 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06553 vss 4010 3907 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06552 4008 4011 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06551 5699 6876 5597 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06550 5597 6877 5699 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06549 vss 6591 5597 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06548 6413 6182 5612 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06547 5612 6183 6413 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06546 vss 5742 5612 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06545 3806 3819 3807 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06544 3807 3805 3806 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06543 vss 5102 3807 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06542 4611 3806 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06541 vss 5502 4471 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06540 4471 4052 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06539 vss 4048 4471 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06538 2250 5069 2251 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06537 2251 2807 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06536 2249 5773 2250 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06535 2387 2388 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06534 2388 6440 2249 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06533 2515 2511 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06532 vss 2512 2515 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06531 2515 2513 3183 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06530 3183 2514 2515 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06529 3127 3555 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06528 3163 3736 3127 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06527 3396 3350 3344 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06526 3341 3349 3396 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06525 3403 3396 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06524 vss 3396 3403 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06523 3346 3348 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06522 vss 3397 3348 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06521 3350 3349 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06520 vss 5054 3349 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06519 3343 3347 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06518 3344 6976 3343 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06517 3347 3349 3346 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06516 3345 3350 3347 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06515 vss 3344 3345 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06514 vss 3403 3342 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06513 3342 6976 3341 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06512 41 120 115 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06511 vss 392 41 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06510 42 43 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06509 vss 42 44 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06508 115 45 42 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06507 392 115 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06506 vss 115 392 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06505 44 45 43 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06504 43 120 118 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06503 vss 3259 120 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06502 45 120 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06501 vss 243 119 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06500 118 119 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06499 5182 6806 5181 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06498 5181 6910 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06497 5261 5524 5182 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06496 vss 6480 6012 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06495 6012 6682 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06494 6464 6012 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06493 3505 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06492 3622 4233 3505 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06491 1506 2946 1418 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06490 1418 2950 1506 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06489 vss 2111 1418 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06488 1505 1506 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06487 1361 2799 1362 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06486 1362 4051 1361 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06485 vss 3813 1362 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06484 1360 1361 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06483 5534 5112 4808 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06482 4808 5113 5534 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06481 vss 4937 4808 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06480 3126 3552 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06479 3152 3165 3126 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06478 vss 6182 6631 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06477 6631 6188 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06476 vss 6183 6631 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06475 4863 4857 4764 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06474 4764 4859 4863 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06473 vss 6867 4764 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06472 6602 6603 6503 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06471 6503 6600 6602 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06470 vss 6601 6503 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06469 6801 6602 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06468 916 1517 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06467 917 1518 916 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06466 1331 1339 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06465 1330 1329 1331 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06464 1653 3740 1654 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06463 1654 2553 1653 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06462 vss 2314 1654 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06461 1652 1653 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06460 2679 5069 2680 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06459 2680 2807 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06458 3814 5992 2679 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06457 2696 2833 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06456 3456 2834 2696 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06455 2042 2299 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06454 2303 2489 2042 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06453 2219 2306 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06452 2307 2492 2219 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06451 vss 5499 5500 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06450 5499 5498 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06449 5500 5510 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06448 5462 6423 5463 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06447 5463 6374 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06446 5461 6375 5462 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06445 5700 5501 5461 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06444 6066 6204 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06443 6900 6203 6066 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06442 4768 6806 4769 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06441 4769 6910 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06440 4866 4914 4768 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06439 308 598 309 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06438 309 307 308 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06437 vss 470 309 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06436 588 308 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06435 2075 2628 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06434 2194 2625 2075 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06433 6823 6876 6822 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06432 6822 6877 6823 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06431 vss 6820 6822 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06430 6821 6823 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06429 6419 6417 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06428 6914 6418 6419 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06427 vss 5489 5491 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06426 5491 5490 5492 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06425 6176 5492 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06424 vss 5140 5143 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06423 5143 5141 5142 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06422 5570 5142 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06421 vss 5773 4337 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06420 4337 5341 4498 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06419 4497 4498 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06418 3913 4461 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06417 4021 4020 3913 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06416 1666 1667 1668 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06415 1668 1676 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06414 1670 2331 1666 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06413 3812 5069 3815 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06412 3815 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06411 3813 3818 3812 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06410 6519 6629 6518 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06409 6518 6819 6630 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06408 vss 6627 6519 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06407 6628 6630 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06406 5476 5955 5475 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06405 5475 5867 5477 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06404 vss 5485 5476 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06403 5474 5477 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06402 5922 5919 5921 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06401 5921 6129 5920 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06400 vss 5925 5922 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06399 5918 5920 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06398 1435 1541 1434 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06397 1434 2986 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06396 1433 2550 1435 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06395 2512 1542 1433 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06394 5188 6423 5189 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06393 5189 6374 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06392 5187 6375 5188 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06391 5269 5268 5187 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06390 6546 6691 6547 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06389 6547 6692 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06388 6545 6695 6546 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06387 6696 6693 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06386 6693 6921 6545 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06385 1342 1340 1341 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06384 1341 3408 1342 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06383 vss 2521 1341 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06382 1699 1342 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06381 327 331 328 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06380 vss 779 327 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06379 330 488 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06378 328 329 330 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06377 vss 488 331 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06376 329 779 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06375 vss 4456 4223 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06374 4223 4477 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06373 5300 4223 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06372 vss 2838 4088 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06371 2838 4524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06370 4088 3263 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06369 5610 6376 5611 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06368 5611 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06367 5609 5992 5610 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06366 6212 6440 5609 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06365 5616 5749 5615 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06364 5615 5748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06363 5614 6893 5616 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06362 5750 6440 5614 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06361 6229 6235 6230 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06360 6082 6237 6229 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06359 6442 6229 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06358 vss 6229 6442 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06357 6085 6236 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06356 vss 6232 6236 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06355 6235 6237 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06354 vss 6984 6237 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06353 6083 6233 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06352 6230 6976 6083 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06351 6233 6237 6085 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06350 6084 6235 6233 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06349 vss 6230 6084 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06348 vss 6442 6081 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06347 6081 6976 6082 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06346 5130 5127 5131 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06345 5131 5132 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06344 5128 5343 5130 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06343 5141 5129 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06342 5129 5342 5128 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06341 3366 3449 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06340 4233 3455 3366 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06339 3365 3863 4233 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06338 vss 4071 3365 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06337 3365 3458 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06336 vss 2897 2899 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06335 2899 2896 2898 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06334 2895 2898 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06333 1575 1578 1457 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06332 1457 1757 1575 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06331 vss 4241 1457 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06330 4165 4166 4855 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06329 vss 4163 4165 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06328 4167 4649 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06327 4855 4164 4167 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06326 vss 4649 4166 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06325 4164 4163 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06324 vss 1505 704 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06323 704 1652 775 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06322 774 775 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06321 vss 3201 3093 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06320 3093 3591 3196 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06319 3195 3196 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06318 vss 2086 1650 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06317 1650 1649 1651 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06316 5949 1651 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06315 5945 6791 5946 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06314 5944 5943 5945 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06313 5946 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06312 5942 5945 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06311 vss 6637 5944 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06310 5944 6619 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06309 5418 5425 5417 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06308 vss 6665 5418 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06307 5419 5421 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06306 vss 5419 5420 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06305 5417 5424 5419 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06304 6665 5417 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06303 vss 5417 6665 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06302 5420 5424 5421 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06301 5421 5425 5422 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06300 vss 6580 5425 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06299 5424 5425 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06298 vss 5857 5423 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06297 5422 5423 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06296 6894 6904 6895 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06295 vss 6893 6894 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06294 6896 6898 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06293 vss 6896 6897 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06292 6895 6901 6896 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06291 6893 6895 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06290 vss 6895 6893 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06289 6897 6901 6898 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06288 6898 6904 6899 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06287 vss 6984 6904 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06286 6901 6904 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06285 vss 6900 6902 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06284 6899 6902 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06283 6688 6934 6543 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06282 vss 6694 6689 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06281 6543 6689 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06280 6144 6190 5930 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06279 5930 6191 6144 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06278 vss 5965 5930 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06277 1623 1624 6119 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06276 vss 6807 1623 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06275 1625 6590 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06274 6119 1622 1625 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06273 vss 6590 1624 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06272 1622 6807 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06271 594 1655 595 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06270 593 603 594 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06269 595 596 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06268 591 594 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06267 vss 592 593 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06266 593 607 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06265 vss 5069 2694 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06264 2694 2830 2831 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06263 3649 2831 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06262 4315 4413 4405 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06261 vss 4918 4315 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06260 4406 4409 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06259 vss 4406 4316 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06258 4405 4412 4406 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06257 4918 4405 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06256 vss 4405 4918 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06255 4316 4412 4409 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06254 4409 4413 4317 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06253 vss 6580 4413 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06252 4412 4413 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06251 vss 4410 4411 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06250 4317 4411 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06249 vss 482 318 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_06248 318 478 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_06247 766 317 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06246 318 477 317 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_06245 317 480 318 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_06244 1323 4176 1324 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06243 1324 1322 1323 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06242 vss 2747 1324 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06241 vss 5346 5228 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06240 5228 5559 5347 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06239 5345 5347 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06238 2218 2307 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06237 2304 2303 2218 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06236 2217 2479 2304 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06235 vss 2319 2217 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06234 2217 2483 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06233 5211 5749 5212 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06232 5212 5748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06231 5210 6885 5211 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06230 5315 5316 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06229 5316 6440 5210 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06228 6508 6615 6613 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06227 vss 6850 6508 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06226 6509 6839 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06225 6613 6612 6509 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06224 vss 6839 6615 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06223 6612 6850 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06222 4672 4673 4674 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06221 4674 4671 4672 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06220 vss 5965 4674 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06219 vss 6420 6423 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06218 6423 6421 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06217 vss 6422 6423 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06216 4349 4396 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06215 4395 4394 4349 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06214 612 614 611 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06213 vss 1513 612 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06212 613 619 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06211 611 610 613 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06210 vss 619 614 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06209 610 1513 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06208 2157 1194 450 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06207 450 1190 2157 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06206 vss 525 450 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06205 1683 1688 1684 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06204 1684 3593 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06203 1681 2347 1683 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06202 1682 1680 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06201 1680 1679 1681 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06200 3385 3328 3323 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06199 3321 3329 3385 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06198 3573 3385 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06197 vss 3385 3573 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06196 3325 3327 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06195 vss 3565 3327 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06194 3328 3329 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06193 vss 5054 3329 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06192 3322 3326 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06191 3323 6976 3322 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06190 3326 3329 3325 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06189 3324 3328 3326 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06188 vss 3323 3324 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06187 vss 3573 3320 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06186 3320 6976 3321 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06185 1671 1669 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06184 2045 1670 1671 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06183 vss 5735 5737 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06182 5737 5738 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06181 vss 5733 5737 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06180 4452 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06179 vss 6220 4452 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06178 4452 5300 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06177 vss 4572 4452 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06176 3947 4013 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06175 vss 3797 3947 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06174 3947 4217 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06173 vss 5502 3947 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06172 vss 502 366 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06171 366 830 365 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06170 vss 830 367 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06169 365 367 368 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06168 364 365 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06167 368 2048 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06166 vss 6903 6425 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06165 vss 6876 6425 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06164 6425 6877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06163 6424 6425 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06162 vss 4456 3217 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06161 3217 5987 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06160 vss 4477 3217 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06159 3468 6423 3467 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06158 3467 3947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06157 3715 3547 3468 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06156 vss 527 128 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06155 128 830 257 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06154 vss 830 259 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06153 257 259 129 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06152 258 257 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06151 129 2386 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06150 vss 829 720 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06149 720 830 832 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06148 vss 830 834 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06147 832 834 721 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06146 828 832 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06145 721 2793 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06144 vss 988 713 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06143 713 830 814 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06142 vss 830 815 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06141 814 815 714 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06140 810 814 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06139 714 2741 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06138 4339 5773 4340 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06137 4340 5889 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06136 4338 4501 4339 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06135 4502 6440 4338 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06134 vss 4083 3047 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06133 3047 4082 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06132 3046 3047 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06131 3633 3634 3520 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06130 3520 3632 3633 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06129 vss 3636 3520 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06128 3631 3633 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06127 3710 6423 3711 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06126 3711 3947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06125 3951 3709 3710 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06124 vss 636 102 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06123 102 1004 224 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06122 vss 1004 226 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06121 224 226 103 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06120 225 224 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06119 103 917 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06118 vss 825 447 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06117 447 1004 519 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06116 vss 1004 521 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06115 519 521 448 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06114 517 519 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06113 448 1196 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06112 vss 522 388 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06111 388 1004 389 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06110 vss 1004 391 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06109 389 391 390 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06108 387 389 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06107 390 1208 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06106 vss 4676 2681 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06105 2681 3046 2805 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06104 vss 3046 2806 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06103 2805 2806 2682 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06102 2801 2805 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06101 2682 2803 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06100 3825 4726 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06099 5115 5575 3825 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06098 3824 4053 5115 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06097 vss 5992 3824 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06096 3824 5773 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06095 5552 5999 5553 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06094 5553 6000 5552 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06093 vss 6440 5553 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06092 6552 6702 6553 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06091 6553 6701 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06090 6551 6704 6552 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06089 6948 6700 6551 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06088 vss 2553 1943 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06087 1943 2356 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06086 2154 1943 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06085 751 1649 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06084 965 2086 751 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06083 6550 6921 6549 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06082 6549 6917 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06081 6700 6963 6550 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06080 vss 4690 4887 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06079 4690 4688 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06078 4887 4689 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06077 vss 4682 4681 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06076 4681 4679 4680 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06075 4878 4680 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06074 3933 4086 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06073 4073 4281 3933 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06072 vss 4071 4073 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06071 4072 4073 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06070 vss 2361 2150 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06069 2150 4673 2359 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06068 vss 4673 2362 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06067 2359 2362 2153 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06066 2360 2359 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06065 2153 2551 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06064 6557 6704 6556 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06063 6556 6705 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06062 6966 6951 6557 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06061 1705 2544 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06060 1704 2142 1705 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06059 vss 1703 1704 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06058 427 488 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06057 592 779 427 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06056 426 489 592 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06055 vss 491 426 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06054 426 486 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06053 3204 3413 3097 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06052 3097 3414 3204 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06051 vss 5262 3097 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06050 3921 6221 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06049 vss 4261 3921 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06048 3921 4708 4456 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06047 4456 4071 3921 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06046 1102 1218 1103 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06045 1103 1732 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06044 1367 4748 1102 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06043 6844 6842 6845 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06042 6845 6843 6846 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06041 vss 6849 6844 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06040 6841 6846 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06039 5854 6591 5855 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06038 5855 6616 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06037 5853 6905 5854 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06036 5914 5917 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06035 5917 6807 5853 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06034 6132 5967 5928 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06033 5928 5993 6132 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06032 vss 5927 5928 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06031 5324 5947 5191 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06030 5191 5949 5324 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06029 vss 5964 5191 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06028 734 2194 735 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06027 735 857 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06026 733 1953 734 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06025 2787 3836 733 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06024 vss 1995 2406 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06023 1995 3460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06022 2406 2852 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06021 5985 5986 5988 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06020 5988 6214 5985 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06019 vss 6893 5988 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06018 2640 2722 2938 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06017 vss 2720 2640 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06016 2641 2919 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06015 2938 2719 2641 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06014 vss 2919 2722 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06013 2719 2720 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06012 5007 6791 5006 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06011 5005 5008 5007 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06010 5006 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06009 5003 5007 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06008 vss 6637 5005 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06007 5005 5004 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06006 3801 4275 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06005 vss 3800 3801 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06004 3801 4708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06003 vss 6224 3801 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06002 4463 3801 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06001 vss 3204 3096 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06000 3096 3596 3203 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05999 3202 3203 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05998 3057 4509 3059 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05997 3059 3062 3058 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05996 vss 3060 3057 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05995 3632 3058 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05994 5872 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05993 6629 6431 5872 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05992 5871 5959 6629 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05991 vss 6182 5871 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05990 5871 6183 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05989 6923 6932 6926 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05988 6924 6933 6923 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05987 6934 6923 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05986 vss 6923 6934 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05985 6929 6931 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05984 vss 6930 6931 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05983 6932 6933 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05982 vss 6984 6933 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05981 6925 6928 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05980 6926 6976 6925 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05979 6928 6933 6929 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05978 6927 6932 6928 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05977 vss 6926 6927 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05976 vss 6934 6922 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05975 6922 6976 6924 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05974 6594 6585 6497 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05973 6497 6586 6594 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05972 vss 6867 6497 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05971 vss 2142 1809 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05970 1809 2544 1930 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05969 1929 1930 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05968 vss 4687 2659 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05967 2659 3740 2759 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05966 2758 2759 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05965 796 2124 759 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05964 758 2122 796 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05963 759 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05962 793 796 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05961 vss 794 758 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05960 758 801 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05959 vss 5773 3844 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05958 3844 4265 3845 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05957 4082 3845 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05956 vss 5144 4341 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05955 4341 4523 4516 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05954 4517 4516 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05953 1931 986 989 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05952 989 987 1931 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05951 vss 988 989 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05950 vss 3174 3085 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05949 3085 3182 3175 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05948 3570 3175 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05947 3561 5949 3479 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05946 3479 5947 3561 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05945 vss 3969 3479 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05944 2900 2908 2901 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05943 vss 3376 2900 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05942 2902 2903 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05941 vss 2902 2904 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05940 2901 2907 2902 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05939 3376 2901 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05938 vss 2901 3376 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05937 2904 2907 2903 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05936 2903 2908 2905 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05935 vss 3160 2908 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05934 2907 2908 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05933 vss 3152 2906 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05932 2905 2906 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05931 vss 3010 2244 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05930 2244 3006 2376 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05929 2375 2376 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05928 vss 6917 5110 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05927 5110 6919 5111 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05926 5113 5111 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05925 vss 3818 2191 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05924 2191 2615 2190 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05923 2195 2190 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05922 3789 4213 3791 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05921 3791 4212 3789 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05920 vss 4696 3791 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05919 2493 3741 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05918 2492 2739 2493 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05917 vss 2733 2492 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05916 1065 1501 1066 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05915 1066 1320 1157 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05914 vss 2314 1065 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05913 1156 1157 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05912 6311 6314 6585 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05911 vss 6310 6311 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05910 6313 6778 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05909 6585 6312 6313 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05908 vss 6778 6314 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05907 6312 6310 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05906 5903 5791 5628 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05905 5628 5792 5903 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05904 vss 6250 5628 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05903 1317 2755 1318 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05902 1318 3586 1317 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05901 vss 2111 1318 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05900 3201 3199 3095 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05899 3095 3618 3201 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05898 vss 5959 3095 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05897 634 1194 635 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05896 635 1190 634 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05895 vss 633 635 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05894 918 634 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05893 3444 3634 3443 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05892 3443 3632 3444 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05891 vss 3442 3443 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05890 4947 3444 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05889 2089 2303 2091 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05888 2090 2479 2089 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05887 2091 2307 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05886 2088 2089 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05885 vss 2319 2090 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05884 2090 2483 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05883 3121 3260 3252 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05882 vss 3460 3121 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05881 3254 3257 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05880 vss 3254 3122 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05879 3252 3261 3254 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05878 3460 3252 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05877 vss 3252 3460 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05876 3122 3261 3257 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05875 3257 3260 3123 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05874 vss 3259 3260 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05873 3261 3260 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05872 vss 3459 3258 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05871 3123 3258 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05870 710 811 803 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05869 vss 988 710 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05868 804 806 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05867 vss 804 711 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05866 803 809 804 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05865 988 803 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05864 vss 803 988 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05863 711 809 806 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05862 806 811 712 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05861 vss 3160 811 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05860 809 811 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05859 vss 810 808 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05858 712 808 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05857 4606 5268 4607 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05856 4607 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05855 4605 5992 4606 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05854 4699 4698 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05853 4698 6440 4605 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05852 4507 4726 4266 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05851 4266 4265 4507 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05850 vss 5773 4266 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05849 3746 3753 3747 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05848 3744 3754 3746 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05847 3972 3746 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05846 vss 3746 3972 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05845 3751 3752 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05844 vss 3750 3752 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05843 3753 3754 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05842 vss 5054 3754 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05841 3745 3748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05840 3747 6976 3745 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05839 3748 3754 3751 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05838 3749 3753 3748 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05837 vss 3747 3749 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05836 vss 3972 3743 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05835 3743 6976 3744 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05834 370 376 369 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05833 vss 663 370 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05832 371 372 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05831 vss 371 373 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05830 369 377 371 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05829 663 369 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05828 vss 369 663 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05827 373 377 372 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05826 372 376 375 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05825 vss 3259 376 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05824 377 376 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05823 vss 661 374 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05822 375 374 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05821 970 2498 969 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05820 969 1649 970 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05819 vss 1172 969 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05818 968 970 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05817 vss 6224 5112 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05816 5112 4708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05815 vss 4524 5112 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05814 2043 2299 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05813 2095 2492 2043 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05812 3948 5967 3724 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05811 3724 5993 3948 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05810 vss 3969 3724 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05809 3316 3717 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05808 3315 3561 3316 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05807 vss 4611 3621 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05806 3621 4066 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05805 vss 3618 3621 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05804 5443 6806 5441 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05803 5441 6910 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05802 5442 5670 5443 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05801 vss 1704 2344 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05800 2344 1700 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05799 vss 1699 2344 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05798 2614 2615 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05797 2834 3818 2614 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05796 2494 3741 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05795 2511 2739 2494 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05794 6939 6945 6940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05793 6936 6947 6939 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05792 6963 6939 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05791 vss 6939 6963 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05790 6943 6944 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05789 vss 6946 6944 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05788 6945 6947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05787 vss 6984 6947 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05786 6938 6942 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05785 6940 6976 6938 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05784 6942 6947 6943 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05783 6941 6945 6942 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05782 vss 6940 6941 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05781 vss 6963 6937 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05780 6937 6976 6936 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05779 5252 6876 5174 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05778 5174 6877 5252 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05777 vss 5524 5174 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05776 5254 5252 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05775 3916 4051 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05774 4052 4613 3916 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05773 3372 3658 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05772 3371 4286 3372 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05771 2649 3186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05770 2739 5804 2649 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05769 3039 4737 3038 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05768 3038 3042 3039 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05767 vss 3044 3038 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05766 vss 5026 4650 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05765 4650 5014 4651 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05764 4649 4651 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05763 5225 5337 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05762 5340 5338 5225 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05761 vss 5336 5340 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05760 6232 5340 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05759 1086 1925 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05758 1196 1694 1086 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05757 3585 3737 3488 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05756 3488 3738 3585 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05755 vss 4308 3488 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05754 3586 3585 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05753 1424 1679 1423 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05752 1423 1687 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05751 1914 1911 1424 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05750 950 1169 949 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05749 949 2728 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05748 1151 1727 950 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05747 1363 5069 1364 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05746 1364 2830 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05745 4051 6440 1363 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05744 1451 5069 1450 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05743 1450 2830 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05742 1449 2799 1451 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05741 1559 6440 1449 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05740 2306 3740 2101 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05739 2101 2512 2306 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05738 vss 2314 2101 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05737 1627 1888 1626 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05736 1626 2304 1627 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05735 vss 1884 1626 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05734 5939 6423 5940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05733 5940 6374 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05732 5938 6375 5939 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05731 5937 5936 5938 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05730 3472 3553 3473 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05729 3473 3757 3554 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05728 vss 3953 3472 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05727 3552 3554 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05726 6366 6363 6365 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05725 6365 6364 6367 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05724 vss 6632 6366 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05723 6362 6367 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05722 4817 4946 4818 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05721 4818 4948 4949 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05720 vss 4947 4817 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05719 4945 4949 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05718 2529 5725 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05717 2530 3186 2529 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05716 vss 2758 2530 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05715 vss 2044 1912 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05714 vss 2045 1912 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05713 1912 2046 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05712 5721 1912 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05711 3197 3199 3094 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05710 3094 3618 3197 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05709 vss 5958 3094 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05708 vss 4509 1831 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05707 1831 1986 1984 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05706 1985 1984 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05705 vss 868 2352 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05704 868 4748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05703 2352 4524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05702 4152 4150 4155 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05701 4155 4153 4154 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05700 vss 6118 4152 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05699 4151 4154 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05698 1374 2506 1375 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05697 1375 1372 1373 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05696 vss 1985 1374 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05695 3042 1373 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05694 5015 5524 5016 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05693 5016 5914 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05692 5013 5670 5015 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05691 5014 5012 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05690 5012 6665 5013 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05689 3117 3849 3118 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05688 3118 3866 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05687 4068 3664 3117 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05686 vss 6919 5980 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05685 5980 6434 5979 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05684 6186 5979 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05683 vss 4441 2660 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05682 2660 3740 2760 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05681 2952 2760 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05680 160 219 489 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05679 vss 784 160 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05678 161 488 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05677 489 218 161 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05676 vss 488 219 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05675 218 784 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05674 vss 1177 1080 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05673 1080 1332 1179 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05672 1178 1179 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05671 6483 6490 6484 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05670 6482 6492 6483 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05669 6480 6483 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05668 vss 6483 6480 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05667 6488 6489 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05666 vss 6726 6489 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05665 6490 6492 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05664 vss 6984 6492 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05663 6485 6487 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05662 6484 6976 6485 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05661 6487 6492 6488 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05660 6486 6490 6487 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05659 vss 6484 6486 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05658 vss 6480 6481 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05657 6481 6976 6482 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05656 3445 3364 3358 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05655 3355 3363 3445 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05654 4239 3445 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05653 vss 3445 4239 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05652 3361 3362 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05651 vss 3640 3362 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05650 3364 3363 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05649 vss 6984 3363 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05648 3357 3360 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05647 3358 6976 3357 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05646 3360 3363 3361 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05645 3359 3364 3360 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05644 vss 3358 3359 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05643 vss 4239 3356 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05642 3356 6976 3355 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05641 vss 3589 3490 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05640 3490 3776 3590 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05639 3591 3590 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05638 vss 2507 2510 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05637 2510 2508 2509 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05636 3566 2509 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05635 1767 2125 1768 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05634 1768 1991 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05633 1765 4094 1767 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05632 2180 1766 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05631 1766 5363 1765 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05630 vss 2987 2989 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05629 2989 3610 2988 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05628 2986 2988 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05627 2097 3167 2098 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05626 2098 2495 2097 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05625 vss 2111 2098 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05624 6493 6582 6573 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05623 vss 6905 6493 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05622 6574 6575 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05621 vss 6574 6495 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05620 6573 6578 6574 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05619 6905 6573 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05618 vss 6573 6905 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05617 6495 6578 6575 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05616 6575 6582 6494 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05615 vss 6580 6582 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05614 6578 6582 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05613 vss 6589 6579 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05612 6494 6579 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05611 6093 6705 6094 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05610 6094 6690 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05609 6092 6951 6093 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05608 6959 6241 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05607 6241 6703 6092 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05606 599 1513 601 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05605 601 640 600 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05604 vss 2314 599 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05603 598 600 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05602 6907 6918 6908 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05601 vss 6906 6907 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05600 6909 6912 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05599 vss 6909 6911 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05598 6908 6916 6909 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05597 6906 6908 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05596 vss 6908 6906 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05595 6911 6916 6912 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05594 6912 6918 6913 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05593 vss 6984 6918 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05592 6916 6918 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05591 vss 6914 6915 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05590 6913 6915 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05589 6316 6318 6792 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05588 vss 6581 6316 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05587 6317 6590 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05586 6792 6315 6317 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05585 vss 6590 6318 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05584 6315 6581 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05583 6475 6714 6474 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05582 6474 6473 6475 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05581 vss 6471 6474 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05580 vss 3849 2275 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05579 2275 4088 2416 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05578 2415 2416 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05577 1689 1688 1690 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05576 1690 3593 1691 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05575 vss 2347 1689 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05574 1687 1691 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05573 4312 4393 4386 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05572 vss 5026 4312 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05571 4387 4390 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05570 vss 4387 4314 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05569 4386 4392 4387 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05568 5026 4386 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05567 vss 4386 5026 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05566 4314 4392 4390 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05565 4390 4393 4313 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05564 vss 6580 4393 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05563 4392 4393 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05562 vss 4395 4391 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05561 4313 4391 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05560 1088 1206 1198 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05559 vss 3790 1088 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05558 1199 1200 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05557 vss 1199 1090 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05556 1198 1204 1199 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05555 3790 1198 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05554 vss 1198 3790 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05553 1090 1204 1200 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05552 1200 1206 1089 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05551 vss 3259 1206 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05550 1204 1206 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05549 vss 1203 1205 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05548 1089 1205 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05547 5681 5723 5177 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05546 5177 5721 5681 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05545 vss 5927 5177 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05544 6837 6840 6847 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05543 vss 6835 6837 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05542 6838 6839 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05541 6847 6836 6838 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05540 vss 6839 6840 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05539 6836 6835 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05538 vss 5063 5490 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05537 5063 5065 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05536 5490 5062 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05535 5178 5258 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05534 5431 5444 5178 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05533 5184 5264 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05532 5263 5262 5184 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05531 584 586 587 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05530 585 2086 584 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05529 587 946 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05528 1312 584 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05527 vss 588 585 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05526 585 774 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05525 5518 5986 5517 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05524 5517 6214 5518 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05523 vss 6874 5517 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05522 4614 4616 4617 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05521 4617 6951 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05520 4615 4613 4614 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05519 4722 4717 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05518 4717 5772 4615 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05517 vss 6715 6472 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_05516 6472 6962 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_05515 6704 6470 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05514 6472 6713 6470 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_05513 6470 6469 6472 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_05512 323 319 321 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05511 321 320 323 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05510 vss 328 321 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05509 3497 5737 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05508 3606 3608 3497 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05507 3135 5116 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05506 3618 3218 3135 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05505 2213 2292 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05504 vss 2304 2213 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05503 2213 2291 2723 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05502 2723 2498 2213 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05501 6398 6172 6054 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05500 6054 6173 6398 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05499 vss 6188 6054 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05498 vss 1002 1003 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05497 1003 1004 1006 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05496 vss 1004 1008 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05495 1006 1008 1005 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05494 1001 1006 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05493 1005 2793 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05492 vss 1191 991 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05491 991 1004 992 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05490 vss 1004 994 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05489 992 994 995 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05488 990 992 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05487 995 2741 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05486 vss 1182 351 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05485 351 1004 353 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05484 vss 1004 352 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05483 353 352 354 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05482 350 353 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05481 354 2048 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05480 vss 633 98 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05479 98 1004 221 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05478 vss 1004 223 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05477 221 223 100 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05476 222 221 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05475 100 914 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05474 4219 4453 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05473 5965 4472 4219 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05472 3503 5116 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05471 5948 3617 3503 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05470 4588 4862 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05469 4665 4587 4588 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05468 3528 4089 3527 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05467 3527 4942 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05466 3526 3866 3528 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05465 4273 3836 3526 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05464 913 2161 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05463 2086 1900 913 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05462 3877 6423 3876 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05461 3876 3947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05460 4153 3946 3877 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05459 vss 3403 3400 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05458 3400 3976 3399 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05457 vss 3976 3402 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05456 3399 3402 3398 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05455 3397 3399 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05454 3398 3401 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05453 vss 3190 2661 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05452 2661 3976 2762 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05451 vss 3976 2765 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05450 2762 2765 2662 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05449 2961 2762 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05448 2662 2763 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05447 vss 2979 2980 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05446 2980 3976 2983 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05445 vss 3976 2984 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05444 2983 2984 2982 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05443 2977 2983 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05442 2982 2981 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05441 vss 525 125 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05440 125 1004 253 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05439 vss 1004 256 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05438 253 256 127 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05437 255 253 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05436 127 2386 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05435 6564 6952 6563 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05434 6563 6714 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05433 6562 6974 6564 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05432 6713 6963 6562 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05431 423 482 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05430 vss 478 423 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05429 423 477 961 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05428 961 480 423 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05427 2211 2289 2291 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05426 vss 2298 2211 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05425 2212 2308 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05424 2291 2288 2212 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05423 vss 2308 2289 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05422 2288 2298 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05421 947 1289 948 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05420 948 1158 947 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05419 vss 946 948 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05418 4216 4220 4218 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05417 4218 6600 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05416 4217 4485 4216 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05415 5179 5263 5180 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05414 5180 5259 5260 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05413 vss 5261 5179 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05412 5258 5260 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05411 vss 845 732 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05410 732 2394 848 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05409 vss 2394 850 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05408 848 850 731 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05407 1563 848 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05406 731 849 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05405 vss 4935 2175 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05404 2175 4094 2393 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05403 vss 4094 2395 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05402 2393 2395 2178 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05401 2394 2393 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05400 2178 4241 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05399 5893 6442 5891 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05398 vss 6714 5892 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05397 5891 5892 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05396 6554 6974 6555 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05395 6555 6917 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05394 6703 6963 6554 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05393 849 4524 455 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05392 vss 4748 538 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05391 455 538 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05390 3109 3818 3108 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05389 3108 5069 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05388 3107 5773 3109 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05387 3226 6440 3107 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05386 3102 5069 3101 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05385 3101 5068 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05384 3100 5992 3102 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05383 4220 6440 3100 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05382 vss 3391 1665 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05381 1665 2326 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05380 1667 1665 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05379 1793 1875 1794 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05378 1794 1877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05377 1792 2727 1793 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05376 2717 1876 1792 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05375 2916 2920 6172 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05374 vss 2915 2916 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05373 2918 2919 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05372 6172 2917 2918 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05371 vss 2919 2920 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05370 2917 2915 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05369 5035 5041 5037 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05368 5037 5036 5038 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05367 vss 5942 5035 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05366 5034 5038 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05365 4844 6791 4760 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05364 4759 5017 4844 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05363 4760 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05362 4843 4844 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05361 vss 6637 4759 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05360 4759 5250 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05359 3810 4489 3811 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05358 3811 4042 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05357 3809 3813 3810 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05356 4453 3808 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05355 3808 4051 3809 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05354 70 68 1649 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05353 vss 69 70 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05352 72 86 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05351 1649 71 72 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05350 vss 86 68 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05349 71 69 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05348 vss 1484 1281 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05347 1281 1287 1282 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05346 1478 1282 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05345 2768 2773 2664 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05344 2663 5953 2768 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05343 2664 4441 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05342 2766 2768 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05341 vss 3199 2663 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05340 2663 3618 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05339 vss 791 709 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05338 709 793 792 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05337 973 792 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05336 vss 2314 1069 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05335 1069 1320 1160 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05334 1298 1160 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05333 5173 5251 5250 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05332 vss 5524 5173 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05331 5172 6116 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05330 5250 5248 5172 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05329 vss 6116 5251 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05328 5248 5524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05327 vss 3460 1770 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05326 1770 3263 1769 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05325 2400 1769 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05324 vss 4485 4222 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05323 4222 4220 4221 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05322 4472 4221 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05321 1476 4524 1477 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05320 1477 4094 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05319 1475 4299 1476 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05318 2412 1590 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05317 1590 5363 1475 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05316 5708 4880 4775 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05315 4775 4881 5708 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05314 vss 5948 4775 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05313 1057 1145 1138 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05312 vss 3382 1057 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05311 1139 1142 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05310 vss 1139 1059 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05309 1138 1143 1139 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05308 3382 1138 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05307 vss 1138 3382 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05306 1059 1143 1142 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05305 1142 1145 1058 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05304 vss 3160 1145 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05303 1143 1145 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05302 vss 3315 1144 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05301 1058 1144 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05300 617 1904 618 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05299 616 3188 617 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05298 618 3217 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05297 615 617 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05296 vss 2746 616 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05295 616 1322 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05294 1669 1527 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05293 vss 1521 1669 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05292 vss 4941 3512 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05291 3512 4942 3628 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05290 4053 3628 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05289 1871 4501 1872 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05288 1872 4088 1983 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05287 vss 3460 1871 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05286 1982 1983 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05285 2477 2727 2476 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05284 2476 2728 2480 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05283 vss 2723 2477 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05282 2720 2480 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05281 668 676 669 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05280 vss 829 668 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05279 670 673 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05278 vss 670 672 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05277 669 675 670 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05276 829 669 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05275 vss 669 829 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05274 672 675 673 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05273 673 676 671 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05272 vss 3259 676 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05271 675 676 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05270 vss 828 674 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05269 671 674 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05268 6374 5502 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05267 vss 5954 6374 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05266 4487 4485 4335 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05265 4335 4737 4487 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05264 vss 4488 4335 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05263 5342 4487 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05262 2668 3226 2669 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05261 2669 2788 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05260 2667 4220 2668 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05259 2782 2783 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05258 2783 4485 2667 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05257 6074 6974 6073 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05256 6073 6917 6215 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05255 vss 6963 6074 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05254 6214 6215 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05253 1379 1580 1378 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05252 1378 1749 1379 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05251 vss 4748 1378 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05250 6859 6860 6858 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05249 vss 6874 6859 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05248 6857 6870 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05247 6858 6856 6857 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05246 vss 6870 6860 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05245 6856 6874 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05244 vss 5993 2779 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05243 2779 2775 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05242 vss 5967 2779 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05241 vss 3601 3602 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05240 3601 3783 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05239 3602 3600 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05238 2942 3737 2943 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05237 2943 3738 2942 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05236 vss 5272 2943 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05235 2950 2942 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05234 5104 5721 4780 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05233 4780 5723 5104 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05232 vss 5964 4780 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05231 3319 3549 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05230 3318 3317 3319 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05229 36 111 107 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05228 vss 504 36 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05227 37 39 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05226 vss 37 38 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05225 107 40 37 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05224 504 107 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05223 vss 107 504 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05222 38 40 39 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05221 39 111 110 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05220 vss 3259 111 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05219 40 111 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05218 vss 239 112 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05217 110 112 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05216 vss 6725 6730 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05215 6730 6728 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05214 6726 6730 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05213 2785 4220 2671 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05212 2670 2998 2785 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05211 2671 5116 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05210 4483 2785 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05209 vss 2999 2670 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05208 2670 2997 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05207 750 1313 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05206 1300 961 750 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05205 5532 5533 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05204 6491 5531 5532 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05203 3469 3714 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05202 3548 3558 3469 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05201 401 863 400 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05200 400 402 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05199 399 6440 401 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05198 1818 2155 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05197 1950 2135 1818 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05196 1817 1947 1950 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05195 vss 2057 1817 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05194 1816 2360 1950 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05193 vss 1946 1816 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05192 5926 6806 5924 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05191 5924 6910 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05190 5925 6665 5926 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05189 5665 5792 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05188 5788 5789 5665 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05187 vss 6966 6969 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05186 6969 6968 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05185 6967 6969 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05184 6559 6705 6558 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05183 6558 6707 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05182 6970 6951 6559 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05181 6920 6919 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05180 6951 6917 6920 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05179 vss 5497 5498 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05178 5497 5508 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05177 5498 5730 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05176 vss 4445 4679 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05175 4445 4444 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05174 4679 4447 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05173 6048 6423 6049 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05172 6049 6374 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05171 6047 6375 6048 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05170 6363 6165 6047 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05169 2234 2344 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05168 2346 2345 2234 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05167 3428 5749 3427 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05166 3427 5748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05165 3617 6440 3428 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05164 4370 5341 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05163 4616 5992 4370 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05162 1554 1580 1442 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05161 1442 1749 1554 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05160 vss 4275 1442 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05159 2521 1554 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05158 2232 3186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05157 2333 6187 2232 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05156 1815 1945 1814 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05155 1814 2139 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05154 1947 2138 1815 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05153 6634 6791 6524 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05152 6523 6855 6634 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05151 6524 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05150 6632 6634 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05149 vss 6637 6523 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05148 6523 6858 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05147 vss 4489 4336 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05146 4336 4496 4490 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05145 4488 4490 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05144 2996 3792 2995 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05143 2995 3793 2996 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05142 vss 3423 2995 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05141 434 641 435 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05140 435 3195 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05139 433 629 434 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05138 494 3217 433 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05137 1743 4937 1742 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05136 1742 2352 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05135 1744 4094 1743 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05134 1376 1576 1377 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05133 1377 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05132 1562 4094 1376 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05131 2172 2392 2171 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05130 2171 2170 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05129 2173 2389 2172 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05128 726 3813 727 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05127 727 844 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05126 725 851 726 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05125 1194 3226 725 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05124 912 1171 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05123 911 1727 912 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05122 2642 2725 3174 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05121 vss 2723 2642 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05120 2643 2924 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05119 3174 2724 2643 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05118 vss 2924 2725 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05117 2724 2723 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05116 vss 4883 4776 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05115 4776 4886 4884 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05114 5702 4884 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05113 5042 6423 5043 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05112 5043 6374 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05111 5040 6375 5042 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05110 5041 5039 5040 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05109 4359 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05108 4444 6431 4359 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05107 4358 4441 4444 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05106 vss 6220 4358 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05105 4358 5300 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05104 6051 6360 6050 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05103 6050 6167 6168 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05102 vss 6371 6051 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05101 6166 6168 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05100 4767 4866 4766 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05099 4766 5029 4864 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05098 vss 4863 4767 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05097 4862 4864 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05096 3652 3453 3454 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05095 3454 3451 3652 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05094 vss 3452 3454 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05093 2159 2165 2160 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05092 2160 3004 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05091 2158 2562 2159 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05090 2520 2157 2158 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05089 5196 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05088 5279 6431 5196 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05087 5195 6187 5279 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05086 vss 5954 5195 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05085 5195 5502 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05084 vss 1518 1425 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05083 1425 1517 1519 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05082 3401 1519 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05081 vss 975 977 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05080 977 980 976 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05079 1328 976 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05078 314 335 311 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05077 311 310 314 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05076 vss 607 311 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05075 4225 4275 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05074 vss 4224 4225 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05073 4225 4708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05072 vss 6224 4225 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05071 4929 4225 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05070 vss 1917 2046 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05069 1917 2521 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05068 2046 2535 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05067 5664 6917 5663 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05066 5663 6448 5785 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05065 vss 6682 5664 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05064 6014 5785 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05063 vss 1169 410 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05062 410 581 460 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05061 569 460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05060 vss 1914 1808 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05059 1808 1913 1915 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05058 2044 1915 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05057 vss 2387 135 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05056 135 133 134 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05055 987 134 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05054 1894 3167 1801 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05053 1801 2495 1894 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05052 vss 2111 1801 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05051 1893 1894 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05050 vss 947 699 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05049 699 941 764 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05048 770 764 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05047 vss 2895 2210 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05046 2210 2286 2287 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05045 2716 2287 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05044 1855 2154 1856 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05043 1856 1945 1941 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05042 vss 2122 1855 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05041 2050 1941 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05040 vss 2949 2951 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05039 2949 2953 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05038 2951 2950 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05037 336 784 338 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05036 338 494 337 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05035 vss 2314 336 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05034 335 337 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05033 vss 974 1172 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05032 974 1178 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05031 1172 973 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05030 vss 1900 1802 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05029 1802 2161 1896 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05028 2106 1896 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05027 vss 1758 1738 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05026 1738 1967 1739 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05025 1737 1739 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05024 2094 2095 2096 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05023 2093 2485 2094 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05022 2096 2102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05021 2092 2094 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05020 vss 2319 2093 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05019 2093 2320 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05018 3317 5723 3083 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05017 3083 5721 3317 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05016 vss 3969 3083 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05015 6782 6790 6781 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05014 vss 6807 6782 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05013 6783 6784 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05012 vss 6783 6785 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05011 6781 6789 6783 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05010 6807 6781 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05009 vss 6781 6807 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05008 6785 6789 6784 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05007 6784 6790 6788 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05006 vss 6832 6790 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05005 6789 6790 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05004 vss 6786 6787 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05003 6788 6787 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05002 5600 5718 5709 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05001 vss 5953 5600 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05000 5711 5714 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04999 vss 5711 5601 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04998 5709 5717 5711 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04997 5953 5709 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04996 vss 5709 5953 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04995 5601 5717 5714 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04994 5714 5718 5602 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04993 vss 6832 5718 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04992 5717 5718 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04991 vss 5715 5716 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04990 5602 5716 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04989 5136 5749 5135 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04988 5135 5748 5137 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04987 vss 6440 5136 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04986 5133 5137 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04985 3134 4220 3133 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04984 3133 3226 3214 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04983 vss 4485 3134 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04982 3424 3214 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04981 5641 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04980 6167 6431 5641 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04979 5640 5725 6167 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04978 vss 6182 5640 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04977 5640 6183 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04976 854 863 741 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04975 741 1035 854 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04974 vss 1038 741 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04973 1004 854 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04972 644 651 643 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04971 vss 3796 644 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04970 645 646 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04969 vss 645 647 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04968 643 650 645 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04967 3796 643 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04966 vss 643 3796 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04965 647 650 646 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04964 646 651 649 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04963 vss 3160 651 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04962 650 651 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04961 vss 652 648 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04960 649 648 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04959 4714 5748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04958 4713 5545 4714 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04957 vss 4715 4713 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04956 6188 4713 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04955 2152 2553 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04954 vss 2534 2151 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04953 2998 2521 2152 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04952 2151 2520 2998 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04951 3406 3413 3405 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04950 3405 3414 3406 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04949 vss 5243 3405 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04948 3404 3406 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04947 3941 4088 3942 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04946 3942 4091 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04945 3940 4089 3941 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04944 5889 4090 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04943 4090 4087 3940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04942 3052 5773 3054 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04941 3054 4491 3053 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04940 vss 4524 3052 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04939 3051 3053 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04938 5636 5680 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04937 5682 5681 5636 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04936 1307 1311 4673 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04935 vss 1306 1307 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04934 1310 1309 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04933 4673 1308 1310 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04932 vss 1309 1311 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04931 1308 1306 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04930 5069 3456 2695 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04929 2695 3457 5069 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04928 vss 3455 2695 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04927 1411 1737 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04926 1632 2506 1411 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04925 1410 1882 1632 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04924 vss 1885 1410 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04923 1410 1891 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04922 5185 5264 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04921 5436 5372 5185 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04920 vss 3395 3086 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04919 3086 3976 3177 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04918 vss 3976 3180 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04917 3177 3180 3087 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04916 3337 3177 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04915 3087 3178 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04914 vss 6422 6210 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04913 vss 6421 6210 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04912 6210 6420 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04911 6211 6210 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04910 6795 6876 6796 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04909 6796 6877 6795 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04908 vss 6807 6796 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04907 6794 6795 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04906 195 1900 144 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04905 143 470 195 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04904 144 2161 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04903 302 195 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04902 vss 598 143 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04901 143 307 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04900 3616 3792 3504 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04899 3504 3793 3616 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04898 vss 3802 3504 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04897 3508 3816 3509 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04896 3509 5115 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04895 3969 3814 3508 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04894 vss 3759 3760 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04893 3760 3976 3764 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04892 vss 3976 3762 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04891 3764 3762 3763 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04890 3758 3764 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04889 3763 3761 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04888 vss 3972 3389 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04887 3389 3976 3568 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04886 vss 3976 3569 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04885 3568 3569 3390 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04884 3750 3568 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04883 3390 3570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04882 vss 3979 3891 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04881 3891 3976 3974 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04880 vss 3976 3977 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04879 3974 3977 3892 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04878 3986 3974 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04877 3892 3975 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04876 vss 3573 3387 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04875 3387 3976 3564 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04874 vss 3976 3567 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04873 3564 3567 3386 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04872 3565 3564 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04871 3386 3566 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04870 4173 4414 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04869 4410 4175 4173 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04868 602 1317 604 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04867 604 640 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04866 603 2314 602 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04865 4920 5805 4793 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04864 4793 5756 4920 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04863 vss 4918 4793 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04862 4919 4920 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04861 2059 3006 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04860 2058 3010 2059 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04859 4009 4213 3905 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04858 3905 4212 4009 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04857 vss 4897 3905 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04856 3756 6434 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04855 3757 6919 3756 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04854 3755 5243 3757 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04853 vss 4217 3755 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04852 3755 5502 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04851 5652 6226 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04850 6205 6426 5652 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04849 5651 5804 6205 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04848 vss 6182 5651 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04847 5651 6183 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04846 vss 3790 993 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04845 993 2797 1193 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04844 vss 2797 1195 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04843 1193 1195 996 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04842 1203 1193 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04841 996 1196 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04840 vss 3423 1009 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04839 1009 2797 1011 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04838 vss 2797 1012 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04837 1011 1012 1010 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04836 1007 1011 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04835 1010 1208 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04834 4860 6876 4765 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04833 4765 6877 4860 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04832 vss 4914 4765 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04831 4859 4860 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04830 vss 6850 6507 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04829 6507 6839 6611 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04828 6814 6611 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04827 421 1513 422 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04826 422 640 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04825 476 2314 421 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04824 639 2142 642 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04823 642 2544 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04822 640 3217 639 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04821 25 772 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04820 69 1151 25 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04819 3817 3816 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04818 4048 3814 3817 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04817 4288 4941 4289 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04816 4289 4287 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04815 4284 4286 4288 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04814 4285 4524 4284 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04813 2115 2740 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04812 2116 2520 2115 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04811 vss 2117 2116 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04810 6748 6191 5966 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04809 5966 6190 6748 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04808 vss 5964 5966 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04807 5974 6209 5976 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04806 5976 5975 5977 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04805 vss 5973 5974 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04804 5972 5977 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04803 729 2194 730 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04802 730 845 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04801 728 1953 729 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04800 1212 3836 728 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04799 2685 5069 2684 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04798 2684 2807 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04797 2683 5773 2685 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04796 4485 6440 2683 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04795 vss 2341 2342 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04794 2341 2349 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04793 2342 2535 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04792 2653 2940 2652 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04791 2652 2744 2743 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04790 vss 2938 2653 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04789 2742 2743 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04788 778 1300 705 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04787 705 776 778 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04786 vss 870 705 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04785 1163 778 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04784 vss 5157 2417 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04783 2417 4299 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04782 2418 2417 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04781 2082 2079 2919 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04780 vss 2895 2082 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04779 2083 2080 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04778 2919 2081 2083 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04777 vss 2080 2079 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04776 2081 2895 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04775 6531 6885 6530 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04774 6530 6874 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04773 6529 6893 6531 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04772 6839 6646 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04771 6646 6906 6529 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04770 vss 2534 1702 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04769 1702 2553 1701 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04768 1700 1701 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04767 1356 1580 1355 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04766 1355 1749 1356 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04765 vss 4275 1355 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04764 vss 2492 1800 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04763 1800 2299 1889 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04762 1888 1889 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04761 6026 6113 6115 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04760 vss 6112 6026 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04759 6027 6116 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04758 6115 6114 6027 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04757 vss 6116 6113 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04756 6114 6112 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04755 2658 5725 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04754 2756 3186 2658 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04753 vss 2758 2756 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04752 2755 2756 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04751 vss 2938 2939 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04750 2939 2940 2941 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04749 3975 2941 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04748 vss 5560 5559 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04747 5560 5784 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04746 5559 5749 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04745 vss 3658 3516 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04744 3516 4942 3630 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04743 5068 3630 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04742 vss 2512 2233 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04741 2233 2349 2334 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04740 2519 2334 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04739 2635 2713 2705 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04738 vss 3546 2635 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04737 2707 2708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04736 vss 2707 2636 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04735 2705 2710 2707 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04734 3546 2705 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04733 vss 2705 3546 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04732 2636 2710 2708 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04731 2708 2713 2637 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04730 vss 3160 2713 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04729 2710 2713 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04728 vss 3318 2711 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04727 2637 2711 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04726 4262 5773 4263 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04725 4263 4265 4264 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04724 vss 6440 4262 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04723 4492 4264 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04722 3507 5068 3506 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04721 3506 4062 3623 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04720 vss 5069 3507 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04719 3798 3623 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04718 vss 4286 3529 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04717 3529 3658 3643 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04716 3818 3643 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04715 1413 2161 1412 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04714 1412 2498 1497 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04713 vss 1900 1413 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04712 1640 1497 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04711 1389 2409 1391 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04710 1391 2198 1389 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04709 vss 1587 1391 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04708 5993 2106 2108 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04707 2108 2107 5993 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04706 vss 2109 2108 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04705 5647 5936 5646 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04704 5646 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04703 5645 5992 5647 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04702 5735 5732 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04701 5732 6440 5645 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04700 1415 2736 1500 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04699 1500 2498 1416 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04698 1416 2106 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04697 1414 2535 1500 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04696 vss 3217 1414 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04695 vss 2111 1415 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04694 1498 1500 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04693 51 131 126 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04692 vss 527 51 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04691 52 54 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04690 vss 52 53 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04689 126 55 52 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04688 527 126 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04687 vss 126 527 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04686 53 55 54 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04685 54 131 130 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04684 vss 3259 131 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04683 55 131 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04682 vss 258 132 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04681 130 132 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04680 5727 5954 5494 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04679 5494 5502 5727 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04678 vss 5804 5494 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04677 5320 5986 5214 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04676 5214 6214 5320 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04675 vss 6885 5214 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04674 1866 3866 1867 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04673 1867 2352 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04672 1865 3849 1866 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04671 2399 1980 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04670 1980 3664 1865 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04669 3225 5987 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04668 vss 3221 3225 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04667 3225 4456 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04666 vss 4477 3225 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04665 3045 6727 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04664 3044 3046 3045 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04663 3043 3042 3044 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04662 vss 3245 3043 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04661 3041 3248 3044 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04660 vss 4748 3041 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04659 162 235 228 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04658 vss 500 162 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04657 229 231 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04656 vss 229 164 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04655 228 233 229 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04654 500 228 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04653 vss 228 500 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04652 164 233 231 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04651 231 235 163 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04650 vss 3160 235 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04649 233 235 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04648 vss 237 234 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04647 163 234 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04646 6806 6420 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04645 vss 6222 6806 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04644 6806 6422 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04643 vss 6186 6806 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04642 6930 6935 6548 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04641 6548 6696 6930 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04640 vss 6706 6548 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04639 3781 4213 3782 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04638 3782 4212 3781 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04637 vss 4438 3782 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04636 4682 5954 4683 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04635 4683 5502 4682 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04634 vss 5953 4683 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04633 3713 3950 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04632 3712 3725 3713 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04631 6203 6190 6062 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04630 6062 6191 6203 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04629 vss 6188 6062 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04628 2821 3040 2692 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04627 2692 2820 2821 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04626 vss 3238 2692 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04625 2824 2821 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04624 5444 5949 5445 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04623 5445 5947 5444 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04622 vss 5927 5445 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04621 6096 6917 6095 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04620 6095 6448 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04619 6705 6480 6096 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04618 5097 5986 5098 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04617 5098 6214 5097 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04616 vss 6740 5098 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04615 3793 1989 1452 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04614 1452 1745 3793 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04613 vss 1560 1452 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04612 2987 3413 2985 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04611 2985 3414 2987 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04610 vss 6265 2985 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04609 1619 2897 1621 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04608 1621 2896 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04607 1620 2921 1619 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04606 3878 4151 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04605 3949 3948 3878 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04604 vss 5727 5608 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04603 5608 5728 5729 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04602 6170 5729 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04601 6797 6806 6799 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04600 6799 6910 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04599 6798 6905 6797 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04598 6810 6806 6809 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04597 6809 6910 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04596 6808 6807 6810 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04595 5572 5907 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04594 5791 6440 5572 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04593 6451 6448 6450 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04592 6450 6449 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04591 6701 6917 6451 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04590 6445 6917 6446 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04589 6446 6448 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04588 6702 6682 6445 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04587 416 591 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04586 586 589 416 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04585 4246 5341 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04584 4613 5575 4246 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04583 1075 1209 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04582 1171 1876 1075 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04581 1796 2088 1795 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04580 1795 1882 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04579 1883 2095 1796 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04578 vss 2400 1828 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04577 1828 1975 1976 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04576 3221 1976 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04575 4354 4865 4355 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04574 4355 4675 4415 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04573 vss 4668 4354 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04572 4414 4415 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04571 1508 2946 1419 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04570 1419 2950 1508 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04569 vss 2111 1419 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04568 2923 2925 6190 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04567 vss 2921 2923 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04566 2926 2924 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04565 6190 2922 2926 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04564 vss 2924 2925 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04563 2922 2921 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04562 5868 5953 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04561 5867 5954 5868 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04560 5866 6867 5867 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04559 vss 5951 5866 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04558 5866 5952 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04557 6319 6591 6321 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04556 6321 6616 6320 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04555 vss 6807 6319 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04554 6778 6320 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04553 202 1900 147 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04552 146 607 202 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04551 147 2161 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04550 200 202 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04549 vss 335 146 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04548 146 310 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04547 3029 3036 3030 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04546 3026 3035 3029 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04545 4937 3029 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04544 vss 3029 4937 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04543 3033 3034 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04542 vss 3039 3034 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04541 3036 3035 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04540 vss 3259 3035 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04539 3028 3032 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04538 3030 6976 3028 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04537 3032 3035 3033 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04536 3031 3036 3032 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04535 vss 3030 3031 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04534 vss 4937 3027 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04533 3027 6976 3026 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04532 4903 6220 4697 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04531 4697 5300 4903 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04530 vss 4696 4697 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04529 5915 6876 5916 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04528 5916 6877 5915 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04527 vss 6905 5916 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04526 1422 1517 1421 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04525 1421 1662 1516 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04524 vss 1518 1422 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04523 1695 1516 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04522 6002 6691 6001 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04521 6003 6440 6002 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04520 6001 6921 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04519 6182 6002 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04518 vss 5999 6003 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04517 6003 6000 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04516 3598 4213 3493 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04515 3493 4212 3598 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04514 vss 4205 3493 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04513 1807 2375 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04512 1905 1904 1807 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04511 vss 2382 1905 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04510 3768 3777 3769 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04509 vss 5963 3768 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04508 3770 3772 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04507 vss 3770 3771 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04506 3769 3774 3770 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04505 5963 3769 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04504 vss 3769 5963 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04503 3771 3774 3772 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04502 3772 3777 3773 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04501 vss 5054 3777 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04500 3774 3777 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04499 vss 4200 3775 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04498 3773 3775 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04497 3495 5737 3494 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04496 3494 3598 3599 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04495 vss 3608 3495 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04494 3596 3599 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04493 vss 1395 1387 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04492 1387 2400 1386 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04491 1385 1386 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04490 vss 5748 5547 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04489 5547 5545 5546 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04488 5544 5546 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04487 1870 2407 1869 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04486 1869 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04485 1868 4094 1870 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04484 1979 1981 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04483 1981 3664 1868 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04482 1839 2125 1838 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04481 1838 1991 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04480 1837 4094 1839 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04479 2207 5363 1837 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04478 1994 2629 1840 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04477 1840 2418 1994 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04476 vss 2208 1840 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04475 1992 1994 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04474 vss 2489 1799 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04473 1799 2299 1887 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04472 1885 1887 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04471 vss 1727 951 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04470 951 1171 952 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04469 2727 952 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04468 vss 5963 2497 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04467 2497 3186 2496 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04466 2495 2496 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04465 5125 2999 2559 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04464 2559 2997 5125 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04463 vss 2998 2559 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04462 4703 5753 4702 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04461 4702 5767 4703 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04460 vss 4914 4702 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04459 2548 2545 2549 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04458 2549 3602 2547 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04457 vss 2546 2548 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04456 2544 2547 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04455 2954 5953 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04454 2953 3186 2954 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04453 vss 2952 2953 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04452 vss 5575 5555 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04451 5555 5877 5554 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04450 5999 5554 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04449 2612 5157 2611 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04448 2611 3263 2613 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04447 vss 5363 2612 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04446 2807 2613 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04445 1782 2407 1783 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04444 1783 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04443 1781 4094 1782 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04442 2198 3664 1781 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04441 vss 5758 5620 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04440 5620 5766 5760 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04439 5759 5760 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04438 2109 2116 2110 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04437 2110 2514 2109 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04436 vss 2323 2110 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04435 1842 2727 1841 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04434 1841 1877 1878 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04433 vss 1876 1842 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04432 2080 1878 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04431 1036 6469 1037 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04430 1037 1039 1036 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04429 vss 1578 1037 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04428 1035 1036 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04427 3900 4001 3993 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04426 vss 5725 3900 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04425 3995 3997 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04424 vss 3995 3901 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04423 3993 4000 3995 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04422 5725 3993 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04421 vss 3993 5725 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04420 3901 4000 3997 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04419 3997 4001 3902 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04418 vss 5054 4001 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04417 4000 4001 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04416 vss 4002 3998 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04415 3902 3998 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04414 142 200 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04413 vss 322 142 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04412 142 191 576 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04411 576 2498 142 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04410 5203 5501 5204 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04409 5204 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04408 5202 5992 5203 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04407 5297 5298 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04406 5298 6440 5202 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04405 3090 5958 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04404 3188 3186 3090 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04403 vss 3187 3188 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04402 3009 5116 3008 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04401 3008 3227 3011 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04400 vss 3218 3009 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04399 3006 3011 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04398 3353 3831 3354 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04397 3354 3629 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04396 3352 4253 3353 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04395 3438 3437 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04394 3437 3827 3352 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04393 3392 3740 3394 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04392 3393 5372 3392 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04391 3394 4897 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04390 3391 3392 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04389 vss 3737 3393 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04388 3393 3738 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04387 444 516 509 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04386 vss 3607 444 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04385 510 513 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04384 vss 510 446 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04383 509 514 510 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04382 3607 509 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04381 vss 509 3607 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04380 446 514 513 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04379 513 516 445 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04378 vss 3259 516 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04377 514 516 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04376 vss 657 515 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04375 445 515 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04374 5319 5112 5114 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04373 5114 5113 5319 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04372 vss 5134 5114 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04371 4814 4941 4815 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04370 4815 4942 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04369 4813 5349 4814 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04368 5545 4943 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04367 4943 6440 4813 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04366 4287 4748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04365 vss 4094 4287 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04364 5858 5918 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04363 5857 5856 5858 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04362 5183 5264 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04361 5919 5902 5183 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04360 vss 6225 5566 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04359 5566 5567 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04358 5573 5566 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04357 1070 1161 2138 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04356 vss 1163 1070 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04355 1071 1309 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04354 2138 1162 1071 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04353 vss 1309 1161 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04352 1162 1163 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04351 4913 5805 4791 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04350 4791 5756 4913 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04349 vss 5026 4791 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04348 4911 4913 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04347 1673 2124 1674 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04346 1672 2122 1673 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04345 1674 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04344 1913 1673 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04343 vss 1682 1672 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04342 1672 1911 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04341 3368 3458 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04340 3453 3863 3368 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04339 3367 3455 3453 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04338 vss 3456 3367 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04337 3367 3457 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04336 4462 5112 4242 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04335 4242 5113 4462 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04334 vss 4241 4242 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04333 932 3263 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04332 1233 3460 932 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04331 1237 1588 1127 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04330 1127 1239 1237 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04329 vss 1576 1127 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04328 1236 1237 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04327 2550 3199 2552 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04326 2552 3618 2550 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04325 vss 5804 2552 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04324 vss 2749 2940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04323 2940 2750 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04322 vss 2752 2940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04321 vss 3421 2561 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04320 2561 2797 2564 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04319 vss 2797 2565 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04318 2564 2565 2563 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04317 2560 2564 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04316 2563 2741 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04315 vss 3604 1431 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04314 1431 2797 1539 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04313 vss 2797 1540 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04312 1539 1540 1432 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04311 1549 1539 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04310 1432 2048 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04309 vss 3607 658 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04308 658 2797 660 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04307 vss 2797 662 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04306 660 662 659 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04305 657 660 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04304 659 914 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04303 vss 3796 653 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04302 653 2797 654 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04301 vss 2797 656 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04300 654 656 655 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04299 652 654 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04298 655 917 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04297 5529 5528 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04296 5585 5978 5529 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04295 397 686 396 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04294 396 395 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04293 986 3021 397 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04292 vss 3434 678 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04291 678 2797 679 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04290 vss 2797 681 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04289 679 681 680 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04288 677 679 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04287 680 2386 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04286 vss 3802 2674 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04285 2674 2797 2794 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04284 vss 2797 2798 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04283 2794 2798 2675 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04282 2792 2794 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04281 2675 2793 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04280 vss 3660 3536 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04279 3536 3663 3661 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04278 3662 3661 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04277 6677 6876 6542 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04276 6542 6877 6677 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04275 vss 6893 6542 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04274 6676 6677 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04273 4481 4572 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04272 vss 4709 4481 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04271 4481 5548 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04270 vss 4477 4481 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04269 4612 4481 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04268 vss 3606 3213 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04267 3213 3212 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04266 3210 3213 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04265 3521 4726 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04264 3636 5575 3521 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04263 2205 4941 2204 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04262 2204 4089 2206 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04261 2206 2412 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04260 2203 2411 2204 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04259 vss 2615 2203 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04258 vss 2415 2205 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04257 2202 2204 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04256 2119 2520 2120 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04255 2120 2331 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04254 2329 2740 2119 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04253 vss 2336 2335 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04252 2335 2342 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04251 2750 2335 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04250 6059 6390 6058 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04249 6058 6184 6181 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04248 vss 6869 6059 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04247 6180 6181 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04246 vss 2583 2584 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04245 2584 2587 2586 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04244 vss 2587 2588 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04243 2586 2588 2585 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04242 2582 2586 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04241 2585 5125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04240 6033 6919 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04239 6129 6434 6033 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04238 6032 6867 6129 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04237 vss 6128 6032 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04236 6032 6127 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04235 2601 2823 2602 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04234 2602 2600 2601 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04233 vss 2817 2602 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04232 vss 500 108 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04231 108 830 236 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04230 vss 830 238 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04229 236 238 109 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04228 237 236 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04227 109 914 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04226 vss 504 113 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04225 113 830 240 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04224 vss 830 241 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04223 240 241 114 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04222 239 240 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04221 114 917 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04220 vss 663 664 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04219 664 830 666 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04218 vss 830 667 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04217 666 667 665 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04216 661 666 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04215 665 1196 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04214 vss 392 116 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04213 116 830 242 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04212 vss 830 244 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04211 242 244 117 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04210 243 242 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04209 117 1208 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04208 6252 6259 6253 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04207 6104 6260 6252 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04206 6263 6252 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04205 vss 6252 6263 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04204 6107 6257 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04203 vss 6256 6257 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04202 6259 6260 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04201 vss 6984 6260 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04200 6105 6254 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04199 6253 6976 6105 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04198 6254 6260 6107 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04197 6106 6259 6254 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04196 vss 6253 6106 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04195 vss 6263 6103 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04194 6103 6976 6104 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04193 4620 4732 4621 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04192 4621 4618 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04191 4619 5115 4620 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04190 4948 4736 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04189 4736 5552 4619 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04188 1110 1953 1111 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04187 1111 2194 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04186 1109 3836 1110 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04185 1572 6440 1109 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04184 vss 571 574 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04183 574 573 575 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04182 776 575 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04181 3938 4088 3939 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04180 3939 4091 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04179 3936 4089 3938 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04178 4086 4087 3936 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04177 3003 3413 3002 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04176 3002 3414 3003 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04175 vss 6727 3002 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04174 vss 4524 4232 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04173 vss 4708 4232 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04172 4232 6224 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04171 4470 4232 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04170 4211 5068 4210 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04169 4210 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04168 4209 5069 4211 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04167 4689 4208 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04166 4208 4308 4209 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04165 3538 3849 3539 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04164 3539 3866 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04163 3537 4524 3538 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04162 3663 3665 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04161 3665 3664 3537 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04160 4031 4275 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04159 vss 4028 4031 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04158 4031 4708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04157 vss 6224 4031 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04156 5321 4031 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04155 vss 1359 1553 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04154 1359 4524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04153 1553 4748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04152 vss 4501 2187 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04151 2187 3229 2189 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04150 2188 2189 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04149 4770 4877 4868 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04148 vss 5039 4770 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04147 4869 4872 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04146 vss 4869 4771 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04145 4868 4875 4869 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04144 5039 4868 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04143 vss 4868 5039 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04142 4771 4875 4872 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04141 4872 4877 4772 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04140 vss 5054 4877 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04139 4875 4877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04138 vss 4873 4874 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04137 4772 4874 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04136 1446 1968 1445 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04135 1445 1558 1557 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04134 vss 1559 1446 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04133 1724 1557 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04132 2149 2356 2148 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04131 2148 2553 2147 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04130 vss 2331 2149 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04129 2146 2147 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04128 3779 4909 3778 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04127 3778 3781 3780 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04126 vss 3788 3779 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04125 3776 3780 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04124 vss 2506 622 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04123 622 1737 623 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04122 2498 623 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04121 4238 5112 4237 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04120 4237 5113 4238 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04119 vss 4235 4237 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04118 vss 3234 3113 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04117 3113 3233 3235 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04116 3231 3235 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04115 1382 3849 1383 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04114 1383 3866 1384 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04113 vss 3664 1382 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04112 1965 1384 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04111 3500 3616 3499 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04110 3499 5745 3611 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04109 vss 4018 3500 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04108 3610 3611 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04107 1864 1973 1863 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04106 1863 1972 1974 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04105 vss 3442 1864 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04104 1971 1974 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04103 3309 3314 3373 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04102 vss 3547 3309 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04101 3310 3312 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04100 vss 3310 3311 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04099 3373 3313 3310 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04098 3547 3373 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04097 vss 3373 3547 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04096 3311 3313 3312 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04095 3312 3314 3374 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04094 vss 6580 3314 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04093 3313 3314 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04092 vss 3548 3375 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04091 3374 3375 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04090 1873 1989 1874 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04089 1874 1988 1987 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04088 vss 1990 1873 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04087 2623 1987 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04086 2646 2944 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04085 2734 3572 2646 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04084 vss 2733 2734 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04083 2678 5069 2677 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04082 2677 2830 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04081 2676 2799 2678 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04080 3414 2800 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04079 2800 6440 2676 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04078 3955 6791 3882 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04077 3881 4157 3955 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04076 3882 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04075 3953 3955 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04074 vss 6637 3881 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04073 3881 4643 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04072 165 254 246 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04071 vss 522 165 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04070 248 249 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04069 vss 248 166 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04068 246 251 248 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04067 522 246 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04066 vss 246 522 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04065 166 251 249 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04064 249 254 167 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04063 vss 3259 254 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04062 251 254 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04061 vss 387 252 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04060 167 252 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04059 1532 1534 1429 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04058 1429 3210 1532 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04057 vss 2349 1429 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04056 1530 1532 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04055 6448 6963 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04054 vss 6974 6448 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04053 4678 4676 4677 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04052 4677 6600 4678 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04051 vss 6601 4677 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04050 4675 4678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04049 5023 6876 5024 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04048 5024 6877 5023 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04047 vss 5670 5024 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04046 5022 5023 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04045 5800 5791 5574 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04044 5574 5792 5800 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04043 vss 5573 5574 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04042 4215 4213 4214 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04041 4214 4212 4215 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04040 vss 4687 4214 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04039 4520 4083 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04038 vss 4075 4520 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04037 4520 4082 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04036 vss 6242 4520 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04035 356 363 355 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04034 vss 502 356 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04033 357 358 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04032 vss 357 359 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04031 355 362 357 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04030 502 355 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04029 vss 355 502 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04028 359 362 358 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04027 358 363 360 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04026 vss 3160 363 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04025 362 363 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04024 vss 364 361 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04023 360 361 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04022 vss 6682 6684 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04021 vss 6694 6684 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04020 6684 6934 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04019 6680 6684 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04018 1444 1968 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04017 2349 1559 1444 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04016 vss 2292 2084 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04015 2084 2304 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04014 2921 2085 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04013 2084 2291 2085 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04012 2085 2498 2084 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04011 1797 2092 1798 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04010 1798 1884 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04009 1886 2303 1797 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04008 3909 4452 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04007 4013 4051 3909 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04006 5099 5552 5100 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04005 5100 5329 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04004 5264 5116 5099 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04003 590 1652 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04002 589 1508 590 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04001 6962 6974 6964 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04000 vss 6963 6965 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03999 6964 6965 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03998 1748 2399 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03997 1973 1757 1748 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03996 1119 1975 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03995 1972 1234 1119 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03994 4010 3792 3496 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03993 3496 3793 4010 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03992 vss 3604 3496 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03991 1408 1635 1407 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03990 1407 1490 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03989 1491 1498 1408 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03988 1403 1483 1404 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03987 1404 1627 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03986 1484 1482 1403 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03985 3184 2519 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03984 vss 2536 3184 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03983 3184 2522 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03982 vss 2518 3184 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03981 1369 2787 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03980 vss 6469 1369 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03979 1369 1745 1565 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03978 1565 1989 1369 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03977 5960 6423 5962 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03976 5962 6374 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03975 5961 6375 5960 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03974 6177 6522 5961 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03973 2605 2603 2606 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03972 2606 3242 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03971 2820 2604 2605 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03970 2556 4220 2557 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03969 2557 3226 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03968 3186 4485 2556 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03967 5662 6917 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03966 5772 6963 5662 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03965 1357 1580 1358 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03964 1358 1749 1357 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03963 vss 4524 1358 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03962 2534 1357 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03961 698 947 697 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03960 697 941 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03959 933 1169 698 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03958 1790 2727 1791 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03957 1791 1877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03956 2286 1876 1790 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03955 5933 6347 5935 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03954 5935 5932 5934 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03953 vss 5937 5933 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03952 5931 5934 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03951 6056 6177 6055 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03950 6055 6176 6179 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03949 vss 6393 6056 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03948 6175 6179 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03947 5206 6226 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03946 5493 6426 5206 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03945 5205 5299 5493 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03944 vss 6220 5205 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03943 5205 5300 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03942 3022 5068 3020 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03941 3020 3023 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03940 3021 5069 3022 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03939 1472 3866 1473 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03938 1473 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03937 1471 3849 1472 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03936 1587 3664 1471 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03935 3767 6434 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03934 3766 6919 3767 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03933 3765 4308 3766 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03932 vss 4217 3765 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03931 3765 5502 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03930 3854 3853 3855 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03929 3855 3856 3857 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03928 vss 4524 3854 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03927 4075 3857 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03926 5656 5773 5655 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03925 5655 5877 5751 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03924 vss 6440 5656 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03923 6183 5751 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03922 vss 6440 6005 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03921 6005 6238 6006 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03920 6004 6006 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03919 1729 2058 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03918 vss 1740 1729 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03917 1729 1728 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03916 vss 1727 1729 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03915 2156 1729 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03914 627 3193 628 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03913 628 794 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03912 626 624 627 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03911 791 625 626 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03910 1463 3866 1462 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03909 1462 2352 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03908 1461 3849 1463 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03907 1578 3664 1461 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03906 1951 2379 1819 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03905 1819 2381 1951 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03904 vss 4748 1819 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03903 2350 1951 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03902 939 1146 940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03901 940 1156 939 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03900 vss 2086 940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03899 938 939 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03898 5460 6791 5459 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03897 5458 5699 5460 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03896 5459 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03895 5456 5460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03894 vss 6637 5458 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03893 5458 5695 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03892 vss 2604 2257 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03891 2257 2603 2398 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03890 2823 2398 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03889 vss 2951 2555 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03888 2555 2553 2554 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03887 2551 2554 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03886 vss 2345 2132 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03885 2132 2344 2133 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03884 2129 2133 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03883 4744 5349 4743 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03882 4743 5992 4744 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03881 vss 5889 4743 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03880 4061 4275 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03879 vss 4059 4061 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03878 4061 4708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03877 vss 6224 4061 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03876 5538 4061 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03875 1646 2106 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03874 1645 2498 1646 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03873 1644 2736 1645 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03872 vss 2111 1644 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03871 1643 2535 1645 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03870 vss 3217 1643 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03869 vss 5069 3803 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03868 3803 5068 3804 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03867 3805 3804 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03866 vss 2329 2229 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03865 2229 2353 2330 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03864 2517 2330 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03863 5197 5291 5283 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03862 vss 5804 5197 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03861 5285 5286 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03860 vss 5285 5198 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03859 5283 5290 5285 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03858 5804 5283 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03857 vss 5283 5804 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03856 5198 5290 5286 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03855 5286 5291 5199 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03854 vss 6832 5291 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03853 5290 5291 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03852 vss 5292 5288 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03851 5199 5288 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03850 4311 4384 4839 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03849 vss 6665 4311 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03848 4310 5914 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03847 4839 4382 4310 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03846 vss 5914 4384 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03845 4382 6665 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03844 6090 6702 6091 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03843 6091 6701 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03842 6089 6704 6090 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03841 6957 6240 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03840 6240 6700 6089 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03839 2072 2396 2073 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03838 2073 2074 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03837 2071 2070 2072 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03836 2603 2179 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03835 2179 2506 2071 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03834 4230 4703 4231 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03833 4231 4228 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03832 4229 4925 4230 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03831 4226 4227 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03830 4227 4238 4229 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03829 vss 4710 4709 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03828 4710 5349 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03827 4709 4708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03826 vss 3814 3012 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03825 3012 3816 3013 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03824 3010 3013 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03823 4728 5773 4727 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03822 4727 4726 4729 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03821 vss 6440 4728 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03820 4725 4729 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03819 1834 2406 1833 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03818 1833 2407 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03817 1832 5359 1834 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03816 1986 3836 1832 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03815 1757 3263 1756 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03814 vss 3460 1759 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03813 1756 1759 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03812 1479 1480 1401 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03811 1401 1478 1479 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03810 vss 1620 1401 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03809 4324 4437 4429 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03808 vss 5959 4324 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03807 4430 4432 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03806 vss 4430 4325 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03805 4429 4435 4430 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03804 5959 4429 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03803 vss 4429 5959 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03802 4325 4435 4432 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03801 4432 4437 4326 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03800 vss 5054 4437 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03799 4435 4437 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03798 vss 4434 4436 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03797 4326 4436 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03796 4661 4657 4857 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03795 vss 4853 4661 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03794 4660 4658 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03793 4857 4659 4660 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03792 vss 4658 4657 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03791 4659 4853 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03790 6222 6224 6078 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03789 6078 6221 6222 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03788 vss 6702 6078 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03787 429 615 428 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03786 428 493 492 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03785 vss 2314 429 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03784 491 492 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03783 4716 5992 4719 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03782 4719 4726 4718 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03781 vss 6440 4716 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03780 4715 4718 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03779 3142 3369 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03778 3451 3371 3142 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03777 3141 3455 3451 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03776 vss 3456 3141 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03775 3141 3457 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03774 vss 5575 5109 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03773 5109 5341 5108 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03772 5986 5108 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03771 3761 5967 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03770 vss 5993 3761 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03769 4016 4213 3908 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03768 3908 4212 4016 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03767 vss 5064 3908 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03766 5859 5949 5446 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03765 5446 5947 5859 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03764 vss 5965 5446 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03763 1436 1552 1544 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03762 vss 3604 1436 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03761 1545 1548 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03760 vss 1545 1438 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03759 1544 1551 1545 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03758 3604 1544 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03757 vss 1544 3604 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03756 1438 1551 1548 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03755 1548 1552 1437 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03754 vss 3259 1552 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03753 1551 1552 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03752 vss 1549 1550 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03751 1437 1550 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03750 vss 1327 1517 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03749 1327 1326 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03748 1517 1328 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03747 963 960 1518 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03746 vss 961 963 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03745 964 1313 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03744 1518 962 964 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03743 vss 1313 960 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03742 962 961 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03741 4378 4507 4377 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03740 4377 5345 4508 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03739 vss 4505 4378 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03738 4506 4508 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03737 2619 4276 2618 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03736 2618 4089 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03735 2617 4286 2619 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03734 4491 2616 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03733 2616 3866 2617 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03732 5907 5893 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03731 6471 6728 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03730 6226 6480 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03729 6025 6261 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03728 5888 6571 5890 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03727 5890 5889 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03726 5887 5992 5888 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03725 5998 5997 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03724 5997 6440 5887 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03723 4172 6434 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03722 4171 6919 4172 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03721 4170 6265 4171 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03720 vss 4217 4170 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03719 4170 5502 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03718 954 955 1309 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03717 vss 953 954 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03716 957 2999 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03715 1309 956 957 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03714 vss 2999 955 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03713 956 953 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03712 3788 3792 3787 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03711 3787 3793 3788 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03710 vss 3796 3787 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03709 6023 6263 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03708 3658 4299 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03707 vss 5157 3658 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03706 vss 2737 2749 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03705 2749 2535 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03704 vss 2355 2749 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03703 6609 6876 6506 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03702 6506 6877 6609 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03701 vss 6820 6506 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03700 169 3229 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03699 261 845 169 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03698 722 843 836 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03697 vss 3423 722 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03696 837 840 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03695 vss 837 723 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03694 836 842 837 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03693 3423 836 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03692 vss 836 3423 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03691 723 842 840 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03690 840 843 724 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03689 vss 3259 843 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03688 842 843 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03687 vss 1007 841 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03686 724 841 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03685 5486 6434 5484 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03684 5484 6431 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03683 5485 6919 5486 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03682 6498 6593 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03681 6589 6588 6498 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03680 6597 6598 6502 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03679 6502 6600 6597 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03678 vss 6601 6502 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03677 6596 6597 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03676 6544 6691 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03675 6690 6921 6544 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03674 2545 986 443 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03673 443 987 2545 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03672 vss 663 443 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03671 972 4176 971 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03670 971 1322 972 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03669 vss 2747 971 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03668 981 972 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03667 1635 1885 1634 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03666 1634 1891 1635 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03665 vss 1882 1634 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03664 vss 5277 5194 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03663 5194 5279 5278 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03662 6364 5278 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03661 6648 6876 6532 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03660 6532 6877 6648 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03659 vss 6885 6532 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03658 vss 302 304 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_03657 304 312 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_03656 301 303 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03655 304 305 303 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_03654 303 2498 304 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_03653 334 784 333 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03652 333 494 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03651 332 2314 334 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03650 2651 2940 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03649 2741 2938 2651 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03648 3018 3816 3019 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03647 3019 3631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03646 3199 3814 3018 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03645 171 1231 172 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03644 172 1732 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03643 263 4501 171 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03642 1688 986 441 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03641 441 987 1688 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03640 vss 502 441 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03639 6504 6608 6607 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03638 vss 6820 6504 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03637 6505 6814 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03636 6607 6605 6505 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03635 vss 6814 6608 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03634 6605 6820 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03633 3991 4217 3898 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03632 3898 5502 3991 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03631 vss 6727 3898 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03630 vss 3438 3106 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03629 3106 3225 3220 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03628 3976 3220 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03627 4898 6220 4781 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03626 4781 5300 4898 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03625 vss 4897 4781 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03624 4896 4898 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03623 vss 6665 5169 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03622 5169 5914 5246 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03621 5245 5246 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03620 2200 2198 2201 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03619 2201 2207 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03618 2199 3062 2200 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03617 2408 3060 2199 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03616 vss 2841 4087 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03615 2841 5363 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03614 4087 4094 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03613 3742 5299 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03612 3741 3740 3742 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03611 3739 6265 3741 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03610 vss 3737 3739 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03609 3739 3738 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03608 1063 1153 1490 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03607 vss 1647 1063 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03606 1064 1298 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03605 1490 1154 1064 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03604 vss 1298 1153 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03603 1154 1647 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03602 5364 5371 5365 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03601 5239 5373 5364 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03600 5363 5364 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03599 vss 5364 5363 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03598 5242 5370 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03597 vss 5369 5370 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03596 5371 5373 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03595 vss 6984 5373 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03594 5240 5367 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03593 5365 6976 5240 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03592 5367 5373 5242 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03591 5241 5371 5367 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03590 vss 5365 5241 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03589 vss 5363 5238 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03588 5238 6976 5239 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03587 4394 5044 4169 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03586 4169 5045 4394 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03585 vss 5927 4169 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03584 6080 6226 6079 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03583 6079 6691 6227 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03582 vss 6921 6080 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03581 6225 6227 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03580 1353 1580 1354 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03579 1354 1749 1353 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03578 vss 4524 1354 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03577 vss 2520 2322 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03576 2322 2740 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03575 2323 2322 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03574 4773 5269 4774 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03573 4774 4878 4879 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03572 vss 5456 4773 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03571 4876 4879 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03570 2826 2823 2693 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03569 2693 5792 2826 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03568 vss 2824 2693 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03567 2607 1033 1034 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03566 1034 1223 2607 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03565 vss 1732 1034 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03564 1107 1572 1108 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03563 1108 1381 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03562 1106 1367 1107 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03561 2797 1220 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03560 1220 2070 1106 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03559 4365 4453 4364 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03558 4364 4460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03557 4363 4455 4365 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03556 6375 4454 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03555 4454 4472 4363 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03554 vss 965 967 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03553 967 968 966 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03552 3178 966 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03551 757 3217 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03550 787 1904 757 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03549 756 3188 787 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03548 vss 2746 756 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03547 756 1322 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03546 5943 6876 5941 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03545 5941 6877 5943 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03544 vss 6740 5941 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03543 5011 6876 5010 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03542 5010 6877 5011 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03541 vss 6665 5010 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03540 412 2727 411 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03539 411 579 462 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03538 vss 1876 412 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03537 466 462 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03536 3112 5575 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03535 3233 4726 3112 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03534 3111 4053 3233 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03533 vss 5773 3111 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03532 3110 4524 3233 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03531 vss 3229 3110 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03530 5964 3634 3441 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03529 3441 3632 5964 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03528 vss 3442 3441 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03527 1745 2194 1116 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03526 1116 2195 1745 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03525 vss 6440 1116 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03524 5447 5457 5448 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03523 vss 5501 5447 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03522 5449 5452 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03521 vss 5449 5451 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03520 5448 5454 5449 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03519 5501 5448 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03518 vss 5448 5501 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03517 5451 5454 5452 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03516 5452 5457 5450 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03515 vss 6832 5457 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03514 5454 5457 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03513 vss 5453 5455 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03512 5450 5455 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03511 4175 4880 4174 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03510 4174 4881 4175 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03509 vss 5927 4174 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03508 6439 6714 6441 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03507 6441 6440 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03506 6437 6952 6439 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03505 6691 6438 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03504 6438 6963 6437 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03503 vss 2799 2176 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03502 2176 2399 2177 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03501 2174 2177 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03500 vss 3003 3005 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03499 3005 3429 3007 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03498 3004 3007 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03497 4357 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03496 4685 6431 4357 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03495 4356 4438 4685 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03494 vss 6220 4356 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03493 4356 5300 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03492 3077 3151 3144 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03491 vss 3709 3077 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03490 3145 3147 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03489 vss 3145 3078 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03488 3144 3150 3145 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03487 3709 3144 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03486 vss 3144 3709 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03485 3078 3150 3147 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03484 3147 3151 3079 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03483 vss 3160 3151 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03482 3150 3151 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03481 vss 3712 3149 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03480 3079 3149 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03479 2162 3006 2163 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03478 2163 3217 2164 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03477 vss 3010 2162 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03476 2161 2164 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03475 3959 6791 3884 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03474 3883 3962 3959 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03473 3884 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03472 3957 3959 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03471 vss 6637 3883 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03470 3883 4160 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03469 4805 4941 4806 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03468 4806 4942 4934 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03467 vss 5773 4805 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03466 5756 4934 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03465 3839 4286 3838 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03464 3838 4941 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03463 3837 3836 3839 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03462 4250 3835 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03461 3835 4524 3837 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03460 1858 1953 1860 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03459 1860 2194 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03458 1859 2125 1858 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03457 2514 1954 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03456 1954 3836 1859 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03455 5860 5931 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03454 5861 5859 5860 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03453 6417 5967 5613 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03452 5613 5993 6417 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03451 vss 5948 5613 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03450 5270 4673 4323 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03449 4323 4671 5270 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03448 vss 5948 4323 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03447 378 386 379 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03446 vss 825 378 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03445 380 382 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03444 vss 380 381 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03443 379 384 380 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03442 825 379 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03441 vss 379 825 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03440 381 384 382 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03439 382 386 383 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03438 vss 3259 386 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03437 384 386 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03436 vss 517 385 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03435 383 385 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03434 6479 6974 6478 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03433 6478 6477 6479 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03432 vss 6480 6478 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03431 6725 6479 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03430 vss 4695 4604 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03429 4604 5089 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03428 vss 4919 4604 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03427 1334 1340 1335 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03426 1335 3408 1334 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03425 vss 2534 1335 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03424 1333 1334 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03423 5008 6876 5009 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03422 5009 6877 5008 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03421 vss 5670 5009 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03420 2074 4213 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03419 vss 2174 2074 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03418 2074 3051 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03417 vss 2188 2074 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03416 1778 3460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03415 vss 3263 1778 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03414 4590 4876 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03413 4589 4672 4590 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03412 3971 4673 3890 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03411 3890 4671 3971 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03410 vss 3969 3890 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03409 6143 6172 5929 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03408 5929 6173 6143 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03407 vss 5965 5929 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03406 1336 1340 1337 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03405 1337 3408 1336 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03404 vss 2349 1337 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03403 1338 1336 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03402 vss 4087 3535 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03401 3535 3660 3659 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03400 3856 3659 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03399 1447 1968 1448 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03398 1448 1558 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03397 1728 1559 1447 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03396 2049 2544 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03395 2136 2142 2049 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03394 3532 3653 3533 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03393 3533 3654 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03392 3655 3652 3532 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03391 1460 2406 1459 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03390 1459 2412 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03389 1458 5359 1460 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03388 1758 4501 1458 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03387 6978 6986 6979 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03386 6973 6988 6978 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03385 6974 6978 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03384 vss 6978 6974 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03383 6983 6985 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03382 vss 6981 6985 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03381 6986 6988 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03380 vss 6984 6988 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03379 6977 6982 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03378 6979 6976 6977 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03377 6982 6988 6983 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03376 6980 6986 6982 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03375 vss 6979 6980 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03374 vss 6974 6975 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03373 6975 6976 6973 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03372 4646 4918 4648 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03371 4648 5014 4647 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03370 vss 5026 4646 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03369 4658 4647 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03368 vss 4233 4234 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03367 4234 5102 4236 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03366 6422 4236 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03365 1660 1904 1659 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03364 1659 1737 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03363 1661 2375 1660 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03362 vss 2755 2121 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03361 2121 3586 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03360 2135 2121 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03359 2580 5069 2581 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03358 2581 2807 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03357 2587 5773 2580 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03356 2629 5363 2077 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03355 vss 3263 2078 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03354 2077 2078 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03353 2113 3217 2112 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03352 2112 2506 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03351 2114 2501 2113 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03350 2111 2782 2114 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03349 2099 3740 2100 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03348 2100 2512 2099 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03347 vss 2314 2100 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03346 2299 2099 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03345 3238 4083 3115 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03344 3115 4082 3238 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03343 vss 6265 3115 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03342 6501 6594 6500 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03341 6500 6596 6595 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03340 vss 6798 6501 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03339 6593 6595 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03338 vss 2402 2404 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03337 2402 5349 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03336 2404 5157 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03335 3558 6172 3476 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03334 3476 6173 3558 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03333 vss 3969 3476 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03332 4787 5068 4786 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03331 4786 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03330 4785 5069 4787 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03329 5062 4902 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03328 4902 5902 4785 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03327 6468 6466 6467 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03326 6465 6694 6468 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03325 6467 6476 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03324 6463 6468 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03323 vss 6464 6465 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03322 6465 6690 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03321 vss 961 959 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03320 959 1313 958 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03319 1165 958 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03318 2273 2412 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03317 2622 4089 2273 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03316 2274 4941 2622 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03315 vss 2415 2274 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03314 2272 2411 2622 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03313 vss 2615 2272 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03312 1148 1488 1060 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03311 1060 1485 1148 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03310 vss 1490 1060 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03309 1146 1148 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03308 4591 4880 4322 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03307 4322 4881 4591 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03306 vss 5965 4322 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03305 1959 1735 1736 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03304 1736 1950 1959 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03303 vss 2801 1736 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03302 6958 6957 6960 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03301 6960 6959 6961 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03300 vss 6974 6958 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03299 6972 6961 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03298 1041 1039 1040 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03297 1040 1229 1042 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03296 vss 1038 1041 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03295 2604 1042 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03294 1344 2544 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03293 1343 2142 1344 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03292 vss 1353 1343 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03291 vss 1215 1018 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03290 1018 1214 1017 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03289 1210 1017 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03288 vss 682 684 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03287 684 859 683 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03286 844 683 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03285 vss 1491 1284 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03284 1284 1292 1283 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03283 1480 1283 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03282 6626 6876 6517 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03281 6517 6877 6626 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03280 vss 6740 6517 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03279 6624 6626 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03278 4828 4963 4955 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03277 vss 5359 4828 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03276 4957 4960 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03275 vss 4957 4829 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03274 4955 4964 4957 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03273 5359 4955 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03272 vss 4955 5359 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03271 4829 4964 4960 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03270 4960 4963 4830 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03269 vss 6984 4963 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03268 4964 4963 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03267 vss 4961 4962 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03266 4830 4962 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03265 5074 5081 5075 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03264 vss 5742 5074 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03263 5076 5077 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03262 vss 5076 5078 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03261 5075 5082 5076 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03260 5742 5075 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03259 vss 5075 5742 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03258 5078 5082 5077 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03257 5077 5081 5079 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03256 vss 6984 5081 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03255 5082 5081 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03254 vss 5306 5080 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03253 5079 5080 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03252 6640 6876 6394 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03251 6394 6877 6640 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03250 vss 6893 6394 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03249 5911 5909 6128 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03248 vss 5910 5911 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03247 5913 5914 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03246 6128 5912 5913 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03245 vss 5914 5909 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03244 5912 5910 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03243 2265 3866 2264 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03242 2264 4286 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03241 2263 2406 2265 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03240 4509 3836 2263 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03239 vss 1224 1112 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03238 1112 1221 1222 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03237 1365 1222 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03236 1806 2375 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03235 1902 1904 1806 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03234 vss 2382 1902 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03233 2319 1902 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03232 3131 5064 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03231 3172 3740 3131 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03230 3130 5902 3172 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03229 vss 3737 3130 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03228 3130 3738 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03227 6527 6645 6644 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03226 vss 6906 6527 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03225 6528 6893 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03224 6644 6642 6528 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03223 vss 6893 6645 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03222 6642 6906 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03221 5093 5749 5092 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03220 5092 5748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03219 5091 6740 5093 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03218 5089 5090 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03217 5090 6440 5091 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03216 vss 2407 2262 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03215 2262 2404 2405 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03214 2830 2405 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03213 748 1479 747 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03212 747 936 763 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03211 vss 933 748 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03210 769 763 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03209 5047 5056 5048 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03208 vss 5958 5047 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03207 5049 5050 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03206 vss 5049 5051 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03205 5048 5055 5049 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03204 5958 5048 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03203 vss 5048 5958 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03202 5051 5055 5050 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03201 5050 5056 5052 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03200 vss 5054 5056 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03199 5055 5056 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03198 vss 5057 5053 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03197 5052 5053 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03196 4654 4652 4653 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03195 vss 4914 4654 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03194 4656 4658 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03193 4653 4655 4656 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03192 vss 4658 4652 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03191 4655 4914 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03190 4734 6469 4735 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03189 4735 4733 4734 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03188 vss 4731 4735 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03187 4732 4734 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03186 700 768 5044 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03185 vss 766 700 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03184 701 1313 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03183 5044 765 701 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03182 vss 1313 768 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03181 765 766 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03180 vss 4517 4515 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03179 4515 4622 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03178 vss 6000 4515 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03177 6447 5272 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03176 4676 4308 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03175 4176 5243 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03174 2746 5262 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03173 6598 6265 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03172 6603 6727 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03171 4089 3460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03170 vss 2852 4089 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03169 vss 4083 3245 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03168 3245 3246 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03167 vss 4082 3245 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03166 2240 2372 2364 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03165 vss 3421 2240 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03164 2365 2367 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03163 vss 2365 2241 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03162 2364 2369 2365 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03161 3421 2364 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03160 vss 2364 3421 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03159 2241 2369 2367 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03158 2367 2372 2242 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03157 vss 3259 2372 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03156 2369 2372 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03155 vss 2560 2370 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03154 2242 2370 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03153 2958 2965 2959 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03152 2955 2966 2958 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03151 3190 2958 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03150 vss 2958 3190 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03149 2963 2964 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03148 vss 2961 2964 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03147 2965 2966 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03146 vss 3160 2966 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03145 2957 2962 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03144 2959 6976 2957 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03143 2962 2966 2963 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03142 2960 2965 2962 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03141 vss 2959 2960 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03140 vss 3190 2956 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03139 2956 6976 2955 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03138 506 986 442 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03137 442 987 506 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03136 vss 504 442 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03135 1189 506 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03134 4032 3423 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03133 5705 6591 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03132 4853 4914 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03131 3800 3790 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03130 2562 3199 2558 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03129 2558 3618 2562 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03128 vss 5742 2558 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03127 5540 5986 5541 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03126 5541 6214 5540 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03125 vss 6906 5541 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03124 vss 4520 4630 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03123 4630 4521 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03122 vss 4518 4630 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03121 6034 6800 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03120 6786 6132 6034 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03119 6077 6701 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03118 6220 6702 6077 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03117 1843 1880 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03116 2896 1883 1843 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03115 1402 2896 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03114 1875 2897 1402 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03113 4851 6876 4762 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03112 4762 6877 4851 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03111 vss 5026 4762 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03110 4850 4851 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03109 vss 6970 6971 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03108 6971 6972 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03107 6981 6971 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03106 1638 1639 1884 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03105 vss 2097 1638 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03104 1637 1641 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03103 1884 1636 1637 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03102 vss 1641 1639 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03101 1636 2097 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03100 1633 1632 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03099 2897 1886 1633 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03098 6812 6816 6817 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03097 vss 6811 6812 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03096 6815 6814 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03095 6817 6813 6815 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03094 vss 6814 6816 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03093 6813 6811 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03092 4594 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03091 4688 6431 4594 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03090 4593 4687 4688 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03089 vss 6220 4593 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03088 4593 5300 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03087 578 576 580 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03086 580 579 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03085 577 2727 578 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03084 870 1876 577 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03083 3411 3413 3412 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03082 3412 3414 3411 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03081 vss 4308 3412 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03080 3600 3411 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03079 398 4524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03078 845 4748 398 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03077 vss 3858 4276 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03076 3858 4748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03075 4276 4094 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03074 707 2161 706 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03073 706 2498 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03072 2314 1900 707 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03071 406 2615 407 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03070 407 2411 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03069 405 3460 406 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03068 456 1231 457 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03067 457 1732 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03066 682 4748 456 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03065 1296 1299 1483 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03064 vss 1501 1296 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03063 1297 1298 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03062 1483 1295 1297 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03061 vss 1298 1299 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03060 1295 1501 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03059 2516 2535 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03058 2525 2737 2516 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03057 vss 3991 3899 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03056 3899 4452 3992 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03055 4150 3992 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03054 5067 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03053 5065 6685 5067 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03052 5066 5064 5065 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03051 vss 6220 5066 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03050 5066 5300 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03049 vss 4482 4334 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03048 4334 4483 4484 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03047 5154 4484 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03046 1588 2852 1474 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03045 vss 3460 1589 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03044 1474 1589 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03043 1785 1991 1786 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03042 1786 2352 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03041 1784 4094 1785 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03040 1990 5363 1784 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03039 1772 4089 1773 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03038 1773 2352 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03037 1771 4087 1772 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03036 1989 4299 1771 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03035 5542 5748 5543 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03034 5543 5545 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03033 5758 6906 5542 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03032 vss 5993 2385 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03031 2385 5967 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03030 2386 2385 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03029 6402 6401 6403 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03028 6403 6405 6404 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03027 vss 6660 6402 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03026 6400 6404 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03025 vss m_clock 3419 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03024 5334 3419 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03023 vss 3419 5334 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03022 vss 3419 5334 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03021 5334 3419 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03020 vss 5334 5335 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03019 6984 5335 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03018 vss 5335 6984 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03017 vss 5335 6984 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03016 6984 5335 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03015 vss 5334 5333 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03014 5332 5333 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03013 vss 5333 5332 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03012 vss 5333 5332 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03011 5332 5333 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03010 vss 5334 5122 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03009 5121 5122 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03008 vss 5122 5121 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03007 vss 5122 5121 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03006 5121 5122 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03005 vss 5334 5267 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03004 6832 5267 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03003 vss 5267 6832 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03002 vss 5267 6832 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03001 6832 5267 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03000 vss 5334 5266 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02999 6580 5266 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02998 vss 5266 6580 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02997 vss 5266 6580 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02996 6580 5266 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02995 978 918 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02994 vss 3210 978 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02993 978 2537 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02992 vss 919 978 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02991 1176 978 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02990 vss 6974 6218 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02989 6218 6963 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02988 6219 6218 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02987 vss 4708 4730 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02986 4730 6224 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02985 4731 4730 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02984 2645 2944 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02983 2731 3572 2645 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02982 vss 2733 2731 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02981 2730 2731 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02980 1184 1194 1085 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02979 1085 1190 1184 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02978 vss 1182 1085 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02977 1919 1184 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02976 2118 2512 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02975 2513 2511 2118 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02974 vss 2117 2513 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02973 4596 5068 4597 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02972 4597 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02971 4595 5069 4596 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02970 4692 4691 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02969 4691 5243 4595 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02968 5864 5044 5046 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02967 5046 5045 5864 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02966 vss 6188 5046 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02965 1288 1900 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02964 1287 2161 1288 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02963 1286 1490 1287 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02962 vss 1488 1286 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02961 1286 1485 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02960 4047 4275 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02959 vss 4043 4047 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02958 4047 4708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02957 vss 6224 4047 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02956 5327 4047 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02955 4180 6434 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02954 4181 6919 4180 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02953 4179 5272 4181 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02952 vss 4217 4179 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02951 4179 5502 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02950 5591 5692 5684 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02949 vss 5936 5591 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02948 5686 5689 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02947 vss 5686 5592 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02946 5684 5691 5686 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02945 5936 5684 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02944 vss 5684 5936 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02943 5592 5691 5689 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02942 5689 5692 5593 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02941 vss 6580 5692 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02940 5691 5692 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02939 vss 5861 5690 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02938 5593 5690 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02937 vss 4932 6678 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02936 4932 4939 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02935 6678 6422 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02934 693 1953 694 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02933 694 2194 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02932 691 3836 693 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02931 690 692 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02930 692 6440 691 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02929 vss 1779 1046 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02928 1046 1991 1047 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02927 1218 1047 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02926 vss 4299 140 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02925 140 405 139 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02924 138 139 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02923 3792 1746 1747 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02922 1747 1745 3792 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02921 vss 2184 1747 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02920 6121 6791 6029 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02919 6028 6123 6121 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02918 6029 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02917 6118 6121 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02916 vss 6637 6028 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02915 6028 6119 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02914 5874 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02913 6401 6685 5874 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02912 5873 5963 6401 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02911 vss 6182 5873 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02910 5873 6183 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02909 6639 6791 6526 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02908 6525 6640 6639 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02907 6526 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02906 6636 6639 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02905 vss 6637 6525 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02904 6525 6644 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02903 4055 5575 3918 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02902 3917 4053 4055 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02901 3918 4726 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02900 5927 4055 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02899 vss 5992 3917 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02898 3917 5773 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02897 4367 5097 4368 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02896 4368 4463 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02895 4366 4701 4367 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02894 4461 4464 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02893 4464 4462 4366 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02892 419 475 473 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02891 vss 1505 419 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02890 420 1652 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02889 473 472 420 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02888 vss 1652 475 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02887 472 1505 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02886 1067 1647 1068 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02885 1068 1320 1159 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02884 vss 2314 1067 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02883 1158 1159 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02882 2462 2469 2461 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02881 vss 3946 2462 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02880 2463 2465 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02879 vss 2463 2464 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02878 2461 2468 2463 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02877 3946 2461 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02876 vss 2461 3946 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02875 2464 2468 2465 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02874 2465 2469 2466 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02873 vss 3160 2469 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02872 2468 2469 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02871 vss 3949 2467 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02870 2466 2467 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02869 3927 4941 3928 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02868 3928 4942 4067 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02867 vss 5349 3927 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02866 5749 4067 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02865 3842 4276 3843 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02864 3843 4941 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02863 3841 4286 3842 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02862 4726 3840 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02861 3840 4524 3841 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02860 31 105 101 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02859 vss 636 31 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02858 32 34 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02857 vss 32 33 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02856 101 35 32 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02855 636 101 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02854 vss 101 636 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02853 33 35 34 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02852 34 105 104 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02851 vss 3160 105 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02850 35 105 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02849 vss 225 106 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02848 104 106 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02847 772 911 702 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02846 702 769 772 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02845 vss 770 702 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02844 1392 1992 1393 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02843 1393 1394 1392 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02842 vss 2198 1393 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02841 1390 1392 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02840 1827 5992 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02839 1967 4053 1827 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02838 1826 1965 1967 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02837 vss 1982 1826 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02836 1825 3229 1967 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02835 vss 2125 1825 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02834 1113 1732 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02833 2070 1223 1113 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02832 2214 2295 2298 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02831 vss 2489 2214 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02830 2215 2299 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02829 2298 2296 2215 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02828 vss 2299 2295 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02827 2296 2489 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02826 3388 3339 3332 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02825 3331 3340 3388 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02824 3395 3388 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02823 vss 3388 3395 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02822 3336 3338 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02821 vss 3337 3338 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02820 3339 3340 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02819 vss 5054 3340 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02818 3333 3335 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02817 3332 6976 3333 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02816 3335 3340 3336 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02815 3334 3339 3335 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02814 vss 3332 3334 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02813 vss 3395 3330 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02812 3330 6976 3331 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02811 5863 6362 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02810 6139 5862 5863 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02809 vss 3798 3799 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02808 vss 3969 3799 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02807 3799 4611 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02806 3797 3799 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02805 3889 6434 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02804 3967 6919 3889 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02803 3888 5902 3967 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02802 vss 4217 3888 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02801 3888 5502 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02800 5021 6919 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02799 5440 6434 5021 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02798 5020 6867 5440 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02797 vss 5019 5020 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02796 5020 5022 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02795 6097 6476 6098 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02794 6098 6243 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02793 6706 6242 6097 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02792 1536 1534 1430 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02791 1430 3210 1536 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02790 vss 2521 1430 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02789 1533 1536 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02788 2909 2915 2639 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02787 2639 2716 2909 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02786 vss 2717 2639 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02785 3119 5157 3120 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02784 3120 3263 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02783 3458 5363 3119 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02782 4592 5034 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02781 4873 4591 4592 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02780 5956 6806 5957 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02779 5957 6631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02778 5955 6591 5956 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02777 5236 5788 5235 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02776 5235 5570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02775 5361 5359 5236 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02774 1395 1992 1396 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02773 1396 1394 1395 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02772 vss 2198 1396 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02771 3448 3455 3447 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02770 3446 3863 3448 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02769 3447 3449 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02768 3639 3448 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02767 vss 4071 3446 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02766 3446 3458 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02765 3442 2180 1829 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02764 1829 1979 3442 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02763 vss 2193 1829 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02762 2239 3793 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02761 2355 2352 2239 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02760 6370 6806 6373 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02759 6373 6631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02758 6371 6740 6370 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02757 6379 6423 6378 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02756 6378 6374 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02755 6377 6375 6379 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02754 6372 6376 6377 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02753 vss 6906 6536 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02752 6536 6893 6659 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02751 6890 6659 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02750 4810 4946 4809 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02749 4809 5549 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02748 6420 4947 4810 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02747 1124 1234 1123 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02746 1123 1975 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02745 1235 1233 1124 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02744 1306 1300 703 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02743 703 776 1306 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02742 vss 870 703 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02741 vss 2346 2339 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02740 2339 2340 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02739 4881 2339 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02738 66 335 67 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02737 67 310 66 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02736 vss 607 67 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02735 307 66 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02734 3608 3792 3498 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02733 3498 3793 3608 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02732 vss 3607 3498 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02731 1019 1953 1020 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02730 1020 2194 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02729 1560 3836 1019 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02728 vss 6686 6919 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02727 6686 6974 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02726 6919 6963 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02725 941 1146 942 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02724 942 1156 941 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02723 vss 2086 942 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02722 6020 6023 6022 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02721 6022 6261 6021 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02720 vss 6476 6020 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02719 6247 6021 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02718 vss 3866 1754 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02717 1754 4286 1755 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02716 2183 1755 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02715 vss 5363 3066 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02714 3066 4094 3065 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02713 3849 3065 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02712 935 1479 934 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02711 934 936 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02710 2728 933 935 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02709 2475 2727 2474 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02708 2474 2728 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02707 2915 2723 2475 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02706 5637 6342 5638 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02705 5638 5702 5703 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02704 vss 5700 5637 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02703 5701 5703 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02702 4248 4253 4247 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02701 4247 4258 4249 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02700 vss 4616 4248 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02699 4482 4249 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02698 1723 1722 1726 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02697 1726 1724 1725 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02696 vss 1730 1723 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02695 2775 1725 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02694 2819 3037 2691 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02693 2691 2820 2819 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02692 vss 3236 2691 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02691 2817 2819 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02690 vss 4438 3091 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02689 3091 3740 3192 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02688 3191 3192 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02687 1185 1188 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02686 vss 3408 1185 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02685 1185 2770 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02684 vss 1189 1185 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02683 1186 1185 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02682 5761 5753 5617 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02681 5617 5767 5761 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02680 vss 6905 5617 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02679 6357 5949 5950 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02678 5950 5947 6357 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02677 vss 5948 5950 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02676 6455 6461 6456 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02675 6452 6462 6455 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02674 6694 6455 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02673 vss 6455 6694 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02672 6459 6460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02671 vss 6463 6460 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02670 6461 6462 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02669 vss 6984 6462 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02668 6454 6457 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02667 6456 6976 6454 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02666 6457 6462 6459 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02665 6458 6461 6457 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02664 vss 6456 6458 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02663 vss 6694 6453 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02662 6453 6976 6452 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02661 vss 1169 1074 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02660 1074 1313 1170 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02659 2999 1170 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02658 vss 2314 159 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02657 159 493 217 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02656 216 217 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02655 vss 3650 3654 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02654 3650 4080 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02653 3654 3649 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02652 1467 2406 1468 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02651 1468 2407 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02650 1466 5359 1467 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02649 1580 1581 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02648 1581 3836 1466 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02647 5145 5155 5146 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02646 vss 5144 5145 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02645 5147 5149 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02644 vss 5147 5148 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02643 5146 5153 5147 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02642 5144 5146 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02641 vss 5146 5144 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02640 5148 5153 5149 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02639 5149 5155 5150 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02638 vss 6984 5155 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02637 5153 5155 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02636 vss 5151 5152 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02635 5150 5152 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02634 4644 4641 4643 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02633 vss 5026 4644 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02632 4645 5014 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02631 4643 4642 4645 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02630 vss 5014 4641 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02629 4642 5026 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02628 313 314 315 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02627 315 473 316 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02626 vss 476 313 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02625 312 316 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02624 vss 6440 5103 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02623 5103 5349 5105 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02622 5102 5105 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02621 vss 2787 2672 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02620 2672 3617 2789 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02619 2788 2789 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02618 vss 4748 695 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02617 695 4524 696 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02616 857 696 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02615 vss 6440 3024 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02614 3024 5992 3025 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02613 3023 3025 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02612 vss 3818 3820 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02611 3820 5069 3822 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02610 3819 3822 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02609 2542 3199 2541 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02608 2541 3618 2542 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02607 vss 5963 2541 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02606 5478 4899 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02605 vss 4892 5478 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02604 3867 3875 3868 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02603 vss 4094 3867 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02602 3869 3870 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02601 vss 3869 3872 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02600 3868 3873 3869 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02599 4094 3868 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02598 vss 3868 4094 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02597 3872 3873 3870 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02596 3870 3875 3871 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02595 vss 6984 3875 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02594 3873 3875 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02593 vss 4093 3874 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02592 3871 3874 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02591 985 2124 984 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02590 983 2122 985 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02589 984 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02588 980 985 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02587 vss 981 983 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02586 983 982 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02585 vss 5893 5624 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02584 5624 5787 5786 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02583 5784 5786 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02582 vss 5992 4712 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02581 4712 5341 4711 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02580 5753 4711 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02579 vss 2615 459 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02578 459 2411 541 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02577 1033 541 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02576 1988 1779 1780 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02575 1780 4087 1988 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02574 vss 1991 1780 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02573 4182 4190 4183 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02572 vss 6187 4182 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02571 4184 4186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02570 vss 4184 4185 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02569 4183 4189 4184 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02568 6187 4183 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02567 vss 4183 6187 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02566 4185 4189 4186 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02565 4186 4190 4187 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02564 vss 5054 4190 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02563 4189 4190 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02562 vss 4191 4188 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02561 4187 4188 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02560 5661 6921 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02559 5770 6691 5661 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02558 5660 6440 5770 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02557 vss 5999 5660 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02556 5660 6000 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02555 2142 1194 718 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02554 718 1190 2142 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02553 vss 825 718 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02552 2373 2799 2243 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02551 2243 4051 2373 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02550 vss 2790 2243 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02549 2371 2373 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02548 6352 6740 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02547 4163 4918 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02546 4024 3796 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02545 vss 3067 3660 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02544 3067 3263 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02543 3660 3460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02542 vss 3051 1381 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02541 1381 1380 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02540 vss 1749 1381 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02539 2566 2574 2567 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02538 vss 3802 2566 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02537 2568 2570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02536 vss 2568 2571 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02535 2567 2573 2568 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02534 3802 2567 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02533 vss 2567 3802 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02532 2571 2573 2570 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02531 2570 2574 2569 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02530 vss 3259 2574 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02529 2573 2574 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02528 vss 2792 2572 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02527 2569 2572 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02526 vss 3240 3242 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02525 3240 3637 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02524 3242 4083 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02523 781 1904 753 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02522 752 2747 781 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02521 753 3217 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02520 779 781 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02519 vss 4176 752 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02518 752 1322 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02517 3522 4265 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02516 3637 5773 3522 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02515 6811 6820 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02514 4836 5026 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02513 6835 6850 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02512 6112 5524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02511 6695 6694 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02510 6935 6934 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02509 3981 3987 3982 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02508 3894 3989 3981 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02507 3979 3981 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02506 vss 3981 3979 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02505 3897 3988 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02504 vss 3986 3988 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02503 3987 3989 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02502 vss 5054 3989 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02501 3895 3985 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02500 3982 6976 3895 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02499 3985 3989 3897 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02498 3896 3987 3985 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02497 vss 3982 3896 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02496 vss 3979 3893 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02495 3893 6976 3894 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02494 4401 6876 4168 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02493 4168 6877 4401 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02492 vss 4914 4168 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02491 6583 6876 6496 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02490 6496 6877 6583 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02489 vss 6905 6496 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02488 6586 6583 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02487 5101 5329 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02486 5954 5552 5101 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02485 5550 6238 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02484 5551 6440 5550 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02483 1348 2544 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02482 1706 2142 1348 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02481 vss 1356 1706 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02480 4371 4491 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02479 4733 5773 4371 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02478 4224 3604 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02477 5531 5993 5530 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02476 5530 5967 5531 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02475 vss 5964 5530 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02474 1679 1194 1084 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02473 1084 1190 1679 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02472 vss 1182 1084 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02471 3736 4880 3735 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02470 3735 4881 3736 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02469 vss 3969 3735 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02468 vss 5157 4754 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02467 4754 5893 4965 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02466 vss 5893 4833 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02465 4965 4833 4753 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02464 5164 4965 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02463 4753 5372 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02462 vss 3263 3125 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02461 3125 5893 3266 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02460 vss 5893 3267 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02459 3266 3267 3124 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02458 3262 3266 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02457 3124 5262 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02456 vss 4748 4348 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02455 4348 5893 4537 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02454 vss 5893 4538 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02453 4537 4538 4347 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02452 4751 4537 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02451 4347 5243 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02450 vss 4524 4306 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02449 4306 5893 4307 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02448 vss 5893 4309 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02447 4307 4309 4305 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02446 4531 4307 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02445 4305 4308 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02444 6039 6434 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02443 6601 6919 6039 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02442 1514 2755 1420 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02441 1420 3586 1514 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02440 vss 2111 1420 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02439 1513 1514 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02438 982 3408 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02437 vss 2770 982 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02436 982 1189 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02435 vss 1188 982 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02434 4623 4744 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02433 4622 4745 4623 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02432 1629 1630 1882 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02431 vss 1893 1629 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02430 1631 1641 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02429 1882 1628 1631 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02428 vss 1641 1630 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02427 1628 1893 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02426 vss 2852 2703 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02425 2703 5893 2853 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02424 vss 5893 2856 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02423 2853 2856 2702 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02422 2851 2853 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02421 2702 6727 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02420 vss 3460 3461 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02419 3461 5893 3462 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02418 vss 5893 3464 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02417 3462 3464 3463 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02416 3459 3462 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02415 3463 6265 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02414 vss 4299 4301 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02413 4301 5893 4302 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02412 vss 5893 4304 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02411 4302 4304 4303 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02410 4300 4302 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02409 4303 5902 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02408 689 690 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02407 1372 857 689 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02406 vss 4068 3929 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02405 3929 4273 4069 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02404 4503 4069 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02403 3823 5773 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02402 3821 6440 3823 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02401 3510 5992 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02400 3625 6440 3510 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02399 5657 5762 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02398 6024 6748 5657 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02397 4381 4512 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02396 4521 6690 4381 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02395 5017 6876 5018 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02394 5018 6877 5017 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02393 vss 5524 5018 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02392 vss 3178 1663 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02391 1663 2325 1664 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02390 1662 1664 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02389 4268 5773 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02388 4505 4491 4268 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02387 4267 5992 4505 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02386 vss 4726 4267 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02385 4267 4265 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02384 5746 5805 5519 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02383 5519 5756 5746 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02382 vss 6905 5519 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02381 3716 3715 3718 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02380 3718 3967 3719 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02379 vss 4838 3716 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02378 3714 3719 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02377 3729 3728 3731 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02376 3731 4181 3730 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02375 vss 4399 3729 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02374 3727 3730 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02373 5438 5436 5437 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02372 5437 5440 5439 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02371 vss 5442 5438 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02370 5680 5439 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02369 6516 6820 6515 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02368 6515 6839 6623 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02367 vss 6850 6516 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02366 6622 6623 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02365 vss 918 979 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02364 vss 2537 979 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02363 979 919 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02362 1534 979 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02361 vss 5363 1788 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02360 1788 4299 1787 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02359 2407 1787 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02358 1677 1688 1678 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02357 1678 3593 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02356 1675 2347 1677 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02355 1676 1679 1675 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02354 3725 6190 3726 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02353 3726 6191 3725 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02352 vss 3969 3726 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02351 4599 5068 4600 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02350 4600 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02349 4598 5069 4599 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02348 4895 4693 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02347 4693 5372 4598 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02346 306 302 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02345 vss 312 306 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02344 306 305 953 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02343 953 2498 306 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02342 vss 2752 2754 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02341 vss 2750 2754 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02340 2754 2749 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02339 6173 2754 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02338 3738 2799 2673 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02337 2673 4051 3738 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02336 vss 2790 2673 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02335 5326 5112 4807 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02334 4807 5113 5326 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02333 vss 4935 4807 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02332 5719 6876 5603 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02331 5603 6877 5719 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02330 vss 6591 5603 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02329 5952 5719 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02328 vss 1368 1735 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02327 1368 1367 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02326 1735 1565 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02325 5794 5802 5796 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02324 5630 5803 5794 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02323 6682 5794 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02322 vss 5794 6682 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02321 5633 5801 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02320 vss 5800 5801 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02319 5802 5803 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02318 vss 6984 5803 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02317 5631 5797 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02316 5796 6976 5631 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02315 5797 5803 5633 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02314 5632 5802 5797 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02313 vss 5796 5632 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02312 vss 6682 5629 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02311 5629 6976 5630 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02310 3524 5773 3523 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02309 3523 4491 3638 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02308 vss 4275 3524 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02307 4083 3638 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02306 1347 1346 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02305 vss 2778 1347 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02304 1347 2766 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02303 vss 1345 1347 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02302 2553 1347 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02301 93 91 212 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02300 vss 787 93 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02299 94 216 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02298 212 92 94 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02297 vss 216 91 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02296 92 787 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02295 1465 2406 1464 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02294 1464 2412 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02293 1579 5359 1465 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02292 1956 1963 1957 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02291 1820 1964 1956 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02290 4241 1956 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02289 vss 1956 4241 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02288 1824 1962 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02287 vss 1959 1962 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02286 1963 1964 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02285 vss 3259 1964 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02284 1822 1960 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02283 1957 6976 1822 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02282 1960 1964 1824 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02281 1823 1963 1960 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02280 vss 1957 1823 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02279 vss 4241 1821 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02278 1821 6976 1820 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02277 vss 4205 3089 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02276 3089 3740 3185 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02275 3187 3185 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02274 2267 2406 2268 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02273 2268 2407 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02272 3062 3836 2267 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02271 3061 4509 3063 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02270 3063 3062 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02269 4523 3060 3061 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02268 1933 1194 1087 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02267 1087 1190 1933 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02266 vss 1191 1087 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02265 6415 6637 6416 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02264 6416 6675 6415 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02263 vss 6413 6416 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02262 6414 6415 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02261 6035 6142 6133 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02260 vss 6165 6035 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02259 6135 6137 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02258 vss 6135 6036 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02257 6133 6141 6135 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02256 6165 6133 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02255 vss 6133 6165 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02254 6036 6141 6137 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02253 6137 6142 6037 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02252 vss 6832 6142 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02251 6141 6142 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02250 vss 6139 6140 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02249 6037 6140 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02248 417 471 470 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02247 vss 1508 417 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02246 418 1652 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02245 470 468 418 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02244 vss 1652 471 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02243 468 1508 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02242 641 986 439 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02241 439 987 641 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02240 vss 504 439 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02239 4319 4425 4418 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02238 vss 5268 4319 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02237 4419 4421 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02236 vss 4419 4320 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02235 4418 4424 4419 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02234 5268 4418 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02233 vss 4418 5268 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02232 4320 4424 4421 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02231 4421 4425 4321 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02230 vss 5054 4425 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02229 4424 4425 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02228 vss 4589 4423 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02227 4321 4423 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02226 46 124 121 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02225 vss 525 46 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02224 47 48 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02223 vss 47 49 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02222 121 50 47 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02221 525 121 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02220 vss 121 525 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02219 49 50 48 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02218 48 124 122 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02217 vss 3259 124 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02216 50 124 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02215 vss 255 123 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02214 122 123 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02213 2170 4524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02212 vss 4094 2170 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02211 5644 6165 5643 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02210 5643 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02209 5642 5992 5644 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02208 5730 5731 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02207 5731 6440 5642 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02206 5875 6522 5878 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02205 5878 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02204 5876 5992 5875 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02203 5971 5970 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02202 5970 6440 5876 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02201 vss 5525 5523 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02200 5523 5983 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02199 vss 5521 5523 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02198 vss 4708 5880 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02197 5880 4466 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02196 vss 6224 5880 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02195 760 2194 762 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02194 762 857 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02193 761 1953 760 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02192 1029 852 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02191 852 3836 761 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02190 927 1218 928 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02189 928 1732 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02188 926 4239 927 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02187 1169 1013 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02186 1013 4748 926 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02185 3576 3582 3578 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02184 3484 3583 3576 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02183 3759 3576 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02182 vss 3576 3759 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02181 3487 3581 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02180 vss 3758 3581 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02179 3582 3583 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02178 vss 5054 3583 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02177 3485 3579 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02176 3578 6976 3485 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02175 3579 3583 3487 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02174 3486 3582 3579 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02173 vss 3578 3486 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02172 vss 3759 3483 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02171 3483 6976 3484 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02170 26 99 95 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02169 vss 633 26 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02168 27 29 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02167 vss 27 28 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02166 95 30 27 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02165 633 95 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02164 vss 95 633 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02163 28 30 29 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02162 29 99 97 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02161 vss 3160 99 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02160 30 99 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02159 vss 222 96 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02158 97 96 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02157 4587 4673 4318 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02156 4318 4671 4587 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02155 vss 5927 4318 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02154 6123 6876 6030 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02153 6030 6877 6123 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02152 vss 6807 6030 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02151 vss 6876 6213 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02150 6213 6877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02149 6421 6213 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02148 vss 5748 2829 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02147 2829 3049 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02146 2827 2829 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02145 204 319 148 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02144 148 320 204 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02143 vss 328 148 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02142 310 204 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02141 4927 5753 4707 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02140 4707 5767 4927 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02139 vss 5670 4707 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02138 57 3229 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02137 264 4501 57 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02136 1647 3391 1648 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02135 1648 2326 1647 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02134 vss 2111 1648 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02133 4825 5788 4826 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02132 4826 5570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02131 4954 5144 4825 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02130 5568 5788 5571 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02129 5571 5570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02128 5569 5575 5568 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02127 5229 5788 5230 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02126 5230 5570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02125 5556 5992 5229 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02124 2139 2146 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02123 vss 2052 2139 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02122 2139 2051 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02121 vss 2050 2139 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02120 vss 4699 4608 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02119 4608 4921 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02118 vss 4916 4608 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02117 2657 5959 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02116 2747 3186 2657 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02115 vss 3191 2747 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02114 2165 986 451 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02113 451 987 2165 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02112 vss 527 451 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02111 6513 6620 6619 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02110 vss 6740 6513 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02109 6514 6622 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02108 6619 6618 6514 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02107 vss 6622 6620 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02106 6618 6740 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02105 6660 6889 6537 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02104 6537 6661 6660 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02103 vss 6867 6537 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02102 6368 6806 6369 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02101 6369 6631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02100 6627 6820 6368 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02099 2591 2599 2593 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02098 2589 2598 2591 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02097 4235 2591 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02096 vss 2591 4235 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02095 2596 2597 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02094 vss 2601 2597 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02093 2599 2598 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02092 vss 3259 2598 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02091 2592 2594 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02090 2593 6976 2592 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02089 2594 2598 2596 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02088 2595 2599 2594 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02087 vss 2593 2595 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02086 vss 4235 2590 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02085 2590 6976 2589 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02084 5563 5788 5565 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02083 5565 5570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02082 5564 5773 5563 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02081 5138 5140 5139 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02080 5139 5141 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02079 5348 5349 5138 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02078 2260 2406 2261 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02077 2261 2412 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02076 2259 5359 2260 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02075 3234 4748 2259 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02074 2478 2487 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02073 2479 2734 2478 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02072 2488 2487 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02071 2485 2730 2488 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02070 4402 6791 4353 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02069 4352 4401 4402 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02068 4353 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02067 4399 4402 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02066 vss 6637 4352 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02065 4352 4653 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02064 6520 6806 6521 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02063 6521 6631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02062 6842 6850 6520 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02061 597 1652 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02060 596 1505 597 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02059 3515 3831 3514 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02058 3514 3629 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02057 3513 4253 3515 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02056 4212 3827 3513 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02055 5626 6952 5625 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02054 5625 6714 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02053 5787 6963 5626 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02052 1836 1989 1835 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02051 1835 1988 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02050 2196 1990 1836 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02049 6052 6636 6053 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02048 6053 6170 6171 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02047 vss 6372 6052 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02046 6169 6171 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02045 5607 6423 5606 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02044 5606 6374 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02043 5605 6375 5607 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02042 5973 6571 5605 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02041 vss 6440 5627 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02040 5627 5907 5790 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02039 5789 5790 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02038 300 581 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02037 vss 1169 300 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02036 300 301 579 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02035 579 461 300 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02034 5947 2498 1076 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02033 1076 1649 5947 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02032 vss 1172 1076 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02031 624 986 440 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02030 440 987 624 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02029 vss 500 440 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02028 3050 4941 3048 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02027 3048 4942 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02026 3049 5349 3050 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02025 2632 5157 2633 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02024 vss 4299 2634 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02023 2633 2634 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02022 6351 6791 6350 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02021 6349 6348 6351 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02020 6350 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02019 6347 6351 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02018 vss 6637 6349 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02017 6349 6613 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02016 4207 6220 4206 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02015 4206 5300 4207 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02014 vss 4205 4206 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02013 4892 4207 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02012 5336 5116 4816 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02011 4816 5125 5336 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02010 vss 4945 4816 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02009 2255 2396 2256 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02008 2256 2827 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02007 2254 2607 2255 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02006 4946 2397 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02005 2397 2506 2254 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02004 1940 2050 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02003 vss 2146 1940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02002 1940 2052 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02001 vss 2051 1940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02000 4671 1940 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01999 1935 2553 1811 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01998 1811 2356 1935 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01997 vss 2514 1811 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01996 2051 1935 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01995 vss 1188 1187 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01994 vss 2770 1187 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01993 1187 1189 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01992 1340 1187 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01991 vss 3263 866 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01990 866 3460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01989 1234 866 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01988 vss 3064 4286 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01987 3064 5363 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01986 4286 3263 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01985 vss 2533 2536 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01984 2533 2534 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01983 2536 2535 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01982 4849 4847 4761 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01981 4761 4850 4849 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01980 vss 6867 4761 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01979 4372 5773 4374 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01978 4374 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01977 4373 4748 4372 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01976 4499 4500 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01975 4500 6440 4373 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01974 vss 3197 3092 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01973 3092 3202 3194 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01972 3193 3194 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01971 1487 1888 1405 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01970 1405 2304 1487 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01969 vss 1884 1405 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01968 1485 1487 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01967 4755 4834 4847 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01966 vss 4836 4755 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01965 4756 5014 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01964 4847 4835 4756 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01963 vss 5014 4834 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01962 4835 4836 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01961 3511 3625 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01960 vss 3624 3511 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01959 3511 3821 5502 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01958 5502 3639 3511 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01957 vss 4299 3943 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01956 3943 5157 4092 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01955 4091 4092 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01954 vss 1760 1733 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01953 1733 1732 1734 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01952 2155 1734 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01951 vss 2387 137 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01950 137 138 136 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01949 1190 136 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01948 5576 5586 5577 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01947 vss 5575 5576 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01946 5578 5581 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01945 vss 5578 5579 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01944 5577 5583 5578 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01943 5575 5577 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01942 vss 5577 5575 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01941 5579 5583 5581 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01940 5581 5586 5582 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01939 vss 6984 5586 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01938 5583 5586 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01937 vss 5580 5584 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01936 5582 5584 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01935 4344 4533 4525 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01934 vss 4524 4344 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01933 4527 4530 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01932 vss 4527 4345 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01931 4525 4534 4527 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01930 4524 4525 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01929 vss 4525 4524 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01928 4345 4534 4530 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01927 4530 4533 4346 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01926 vss 6984 4533 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01925 4534 4533 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01924 vss 4531 4532 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01923 4346 4532 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01922 vss 6247 6250 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01921 6250 6475 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01920 vss 6245 6250 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01919 1072 1166 1694 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01918 vss 1165 1072 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01917 1073 1304 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01916 1694 1167 1073 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01915 vss 1304 1166 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01914 1167 1165 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01913 629 1194 437 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01912 437 1190 629 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01911 vss 636 437 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01910 74 772 75 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01909 75 86 73 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01908 vss 1151 74 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01907 320 73 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01906 4801 4927 4802 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01905 4802 4929 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01904 4800 5518 4801 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01903 5106 4930 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01902 4930 4928 4800 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01901 3207 3413 3098 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01900 3098 3414 3207 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01899 vss 5262 3098 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01898 3212 3207 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01897 3915 5992 3914 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01896 3914 5877 4037 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01895 vss 6440 3915 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01894 4038 4037 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01893 4796 5749 4795 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01892 4795 5748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01891 4794 6591 4796 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01890 4921 4923 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01889 4923 6440 4794 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01888 1091 1953 1092 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01887 1092 2194 1207 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01886 vss 3836 1091 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01885 2124 1207 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01884 3432 3430 3431 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01883 3431 5759 3433 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01882 vss 3789 3432 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01881 3429 3433 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01880 2224 2317 2499 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01879 vss 2319 2224 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01878 2225 2320 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01877 2499 2318 2225 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01876 vss 2320 2317 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01875 2318 2319 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01874 2056 2356 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01873 2600 2155 2056 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01872 2055 2156 2600 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01871 vss 4673 2055 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01870 2055 4671 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01869 2992 3413 2991 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01868 2991 3414 2992 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01867 vss 5272 2991 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01866 2990 2992 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01865 5520 5986 5522 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01864 5522 6214 5520 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01863 vss 6850 5522 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01862 5521 5520 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01861 5910 6665 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01860 6886 6885 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01859 4028 3421 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01858 3641 4239 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01857 5244 5670 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01856 6861 6874 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01855 2061 5069 2062 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01854 2062 2807 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01853 2060 2583 2061 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01852 2381 2166 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01851 2166 5992 2060 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01850 1399 3866 1400 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01849 1400 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01848 1398 3849 1399 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01847 1975 1397 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01846 1397 3664 1398 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01845 6061 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01844 6184 6431 6061 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01843 6060 6187 6184 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01842 vss 6182 6060 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01841 6060 6183 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01840 452 537 530 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01839 vss 3434 452 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01838 531 534 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01837 vss 531 454 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01836 530 536 531 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01835 3434 530 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01834 vss 530 3434 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01833 454 536 534 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01832 534 537 453 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01831 vss 3259 537 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01830 536 537 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01829 vss 677 535 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01828 453 535 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01827 vss 6420 6637 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01826 6637 6222 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01825 vss 6422 6637 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01824 vss 5789 5549 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01823 5549 5548 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01822 vss 6004 5549 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01821 637 1194 638 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01820 638 1190 637 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01819 vss 636 638 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01818 1188 637 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01817 4928 5112 4240 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01816 4240 5113 4928 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01815 vss 4239 4240 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01814 1776 3866 1777 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01813 1777 1778 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01812 1775 3849 1776 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01811 3229 1774 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01810 1774 3664 1775 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01809 6903 6906 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01808 4059 3434 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01807 6310 6905 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01806 4043 3802 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01805 3140 3451 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01804 3653 5992 3140 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01803 3864 4091 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01802 3863 4286 3864 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01801 vss 4686 4883 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01800 4686 4685 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01799 4883 4692 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01798 5190 5270 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01797 5468 5474 5190 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01796 5908 5907 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01795 6015 6025 5908 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01794 3246 4524 3116 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01793 3116 4273 3246 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01792 vss 4937 3116 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01791 6879 6876 6878 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01790 6878 6877 6879 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01789 vss 6874 6878 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01788 6875 6879 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01787 3132 3184 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01786 6191 3183 3132 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01785 2656 3182 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01784 2793 3174 2656 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01783 vss 6410 6411 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01782 6411 6414 6412 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01781 6418 6412 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01780 5969 5967 5968 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01779 5968 5993 5969 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01778 vss 5965 5968 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01777 vss 6690 5222 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01776 5222 5331 5330 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01775 5329 5330 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01774 3518 5069 3519 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01773 3519 4062 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01772 3517 3658 3518 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01771 4489 5363 3517 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01770 632 3195 631 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01769 631 981 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01768 630 641 632 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01767 975 629 630 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01766 625 1194 436 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01765 436 1190 625 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01764 vss 633 436 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01763 2472 2473 2507 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01762 vss 2712 2472 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01761 2471 2913 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01760 2507 2470 2471 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01759 vss 2913 2473 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01758 2470 2712 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01757 2315 3740 2223 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01756 2223 2520 2315 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01755 vss 2314 2223 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01754 2487 2315 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01753 4886 5954 4777 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01752 4777 5502 4886 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01751 vss 5959 4777 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01750 3139 3853 3138 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01749 3138 3856 3249 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01748 vss 4275 3139 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01747 3248 3249 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01746 4822 4952 4823 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01745 4823 4953 4951 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01744 vss 5154 4822 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01743 5140 4951 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01742 2654 3182 2655 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01741 2655 2779 2745 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01740 vss 3174 2654 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01739 2744 2745 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01738 vss 1789 1991 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01737 1789 2852 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01736 1991 3460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01735 1574 1989 1456 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01734 1456 1745 1574 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01733 vss 1572 1456 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01732 2396 1574 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01731 vss 2534 1717 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01730 1717 2350 1718 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01729 1716 1718 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01728 2948 5953 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01727 2947 3186 2948 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01726 vss 2952 2947 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01725 2946 2947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01724 1503 3391 1417 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01723 1417 2326 1503 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01722 vss 2111 1417 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01721 1501 1503 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01720 vss 3422 4466 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01719 3422 4524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01718 4466 3607 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01717 87 84 86 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01716 vss 615 87 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01715 88 216 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01714 86 85 88 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01713 vss 216 84 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01712 85 615 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01711 1752 3866 1753 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01710 1753 4286 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01709 1750 2406 1752 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01708 1749 1751 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01707 1751 3836 1750 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01706 vss 1559 1443 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01705 1443 1968 1556 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01704 1703 1556 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01703 vss 2520 2523 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01702 2523 2521 2524 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01701 2522 2524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01700 6323 6331 6322 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01699 vss 6522 6323 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01698 6324 6327 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01697 vss 6324 6325 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01696 6322 6330 6324 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01695 6522 6322 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01694 vss 6322 6522 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01693 6325 6330 6327 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01692 6327 6331 6329 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01691 vss 6832 6331 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01690 6330 6331 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01689 vss 6326 6328 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01688 6329 6328 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01687 vss 5363 3055 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01686 3055 3263 3056 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01685 4942 3056 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01684 1280 1480 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01683 vss 1478 1280 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01682 4474 4472 4331 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01681 4331 5125 4474 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01680 vss 4471 4331 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01679 4952 4474 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01678 2540 2773 2539 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01677 2538 5958 2540 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01676 2539 4205 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01675 2537 2540 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01674 vss 3199 2538 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01673 2538 3618 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01672 2715 2915 2638 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01671 2638 2716 2715 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01670 vss 2717 2638 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01669 2712 2715 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01668 3137 4258 3136 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01667 3136 3231 3228 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01666 vss 3438 3137 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01665 3227 3228 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01664 vss 3664 3534 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01663 3534 3866 3656 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01662 3853 3656 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01661 1104 1218 1105 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01660 1105 1732 1219 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01659 vss 4748 1104 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01658 1564 1219 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01657 1710 2349 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01656 1709 2553 1710 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01655 vss 1716 1709 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01654 1708 1709 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01653 341 349 342 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01652 vss 1182 341 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01651 343 345 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01650 vss 343 344 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01649 342 348 343 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01648 1182 342 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01647 vss 342 1182 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01646 344 348 345 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01645 345 349 346 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01644 vss 3160 349 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01643 348 349 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01642 vss 350 347 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01641 346 347 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01640 6038 6175 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01639 6326 6143 6038 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01638 4496 4497 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01637 vss 4499 4496 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01636 4496 4725 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01635 vss 4492 4496 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01634 5218 5523 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01633 5325 5324 5218 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01632 vss 5144 2192 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01631 2192 5359 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01630 2193 2192 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01629 56 405 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01628 133 4299 56 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01627 5186 5701 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01626 5453 5265 5186 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01625 6353 6356 6359 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01624 vss 6352 6353 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01623 6355 6622 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01622 6359 6354 6355 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01621 vss 6622 6356 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01620 6354 6352 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01619 6667 6668 6539 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01618 6539 6676 6667 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01617 vss 6867 6539 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01616 5030 6447 5031 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01615 5031 6600 5030 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01614 vss 6601 5031 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01613 5029 5030 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01612 vss 6422 5981 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01611 vss 6222 5981 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01610 5981 6420 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01609 6867 5981 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01608 4820 5133 4819 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01607 4819 5125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01606 5132 6447 4820 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01605 409 2727 408 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01604 408 579 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01603 573 1876 409 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01602 6392 6806 6391 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01601 6391 6631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01600 6390 6874 6392 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01599 5982 6906 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01598 vss 6420 5982 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01597 5982 6222 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01596 vss 6422 5982 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01595 6208 5982 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01594 4351 4849 4350 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01593 4350 4397 4398 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01592 vss 5025 4351 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01591 4396 4398 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01590 4330 4470 4329 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01589 4329 4469 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01588 4609 6951 4330 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01587 2994 4608 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01586 2993 2996 2994 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01585 4915 5805 4792 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01584 4792 5756 4915 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01583 vss 4914 4792 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01582 4916 4915 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01581 267 3460 173 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01580 173 1583 267 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01579 vss 264 173 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01578 265 267 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01577 2579 2578 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01576 2773 3438 2579 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01575 3721 3720 3722 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01574 3722 3734 3723 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01573 vss 4843 3721 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01572 3717 3723 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01571 6406 6806 6407 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01570 6407 6631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01569 6405 6885 6406 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01568 6663 6876 6538 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01567 6538 6877 6663 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01566 vss 6885 6538 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01565 6661 6663 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01564 4799 5552 4798 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01563 4798 5329 4926 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01562 vss 5116 4799 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01561 6600 4926 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01560 484 2506 424 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01559 425 489 484 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01558 424 1737 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01557 482 484 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01556 vss 491 425 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01555 425 486 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01554 vss 3592 3407 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01553 3407 3404 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01552 3408 3407 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01551 5071 5068 5073 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01550 5073 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01549 5072 5069 5071 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01548 5496 5070 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01547 5070 6265 5072 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01546 4026 4275 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01545 vss 4024 4026 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01544 4026 4708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01543 vss 6224 4026 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01542 4469 4026 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01541 vss 3836 1830 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01540 1830 2406 1978 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01539 2182 1978 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01538 6345 6791 6344 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01537 6343 6609 6345 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01536 6344 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01535 6342 6345 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01534 vss 6637 6343 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01533 6343 6607 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01532 4157 6876 4156 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01531 4156 6877 4157 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01530 vss 5026 4156 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01529 vss 6262 6466 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01528 6262 6261 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01527 6466 6263 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01526 6953 6957 6955 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01525 6955 6959 6954 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01524 vss 6952 6953 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01523 6968 6954 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01522 5277 4895 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01521 vss 4896 5277 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01520 1719 1904 1720 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01519 1720 1737 1721 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01518 vss 2375 1719 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01517 1722 1721 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01516 755 3217 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01515 784 1904 755 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01514 754 2747 784 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01513 vss 4176 754 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01512 754 1322 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01511 3827 4250 3826 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01510 3826 4491 3827 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01509 vss 5349 3826 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01508 vss 3416 3099 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01507 3099 4014 3209 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01506 3208 3209 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01505 5881 5886 5991 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01504 vss 5992 5881 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01503 5882 5884 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01502 vss 5882 5883 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01501 5991 5885 5882 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01500 5992 5991 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01499 vss 5991 5992 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01498 5883 5885 5884 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01497 5884 5886 5995 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01496 vss 6984 5886 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01495 5885 5886 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01494 vss 5994 5996 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01493 5995 5996 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01492 1301 1305 4880 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01491 vss 1300 1301 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01490 1303 1304 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01489 4880 1302 1303 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01488 vss 1304 1305 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01487 1302 1300 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01486 325 323 324 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01485 324 611 326 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01484 vss 332 325 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01483 322 326 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01482 vss 6440 3919 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01481 3919 5773 4063 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01480 4062 4063 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01479 2631 2629 2630 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01478 2630 2632 2631 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01477 vss 4280 2630 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01476 2628 2631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01475 6360 6359 6361 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01474 6361 6624 6360 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01473 vss 6867 6361 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01472 4635 4640 4749 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01471 vss 4748 4635 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01470 4636 4638 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01469 vss 4636 4637 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01468 4749 4639 4636 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01467 4748 4749 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01466 vss 4749 4748 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01465 4637 4639 4638 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01464 4638 4640 4750 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01463 vss 6984 4640 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01462 4639 4640 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01461 vss 4751 4752 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01460 4750 4752 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01459 1055 4094 1054 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01458 1054 2352 1056 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01457 vss 3664 1055 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01456 2615 1056 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01455 1711 2371 1712 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01454 1712 2506 1713 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01453 vss 2782 1711 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01452 1904 1713 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01451 4804 4941 4803 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01450 4803 4942 4931 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01449 vss 5992 4804 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01448 5805 4931 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01447 5483 5954 5482 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01446 5482 5502 5483 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01445 vss 5958 5482 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01444 5176 6919 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01443 5259 6434 5176 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01442 5175 6867 5259 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01441 vss 6115 5175 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01440 5175 5254 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01439 6949 6963 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01438 6950 6959 6949 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01437 vss 6948 6950 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01436 6946 6950 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01435 5516 5805 5515 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01434 5515 5756 5516 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01433 vss 5524 5515 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01432 5733 5516 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01431 2377 2799 2245 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01430 2245 4051 2377 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01429 vss 2384 2245 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01428 2501 2377 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01427 6224 5773 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01426 4282 5575 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01425 6581 6807 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01424 2481 2486 2483 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01423 vss 2734 2481 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01422 2484 2487 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01421 2483 2482 2484 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01420 vss 2487 2486 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01419 2482 2734 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01418 5512 5749 5514 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01417 5514 5748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01416 5513 6874 5512 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01415 5510 5511 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01414 5511 6440 5513 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01413 5464 5473 5465 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01412 vss 6591 5464 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01411 5466 5469 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01410 vss 5466 5467 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01409 5465 5471 5466 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01408 6591 5465 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01407 vss 5465 6591 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01406 5467 5471 5469 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01405 5469 5473 5470 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01404 vss 6832 5473 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01403 5471 5473 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01402 vss 5468 5472 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01401 5470 5472 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01400 5894 6243 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01399 6473 6242 5894 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01398 vss 2358 2361 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01397 2358 2356 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01396 2361 2553 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01395 393 986 394 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01394 394 987 393 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01393 vss 392 394 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01392 1345 393 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01391 1526 1918 1427 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01390 1427 1919 1526 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01389 vss 2521 1427 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01388 1524 1526 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01387 3861 4088 3860 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01386 3860 4091 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01385 3862 4089 3861 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01384 5877 3859 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01383 3859 4087 3862 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01382 5567 6682 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01381 3634 5359 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01380 4280 5144 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01379 3037 4235 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01378 1576 4937 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01377 3040 4935 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01376 vss 5315 5305 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01375 5305 5971 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01374 vss 5312 5305 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01373 5595 5697 5695 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01372 vss 6591 5595 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01371 5596 6616 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01370 5695 5694 5596 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01369 vss 6616 5697 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01368 5694 6591 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01367 5639 5708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01366 6160 6166 5639 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01365 6541 6893 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01364 vss 6893 6670 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01363 vss 6906 6540 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01362 6671 6669 6541 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01361 6540 6670 6671 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01360 6668 6671 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01359 vss 6671 6668 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01358 6669 6906 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01357 4669 6806 4670 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01356 4670 6910 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01355 4668 4918 4669 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01354 4827 5361 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01353 4961 4953 4827 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01352 801 3210 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01351 vss 2537 801 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01350 801 919 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01349 vss 918 801 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01348 3370 4942 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01347 3369 3658 3370 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01346 4261 5992 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01345 539 2194 458 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01344 458 2195 539 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01343 vss 6440 458 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01342 1732 539 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01341 5865 6628 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01340 6150 5864 5865 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01339 3351 5069 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01338 3624 3818 3351 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01337 4018 4213 3912 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01336 3912 4212 4018 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01335 vss 5299 3912 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01334 1285 1641 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01333 1482 1893 1285 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01332 2127 2124 2126 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01331 2123 2122 2127 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01330 2126 2125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01329 2526 2127 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01328 vss 2535 2123 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01327 2123 2737 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01326 6802 6792 6793 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01325 6793 6794 6802 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01324 vss 6867 6793 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01323 vss 1330 1325 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01322 1325 1328 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01321 5045 1325 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01320 6711 6714 6561 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01319 vss 6952 6712 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01318 6561 6712 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01317 2309 2319 2220 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01316 2220 2320 2309 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01315 vss 2485 2220 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01314 2308 2309 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01313 6849 6847 6848 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01312 6848 6851 6849 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01311 vss 6867 6848 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01310 6019 5905 5897 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01309 5896 5906 6019 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01308 6714 6019 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01307 vss 6019 6714 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01306 5901 5904 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01305 vss 5903 5904 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01304 5905 5906 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01303 vss 6984 5906 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01302 5898 5900 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01301 5897 6976 5898 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01300 5900 5906 5901 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01299 5899 5905 5900 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01298 vss 5897 5899 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01297 vss 6714 5895 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01296 5895 6976 5896 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01295 5170 5670 5171 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01294 5171 5914 5247 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01293 vss 6665 5170 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01292 6116 5247 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01291 5088 5045 4684 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01290 4684 5044 5088 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01289 vss 5964 4684 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01288 vss 200 141 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01287 141 322 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01286 571 189 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01285 141 191 189 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01284 189 2498 141 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01283 2912 2914 5723 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01282 vss 2909 2912 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01281 2911 2913 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01280 5723 2910 2911 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01279 vss 2913 2914 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01278 2910 2909 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01277 910 936 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01276 1877 1479 910 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01275 vss 5262 5060 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01274 5060 5309 5059 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01273 vss 5309 5061 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01272 5059 5061 5058 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01271 5057 5059 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01270 5058 5958 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01269 vss 5243 4197 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01268 4197 5309 4198 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01267 vss 5309 4199 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01266 4198 4199 4196 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01265 4434 4198 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01264 4196 5959 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01263 vss 4308 3903 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01262 3903 5309 4004 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01261 vss 5309 4005 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01260 4004 4005 3904 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01259 4002 4004 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01258 3904 5725 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01257 vss 5272 5192 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01256 5192 5309 5273 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01255 vss 5309 5276 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01254 5273 5276 5193 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01253 5715 5273 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01252 5193 5953 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01251 6068 6205 6067 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01250 6067 6667 6206 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01249 vss 6207 6068 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01248 6204 6206 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01247 2809 2815 2810 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01246 2687 2816 2809 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01245 4935 2809 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01244 vss 2809 4935 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01243 2690 2813 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01242 vss 2826 2813 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01241 2815 2816 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01240 vss 3259 2816 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01239 2688 2812 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01238 2810 6976 2688 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01237 2812 2816 2690 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01236 2689 2815 2812 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01235 vss 2810 2689 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01234 vss 4935 2686 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01233 2686 6976 2687 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01232 4812 4946 4811 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01231 4811 5549 4940 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01230 vss 4947 4812 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01229 4939 4940 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01228 6011 6714 6010 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01227 6010 6469 6011 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01226 vss 6442 6010 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01225 3847 4089 3848 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01224 3848 4287 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01223 3846 4286 3847 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01222 4708 3866 3846 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01221 2292 2298 2087 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01220 2087 2301 2292 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01219 vss 2086 2087 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01218 vss 766 413 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01217 413 571 463 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01216 461 463 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01215 vss 6711 6560 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01214 6560 6956 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01213 6707 6708 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01212 6560 6962 6708 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01211 6708 6715 6560 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01210 1098 3217 1099 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01209 1099 1212 1213 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01208 vss 1985 1098 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01207 1558 1213 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01206 1049 1234 1048 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01205 1048 1975 1050 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01204 vss 1233 1049 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01203 1380 1050 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01202 vss 2314 621 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01201 621 640 620 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01200 619 620 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01199 1129 4524 1128 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01198 1128 4094 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01197 1239 5363 1129 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01196 6824 6834 6825 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01195 vss 6850 6824 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01194 6826 6827 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01193 vss 6826 6828 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01192 6825 6833 6826 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01191 6850 6825 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01190 vss 6825 6850 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01189 6828 6833 6827 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01188 6827 6834 6829 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01187 vss 6832 6834 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01186 6833 6834 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01185 vss 6830 6831 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01184 6829 6831 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01183 4865 4855 4763 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01182 4763 4854 4865 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01181 vss 6867 4763 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01180 4148 4149 5004 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01179 vss 5670 4148 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01178 4147 5245 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01177 5004 4146 4147 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01176 vss 5245 4149 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01175 4146 5670 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01174 6692 6682 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01173 vss 6480 6692 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01172 583 946 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01171 581 586 583 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01170 582 2086 581 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01169 vss 588 582 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01168 582 774 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01167 606 608 607 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01166 vss 1317 606 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01165 609 619 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01164 607 605 609 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01163 vss 619 608 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01162 605 1317 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01161 153 772 154 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01160 154 212 213 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01159 vss 1151 153 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01158 486 213 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01157 vss 6187 2228 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01156 2228 3186 2328 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01155 2326 2328 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01154 vss 3595 3492 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01153 3492 4008 3594 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01152 3593 3594 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01151 6333 6341 6332 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01150 vss 6376 6333 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01149 6334 6338 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01148 vss 6334 6335 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01147 6332 6340 6334 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01146 6376 6332 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01145 vss 6332 6376 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01144 6335 6340 6338 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01143 6338 6341 6339 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01142 vss 6832 6341 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01141 6340 6341 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01140 vss 6336 6337 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01139 6339 6337 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01138 5124 6447 5123 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01137 5123 5125 5124 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01136 vss 5544 5123 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01135 5338 5124 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01134 vss 2531 2532 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01133 2531 2530 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01132 2532 3586 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01131 1523 1918 1426 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01130 1426 1919 1523 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01129 vss 2349 1426 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01128 1521 1523 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01127 5216 5320 5217 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01126 5217 5321 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01125 5215 5322 5216 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01124 5528 5323 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01123 5323 5319 5215 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01122 3934 4515 3935 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01121 3935 4506 4081 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01120 vss 4079 3934 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01119 4080 4081 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01118 5654 6212 5653 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01117 5653 5750 5747 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01116 vss 5746 5654 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01115 5745 5747 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01114 5967 2498 2500 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01113 2500 2499 5967 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01112 vss 2517 2500 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01111 6244 6974 6102 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01110 6102 6477 6244 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01109 vss 6714 6102 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01108 6245 6244 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01107 5322 5753 5213 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01106 5213 5767 5322 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01105 vss 6665 5213 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01104 2504 3217 2505 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01103 2505 2506 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01102 2502 2501 2504 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01101 2733 2503 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01100 2503 2782 2502 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01099 vss 5764 5766 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01098 5764 5763 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01097 5766 5998 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01096 4085 4083 3937 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01095 3937 4082 4085 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01094 vss 5902 3937 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01093 4518 4085 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01092 6433 6688 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01091 6685 6692 6433 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01090 vss 1333 1332 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01089 1332 1530 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01088 vss 1524 1332 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01087 3478 6423 3477 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01086 3477 3947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01085 3728 3560 3478 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01084 715 824 817 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01083 vss 1191 715 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01082 818 821 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01081 vss 818 716 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01080 817 823 818 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01079 1191 817 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01078 vss 817 1191 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01077 716 823 821 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01076 821 824 717 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01075 vss 3259 824 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01074 823 824 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01073 vss 990 822 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01072 717 822 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01071 4701 5753 4700 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01070 4700 5767 4701 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01069 vss 4918 4700 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01068 915 968 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01067 914 965 915 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01066 790 2746 708 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01065 708 1322 790 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01064 vss 3188 708 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01063 794 790 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01062 1217 1989 1101 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01061 1101 1745 1217 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01060 vss 1560 1101 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01059 1215 1217 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01058 1741 1967 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01057 1740 1758 1741 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01056 749 1737 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01055 946 2506 749 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01054 5668 6791 5635 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01053 5634 5915 5668 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01052 5635 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01051 5666 5668 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01050 vss 6637 5634 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01049 5634 6777 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01048 3381 6423 3380 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01047 3380 3947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01046 3556 3379 3381 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01045 5870 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01044 6843 6431 5870 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01043 5869 5958 6843 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01042 vss 6182 5869 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01041 5869 6183 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01040 vss 4082 3647 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01039 vss 3662 3647 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01038 3647 4083 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01037 3648 3647 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01036 vss 1564 1568 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01035 vss 1575 1568 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01034 1568 1565 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01033 2803 1568 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01032 5489 5954 5488 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01031 5488 5502 5489 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01030 vss 5963 5488 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01029 4327 5068 4328 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01028 4328 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01027 4455 5069 4327 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01026 4739 5133 4738 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01025 4738 4737 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01024 5343 5272 4739 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01023 2069 2399 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01022 2578 2400 2069 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01021 1541 986 719 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01020 719 987 1541 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01019 vss 829 719 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01018 5224 5773 5223 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01017 5223 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01016 5331 6440 5224 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01015 2608 2610 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01014 3413 2607 2608 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01013 1319 1679 1321 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01012 1321 1687 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01011 1320 3217 1319 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01010 6069 6806 6070 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01009 6070 6631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01008 6207 6893 6069 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01007 6178 5723 5604 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01006 5604 5721 6178 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01005 vss 5948 5604 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01004 2576 3818 2577 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01003 2577 5069 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01002 2575 5349 2576 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01001 2790 6440 2575 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01000 2247 3818 2248 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00999 2248 5069 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00998 2246 5349 2247 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00997 2384 6440 2246 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00996 2270 4941 2271 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00995 2271 4088 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00994 2625 3849 2270 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00993 744 857 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00992 859 3229 744 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00991 743 1982 859 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00990 vss 1965 743 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00989 742 1389 859 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00988 vss 3460 742 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00987 1685 1688 1686 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00986 1686 3593 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00985 1918 2347 1685 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00984 5479 5483 5480 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00983 5480 5478 5481 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00982 vss 5485 5479 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00981 5932 5481 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00980 vss 4889 4778 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00979 4778 4887 4888 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00978 5036 4888 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00977 3640 3641 3525 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00976 3525 3648 3640 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00975 vss 3645 3525 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00974 4747 4633 4627 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00973 4624 4634 4747 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00972 6242 4747 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00971 vss 4747 6242 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00970 4631 4632 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00969 vss 4630 4632 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00968 4633 4634 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00967 vss 6984 4634 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00966 4626 4629 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00965 4627 6976 4626 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00964 4629 4634 4631 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00963 4628 4633 4629 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00962 vss 4627 4628 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00961 vss 6242 4625 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00960 4625 6976 4624 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00959 6429 6434 6428 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00958 6428 6680 6427 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00957 vss 6919 6429 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00956 6426 6427 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00955 2227 2508 2226 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00954 2226 2742 2327 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00953 vss 2507 2227 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00952 2325 2327 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00951 431 624 432 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00950 432 3193 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00949 430 625 431 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00948 493 3217 430 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00947 1226 4748 1115 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00946 1114 1379 1226 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00945 1115 1576 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00944 1224 1226 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00943 vss 1746 1114 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00942 1114 1745 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00941 5505 5954 5503 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00940 5503 5502 5505 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00939 vss 5742 5503 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00938 vss 3865 3866 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00937 3865 5157 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00936 3866 4299 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00935 vss 5773 3450 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00934 3450 5349 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00933 3452 3450 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00932 2186 2182 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00931 2184 2183 2186 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00930 2185 2193 2184 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00929 vss 2180 2185 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00928 2181 2399 2184 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00927 vss 2799 2181 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00926 3887 6434 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00925 3964 6919 3887 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00924 3886 5372 3964 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00923 vss 4217 3886 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00922 3886 5502 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00921 2076 4299 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00920 2208 5363 2076 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00919 944 1289 945 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00918 945 1158 944 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00917 vss 946 945 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00916 943 944 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00915 4889 5954 4779 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00914 4779 5502 4889 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00913 vss 5725 4779 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00912 2699 2849 2842 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00911 vss 2852 2699 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00910 2844 2846 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00909 vss 2844 2700 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00908 2842 2850 2844 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00907 2852 2842 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00906 vss 2842 2852 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00905 2700 2850 2846 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00904 2846 2849 2701 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00903 vss 3259 2849 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00902 2850 2849 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00901 vss 2851 2848 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00900 2701 2848 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00899 6087 6952 6088 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00898 6088 6714 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00897 6086 6974 6087 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00896 6238 6239 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00895 6239 6963 6086 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00894 3785 3795 3784 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00893 3784 4604 3786 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00892 vss 4215 3785 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00891 3783 3786 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00890 76 81 78 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00889 78 328 77 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00888 vss 214 76 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00887 478 77 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00886 vss 2623 2621 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00885 2621 2622 2620 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00884 3457 2620 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00883 vss 2625 2626 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00882 2626 2628 2627 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00881 2833 2627 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00880 vss 2400 2258 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00879 2258 2399 2401 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00878 4213 2401 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00877 vss 2727 2644 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00876 2644 2728 2729 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00875 2924 2729 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00874 5621 5783 5775 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00873 vss 5773 5621 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00872 5777 5779 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00871 vss 5777 5622 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00870 5775 5782 5777 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00869 5773 5775 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00868 vss 5775 5773 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00867 5622 5782 5779 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00866 5779 5783 5623 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00865 vss 6984 5783 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00864 5782 5783 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00863 vss 5778 5781 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00862 5623 5781 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00861 3068 3076 3069 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00860 vss 3263 3068 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00859 3070 3073 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00858 vss 3070 3072 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00857 3069 3075 3070 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00856 3263 3069 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00855 vss 3069 3263 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00854 3072 3075 3073 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00853 3073 3076 3071 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00852 vss 3259 3076 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00851 3075 3076 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00850 vss 3262 3074 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00849 3071 3074 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00848 4925 5986 4797 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00847 4797 6214 4925 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00846 vss 6591 4797 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00845 415 467 1304 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00844 vss 571 415 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00843 414 466 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00842 1304 464 414 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00841 vss 466 467 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00840 464 571 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00839 5649 5749 5650 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00838 5650 5748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00837 5648 6850 5649 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00836 5738 5739 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00835 5739 6440 5648 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00834 5536 5755 5539 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00833 5539 5538 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00832 5537 5540 5536 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00831 5533 5535 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00830 5535 5534 5537 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00829 6348 6876 6346 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00828 6346 6877 6348 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00827 vss 6850 6346 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00826 vss 5495 5728 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00825 5495 5493 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00824 5728 5496 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00823 vss 4611 5127 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00822 5127 4612 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00821 vss 6422 5127 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00820 59 58 191 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00819 vss 607 59 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00818 61 592 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00817 191 60 61 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00816 vss 592 58 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00815 60 607 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00814 6430 6934 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00813 vss 6694 6430 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00812 5978 6173 5487 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00811 5487 6172 5978 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00810 vss 5964 5487 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00809 3482 4696 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00808 3572 3740 3482 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00807 3481 6727 3572 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00806 vss 3737 3481 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00805 3481 3738 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00804 2221 2312 2320 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00803 vss 2730 2221 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00802 2222 2487 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00801 2320 2311 2222 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00800 vss 2487 2312 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00799 2311 2730 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00798 3165 5044 3084 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00797 3084 5045 3165 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00796 vss 3969 3084 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00795 4824 4954 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00794 5151 4952 4824 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00793 5156 5569 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00792 5580 5154 5156 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00791 vss 4704 4610 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00790 4610 4609 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00789 vss 5094 4610 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00788 523 1194 449 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00787 449 1190 523 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00786 vss 522 449 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00785 1346 523 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00784 4071 5349 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00783 3836 4094 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00782 4275 4524 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00781 4501 4748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00780 2799 3263 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00779 3664 2852 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00778 4271 4276 4272 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00777 4272 4941 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00776 4270 4286 4271 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00775 5341 4269 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00774 4269 4275 4270 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00773 930 1991 931 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00772 931 2352 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00771 929 4094 930 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00770 1223 1043 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00769 1043 5363 929 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00768 1032 5749 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00767 1221 1031 1032 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00766 1030 1232 1221 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00765 vss 1029 1030 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00764 1028 1732 1221 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00763 vss 1231 1028 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00762 2054 2782 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00761 2057 2371 2054 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00760 2053 2154 2057 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00759 vss 4673 2053 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00758 2053 4671 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00757 6044 6164 6156 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00756 vss 6740 6044 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00755 6157 6158 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00754 vss 6157 6045 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00753 6156 6163 6157 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00752 6740 6156 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00751 vss 6156 6740 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00750 6045 6163 6158 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00749 6158 6164 6046 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00748 vss 6832 6164 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00747 6163 6164 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00746 vss 6160 6161 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00745 6046 6161 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00744 4460 6186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00743 vss 6220 4460 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00742 4460 4456 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00741 vss 4477 4460 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00740 4042 5987 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00739 vss 6188 4042 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00738 4042 4038 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00737 vss 4212 4042 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00736 5558 5556 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00735 5994 5557 5558 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00734 5562 5564 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00733 5778 5561 5562 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00732 5231 5348 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00731 5354 5788 5231 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00730 3795 3792 3794 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00729 3794 3793 3795 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00728 vss 3790 3794 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00727 2269 2408 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00726 3455 2409 2269 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00725 2698 2836 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00724 3449 2837 2698 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00723 863 3460 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00722 6469 6440 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00721 6476 6714 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00720 6921 6974 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00719 vss 2609 2610 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00718 2609 5893 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00717 2610 3051 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00716 5598 5707 5951 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00715 vss 5705 5598 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00714 5599 6616 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00713 5951 5704 5599 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00712 vss 6616 5707 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00711 5704 5705 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00710 6358 6357 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00709 6830 6841 6358 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00708 6017 6015 6016 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00707 6018 6694 6017 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00706 6016 6263 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00705 6256 6017 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00704 vss 6013 6018 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00703 6018 6014 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00702 6432 6682 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00701 vss 6694 6432 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00700 6432 6480 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00699 vss 6934 6432 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00698 6431 6432 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00697 5028 6806 5027 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00696 5027 6910 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00695 5025 5026 5028 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00694 3502 4226 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00693 3614 3613 3502 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00692 4020 4881 3489 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00691 3489 4880 4020 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00690 vss 5964 3489 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00689 4705 5753 4706 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00688 4706 5767 4705 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00687 vss 5026 4706 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00686 4704 4705 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00685 199 592 145 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00684 145 607 199 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00683 vss 603 145 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00682 196 199 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00681 3828 5992 3829 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00680 3829 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00679 4258 6440 3828 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00678 3440 5773 3439 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00677 3439 4726 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00676 3629 6440 3440 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00675 2624 2622 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00674 2836 2623 2624 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00673 1542 1194 997 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00672 997 1190 1542 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00671 vss 1002 997 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00670 6072 6208 6071 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00669 6071 6424 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00668 6209 6211 6072 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00667 1093 2139 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00666 1208 2138 1093 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00665 vss 2946 2324 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00664 2324 2950 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00663 2356 2324 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00662 3832 5773 3830 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00661 3830 4265 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00660 3831 6440 3832 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00659 6565 6714 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00658 6715 6952 6565 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00657 2125 4748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00656 vss 4524 2125 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00655 1022 1231 1021 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00654 1021 1218 1022 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00653 vss 1732 1021 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00652 1946 1022 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00651 1121 1582 1122 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00650 1122 1236 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00649 1232 2625 1121 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00648 5508 5805 5509 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00647 5509 5756 5508 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00646 vss 5670 5509 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00645 vss 6265 5201 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00644 5201 5309 5293 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00643 vss 5309 5296 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00642 5293 5296 5200 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00641 5292 5293 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00640 5200 5804 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00639 vss 5902 4202 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00638 4202 5309 4203 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00637 vss 5309 4204 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00636 4203 4204 4201 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00635 4200 4203 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00634 4201 5963 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00633 vss 5372 4193 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00632 4193 5309 4192 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00631 vss 5309 4195 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00630 4192 4195 4194 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00629 4191 4192 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00628 4194 6187 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00627 4380 6690 4379 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00626 4379 6011 4511 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00625 vss 4509 4380 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00624 4510 4511 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00623 207 1900 150 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00622 149 328 207 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00621 150 2161 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00620 480 207 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00619 vss 319 149 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00618 149 320 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00617 1079 1176 1078 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00616 1078 1175 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00615 1177 2331 1079 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00614 1175 2746 1077 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00613 1077 1322 1175 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00612 vss 3188 1077 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00611 5226 5341 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00610 5346 5349 5226 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00609 3920 4726 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00608 4254 5773 3920 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00607 1715 2371 1714 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00606 1714 2506 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00605 1727 2782 1715 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00604 1440 2194 1441 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00603 1441 1553 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00602 1439 1953 1440 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00601 2117 3836 1439 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00600 3879 3951 3880 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00599 3880 4171 3952 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00598 vss 5666 3879 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00597 3950 3952 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00596 3475 3556 3474 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00595 3474 3766 3557 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00594 vss 3957 3475 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00593 3555 3557 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00592 vss 6727 5207 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00591 5207 5309 5308 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00590 vss 5309 5310 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00589 5308 5310 5208 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00588 5306 5308 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00587 5208 5742 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00586 6588 6190 5923 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00585 5923 6191 6588 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00584 vss 5927 5923 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00583 4741 5349 4740 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00582 4740 5877 4742 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00581 vss 6440 4741 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00580 5548 4742 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00579 1061 1150 2913 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00578 vss 1280 1061 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00577 1062 1151 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00576 2913 1149 1062 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00575 vss 1151 1150 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00574 1149 1280 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00573 3925 4276 3926 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00572 3926 4941 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00571 3924 4286 3925 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00570 6221 4275 3924 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00569 4279 4276 4278 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00568 4278 4941 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00567 4277 4286 4279 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00566 4281 4275 4277 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00565 2238 2512 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00564 2353 2534 2238 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00563 2237 2521 2353 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00562 vss 2350 2237 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00561 2236 2349 2353 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00560 vss 2520 2236 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00559 1016 1218 1015 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00558 1015 1732 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00557 1014 4239 1016 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00556 1876 4748 1014 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00555 1095 1953 1096 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00554 1096 2194 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00553 1094 4239 1095 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00552 1209 3836 1094 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00551 vss 4094 3945 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00550 3945 5893 4097 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00549 vss 5893 4098 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00548 4097 4098 3944 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00547 4093 4097 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00546 3944 5272 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00545 1696 1925 1698 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00544 1698 1695 1697 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00543 vss 1694 1696 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00542 1944 1697 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00541 vss 2314 339 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00540 339 494 340 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00539 488 340 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00538 4259 4258 4260 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00537 4260 5551 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00536 4256 4253 4259 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00535 4257 4255 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00534 4255 4254 4256 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00533 vss 2138 2141 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00532 2141 2139 2140 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00531 2981 2140 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00530 5314 5805 5209 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00529 5209 5756 5314 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00528 vss 6665 5209 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00527 5312 5314 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00526 5427 5435 5426 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00525 vss 5524 5427 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00524 5428 5430 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00523 vss 5428 5429 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00522 5426 5434 5428 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00521 5524 5426 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00520 vss 5426 5524 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00519 5429 5434 5430 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00518 5430 5435 5432 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00517 vss 6580 5435 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00516 5434 5435 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00515 vss 5431 5433 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00514 5432 5433 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00513 6380 6389 6381 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00512 vss 6874 6380 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00511 6382 6385 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00510 vss 6382 6383 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00509 6381 6387 6382 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00508 6874 6381 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00507 vss 6381 6874 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00506 6383 6387 6385 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00505 6385 6389 6386 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00504 vss 6832 6389 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00503 6387 6389 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00502 vss 6384 6388 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00501 6386 6388 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00500 5000 5001 5019 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00499 vss 5244 5000 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00498 5002 5245 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00497 5019 4999 5002 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00496 vss 5245 5001 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00495 4999 5244 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00494 2997 1312 1314 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00493 1314 1313 2997 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00492 vss 1661 1314 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00491 vss 6440 1026 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00490 1026 5748 1025 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00489 1031 1025 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00488 4897 3573 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00487 5064 3979 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00486 5299 3972 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00485 4696 3759 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00484 6956 6963 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00483 vss 2352 1810 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00482 1810 3793 1934 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00481 2331 1934 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00480 1845 2161 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00479 1880 1900 1845 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00478 1844 1884 1880 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00477 vss 1888 1844 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00476 1844 2304 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00475 936 938 937 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00474 937 943 936 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00473 vss 1876 937 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00472 6063 6202 6194 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00471 vss 6571 6063 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00470 6196 6200 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00469 vss 6196 6064 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00468 6194 6201 6196 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00467 6571 6194 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00466 vss 6194 6571 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00465 6064 6201 6200 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00464 6200 6202 6065 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00463 vss 6984 6202 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00462 6201 6202 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00461 vss 6197 6198 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00460 6065 6198 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00459 3962 6876 3885 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00458 3885 6877 3962 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00457 vss 4918 3885 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00456 6791 6877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00455 vss 6876 6791 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00454 3613 4671 3501 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00453 3501 4673 3613 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00452 vss 5964 3501 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00451 1529 1534 1428 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00450 1428 3210 1529 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00449 vss 2534 1428 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00448 1527 1529 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00447 vss 6952 6435 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00446 6435 6714 6436 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00445 6434 6436 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00444 4283 4281 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00443 vss 4280 4283 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00442 4283 4285 6000 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00441 6000 4282 4283 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00440 5134 6242 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00439 4441 2979 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00438 4687 3190 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00437 4438 3403 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00436 4205 3395 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00435 1853 2542 1854 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00434 1854 3208 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00433 1852 1931 1853 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00432 2535 1932 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00431 1932 1933 1852 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00430 6882 6884 6883 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00429 vss 6885 6882 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00428 6881 6890 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00427 6883 6880 6881 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00426 vss 6890 6884 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00425 6880 6885 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00424 5087 5749 5086 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00423 5086 5748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00422 5085 6820 5087 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00421 5084 5083 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00420 5083 6440 5085 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00419 2197 2194 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00418 vss 2195 2197 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00417 2197 2196 4079 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00416 4079 2202 2197 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00415 5659 6921 5658 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00414 5658 6917 5768 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00413 vss 6963 5659 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00412 5767 5768 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00411 4015 3792 3417 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00410 3417 3793 4015 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00409 vss 3421 3417 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00408 1294 1737 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00407 1292 2506 1294 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00406 1293 1483 1292 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00405 vss 1645 1293 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00404 1293 1492 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00403 6040 6169 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00402 6336 6144 6040 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00401 920 925 998 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00400 vss 1002 920 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00399 921 923 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00398 vss 921 922 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00397 998 924 921 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00396 1002 998 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00395 vss 998 1002 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00394 922 924 923 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00393 923 925 999 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00392 vss 3259 925 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00391 924 925 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00390 vss 1001 1000 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00389 999 1000 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00388 vss 4905 5504 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00387 4905 4903 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00386 5504 4906 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00385 vss 5297 4909 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00384 4909 5084 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00383 vss 4911 4909 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00382 vss 2381 2382 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00381 2382 2379 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00380 vss 3015 2382 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00379 740 1965 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00378 vss 3229 739 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00377 1038 1982 740 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00376 739 857 1038 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00375 2301 2319 2216 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00374 2216 2483 2301 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00373 vss 2479 2216 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00372 3377 6423 3378 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00371 3378 3947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00370 3553 3376 3377 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00369 4662 6876 4663 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00368 4663 6877 4662 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00367 vss 4918 4663 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00366 4854 4662 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00365 vss 1923 1925 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00364 1923 2129 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00363 1925 2340 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00362 2650 3572 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00361 2740 2944 2650 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00360 1921 2521 1849 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00359 1848 2534 1921 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00358 1849 2512 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00357 2336 1921 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00356 vss 1918 1848 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00355 1848 1919 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00354 3384 6423 3383 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00353 3383 3947 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00352 3720 3382 3384 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00351 4342 5144 4343 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00350 4343 4523 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00349 4953 6440 4342 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00348 1082 1186 1081 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00347 1081 1323 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00346 1329 2331 1082 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00345 1125 4094 1126 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00344 1126 2352 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00343 1394 3664 1125 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00342 1100 1214 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00341 3737 1215 1100 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00340 2945 3186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00339 2944 5742 2945 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00338 vss 1907 1911 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00337 1907 2333 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00336 1911 3391 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00335 3595 3413 3410 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00334 3410 3414 3595 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00333 vss 5372 3410 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00332 6409 6806 6408 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00331 6408 6631 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00330 6410 6906 6409 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00329 vss 5505 5506 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00328 5506 5504 5507 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00327 5975 5507 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00326 vss 5127 4821 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00325 4821 5132 4950 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00324 5561 4950 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00323 vss 5342 5227 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00322 5227 5343 5344 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00321 5557 5344 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00320 vss 2993 2780 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00319 2780 2990 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00318 2778 2780 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00317 737 2830 738 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00316 738 860 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00315 736 5069 737 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00314 851 6440 736 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00313 687 2830 688 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00312 688 1385 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00311 685 5069 687 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00310 686 6440 685 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00309 4724 4731 4723 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00308 4723 4722 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00307 4720 4947 4724 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00306 6852 6876 6853 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00305 6853 6877 6852 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00304 vss 6850 6853 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00303 6851 6852 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00302 6869 6866 6868 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00301 6868 6875 6869 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00300 vss 6867 6868 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00299 6396 6791 6395 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00298 6397 6648 6396 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00297 6395 6678 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00296 6393 6396 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00295 vss 6637 6397 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00294 6397 6883 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00293 6804 6808 6803 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00292 6803 6801 6805 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00291 vss 6802 6804 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00290 6800 6805 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00289 3236 4083 3114 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00288 3114 4082 3236 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00287 vss 5272 3114 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00286 3016 3816 3017 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00285 3017 3227 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00284 3014 5116 3016 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00283 3015 3218 3014 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00282 2392 4748 2253 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00281 vss 4235 2391 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00280 2253 2391 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00279 4783 5068 4784 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00278 4784 5102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00277 4782 5069 4783 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00276 4899 4901 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00275 4901 5262 4782 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00274 6871 6893 6873 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00273 6873 6885 6872 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00272 vss 6906 6871 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00271 6870 6872 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00270 3852 5341 3851 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00269 3850 3853 3852 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00268 3851 5575 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00267 6876 3852 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00266 vss 3849 3850 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00265 3850 3856 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00264 2772 2773 2666 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00263 2665 5959 2772 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00262 2666 4438 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00261 2770 2772 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00260 vss 3199 2665 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00259 2665 3618 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00258 1052 4524 1051 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00257 1051 4094 1053 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00256 vss 5363 1052 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00255 1779 1053 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00254 2411 2629 2209 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00253 2209 2418 2411 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00252 vss 2208 2209 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00251 1847 2102 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00250 1891 2095 1847 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00249 1846 2485 1891 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00248 vss 2319 1846 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00247 1846 2320 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00246 6008 6448 6007 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00245 6007 6449 6009 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00244 vss 6917 6008 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00243 6013 6009 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00242 4745 5773 4746 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00241 4746 5575 4745 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00240 vss 5889 4746 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00239 2266 2412 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00238 3060 2406 2266 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00237 1024 1031 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00236 1214 5749 1024 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00235 1023 1732 1214 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00234 vss 1231 1023 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00233 1023 1218 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00232 vss 2198 1470 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00231 1470 2409 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00230 1583 1586 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00229 1470 1587 1586 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00228 1586 2799 1470 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00227 vss 1893 1406 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00226 1406 1641 1489 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00225 1488 1489 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00224 1290 1645 1291 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00223 1291 1492 1290 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00222 vss 1483 1291 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00221 1289 1290 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00220 2927 2935 2928 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00219 vss 3560 2927 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00218 2929 2931 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00217 vss 2929 2930 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00216 2928 2933 2929 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00215 3560 2928 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00214 vss 2928 3560 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00213 2930 2933 2931 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00212 2931 2935 2932 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00211 vss 3160 2935 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00210 2933 2935 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00209 vss 3563 2934 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00208 2932 2934 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00207 1118 1985 1117 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00206 1117 1235 1230 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00205 vss 1579 1118 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00204 1229 1230 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00203 2506 1231 1027 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00202 1027 1218 2506 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00201 vss 1732 1027 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00200 vss 2936 2648 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00199 2648 3172 2738 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00198 2737 2738 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00197 5232 5360 5351 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00196 vss 5349 5232 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00195 5352 5355 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00194 vss 5352 5233 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00193 5351 5357 5352 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00192 5349 5351 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00191 vss 5351 5349 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00190 5233 5357 5355 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00189 5355 5360 5234 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00188 vss 6984 5360 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00187 5357 5360 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00186 vss 5354 5358 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00185 5234 5358 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00184 6862 6865 6866 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00183 vss 6861 6862 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00182 6864 6870 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00181 6866 6863 6864 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00180 vss 6870 6865 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00179 6863 6861 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00178 63 62 305 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00177 vss 470 63 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00176 65 196 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00175 305 64 65 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00174 vss 196 62 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00173 64 470 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00172 4602 5039 4603 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00171 4603 5877 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00170 4601 5992 4602 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00169 4695 4694 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00168 4694 6440 4601 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00167 158 787 157 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00166 157 493 215 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00165 vss 2314 158 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00164 319 215 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00163 497 986 438 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00162 438 987 497 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00161 vss 500 438 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00160 919 497 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00159 1861 2610 1862 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00158 1862 1971 1970 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00157 vss 2607 1861 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00156 1968 1970 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00155 3169 3740 3129 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00154 3128 5902 3169 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00153 3129 5064 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00152 3167 3169 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00151 vss 3737 3128 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00150 3128 3738 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00149 2231 2512 2230 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00148 2230 2511 2332 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00147 vss 2331 2231 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00146 2518 2332 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00145 3531 4748 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00144 3645 3662 3531 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00143 3530 5372 3645 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00142 vss 4083 3530 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00141 3530 4082 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00140 5158 5167 5159 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00139 vss 5157 5158 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00138 5160 5162 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00137 vss 5160 5163 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00136 5159 5166 5160 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00135 5157 5159 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00134 vss 5159 5157 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00133 5163 5166 5162 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00132 5162 5167 5161 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00131 vss 6984 5167 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00130 5166 5167 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00129 vss 5164 5165 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00128 5161 5165 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00127 3416 3413 3415 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00126 3415 3414 3416 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00125 vss 5902 3415 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00124 2063 2068 2167 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00123 vss 2583 2063 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00122 2064 2065 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00121 vss 2064 2066 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00120 2167 2067 2064 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00119 2583 2167 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00118 vss 2167 2583 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00117 2066 2067 2065 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00116 2065 2068 2168 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00115 vss 3259 2068 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00114 2067 2068 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00113 vss 2582 2169 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00112 2168 2169 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00111 5237 5570 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00110 5369 5788 5237 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00109 3589 3413 3409 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00108 3409 3414 3589 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00107 vss 5243 3409 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00106 3480 3727 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00105 3563 3971 3480 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00104 6041 6154 6145 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00103 vss 6820 6041 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00102 6149 6148 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00101 vss 6149 6042 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00100 6145 6153 6149 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00099 6820 6145 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00098 vss 6145 6820 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00097 6042 6153 6148 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00096 6148 6154 6043 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00095 vss 6832 6154 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00094 6153 6154 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00093 vss 6150 6151 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00092 6043 6151 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00091 5126 5125 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00090 5337 6447 5126 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00089 1657 2356 1658 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00088 1656 2314 1657 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00087 1658 2111 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00086 1655 1657 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00085 vss 3740 1656 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00084 1656 2553 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00083 2546 3199 2543 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00082 2543 3618 2546 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00081 vss 5725 2543 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00080 403 2195 404 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00079 404 2194 403 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00078 vss 1033 404 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00077 402 403 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00076 1803 1898 2107 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00075 vss 1905 1803 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00074 1804 2320 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00073 2107 1897 1804 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00072 vss 2320 1898 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00071 1897 1905 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00070 6057 6178 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00069 6384 6180 6057 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00068 4369 4610 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00067 4465 5088 4369 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00066 5095 5986 5096 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00065 5096 6214 5095 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00064 vss 6820 5096 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00063 5094 5095 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00062 5527 5753 5526 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00061 5526 5767 5527 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00060 vss 5524 5526 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00059 5525 5527 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00058 3834 5992 3833 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00057 3833 4265 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00056 4253 6440 3834 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00055 2409 5359 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00054 vss 5144 2409 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00053 1388 1991 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00052 1746 1779 1388 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00051 6399 6400 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00050 6652 6398 6399 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00049 3435 5069 3436 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00048 3436 5068 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00047 3816 5575 3435 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00046 4333 5992 4332 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00045 4332 4726 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00044 5116 6440 4333 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00043 3103 5068 3104 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00042 3104 4062 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00041 3218 5069 3103 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00040 1469 4089 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00039 1582 2412 1469 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00038 1120 1582 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00037 1231 2625 1120 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00036 2347 3199 2235 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00035 2235 3618 2347 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00034 vss 6187 2235 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00033 2937 3186 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00032 2936 5963 2937 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00031 2647 3172 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00030 2736 2936 2647 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00029 vss 6591 6499 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00028 6499 6616 6592 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00027 6590 6592 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00026 vss 1708 1707 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00025 1707 1706 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00024 2052 1707 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00023 1857 2553 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00022 1945 2356 1857 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00021 83 772 82 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00020 82 212 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00019 81 1151 83 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00018 80 772 79 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00017 79 86 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00016 209 1151 80 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00015 6717 6723 6718 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00014 6567 6724 6717 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00013 6952 6717 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00012 vss 6717 6952 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00011 6570 6721 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00010 vss 6967 6721 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00009 6723 6724 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00008 vss 6984 6724 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00007 6568 6720 vss vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00006 6718 6976 6568 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00005 6720 6724 6570 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00004 6569 6723 6720 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00003 vss 6718 6569 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00002 vss 6952 6566 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00001 6566 6976 6567 vss sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
.ends m65_cts_r_ext

