* Spice description of noa3ao322_x4
* Spice driver version -663785701
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:15

* INTERF i0 i1 i2 i3 i4 i5 i6 nq vdd vss 


.subckt noa3ao322_x4 13 7 8 6 5 4 9 14 3 17 
* NET 3 = vdd
* NET 4 = i5
* NET 5 = i4
* NET 6 = i3
* NET 7 = i1
* NET 8 = i2
* NET 9 = i6
* NET 13 = i0
* NET 14 = nq
* NET 17 = vss
Mtr_00020 2 4 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00019 1 5 15 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00018 15 6 15 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00017 2 8 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00016 15 9 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00015 3 7 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.87U AS=0.4488P AD=0.4488P PS=4.22U PD=4.22U 
Mtr_00014 2 13 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.87U AS=0.4488P AD=0.4488P PS=4.22U PD=4.22U 
Mtr_00013 14 16 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 3 16 14 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 3 15 16 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00010 14 16 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00009 17 4 10 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.68U AS=0.1632P AD=0.1632P PS=1.84U PD=1.84U 
Mtr_00008 10 5 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.68U AS=0.1632P AD=0.1632P PS=1.84U PD=1.84U 
Mtr_00007 17 6 10 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.68U AS=0.1632P AD=0.1632P PS=1.84U PD=1.84U 
Mtr_00006 12 13 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.36U AS=0.3264P AD=0.3264P PS=3.2U PD=3.2U 
Mtr_00005 11 7 12 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.36U AS=0.3264P AD=0.3264P PS=3.2U PD=3.2U 
Mtr_00004 17 16 14 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00003 15 8 11 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.36U AS=0.3264P AD=0.3264P PS=3.2U PD=3.2U 
Mtr_00002 10 9 15 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.02U AS=0.2448P AD=0.2448P PS=2.52U PD=2.52U 
Mtr_00001 17 15 16 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
C16 2 17 1.24896e-15
C15 3 17 4.5163e-15
C14 4 17 1.77053e-15
C13 5 17 1.73747e-15
C12 6 17 1.78042e-15
C11 7 17 1.69828e-15
C10 8 17 1.39425e-15
C9 9 17 1.35774e-15
C8 10 17 5.43814e-16
C5 13 17 1.70741e-15
C4 14 17 2.15173e-15
C3 15 17 2.88659e-15
C2 16 17 2.06732e-15
C1 17 17 4.17598e-15
.ends noa3ao322_x4

