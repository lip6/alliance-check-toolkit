* or21nand_x0
.subckt or21nand_x0 vdd vss nq i0 i1 i2
Mi0_nmos _net0 i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi0_pmos vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi1_nmos vss i1 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi1_pmos _net1 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mi2_nmos _net0 i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mi2_pmos nq i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends or21nand_x0
