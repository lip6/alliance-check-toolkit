* Spice description of mac_cts_r_ext_ihp
* Spice driver version 1906871213
* Date ( dd/mm/yyyy hh:mm:ss ): 30/09/2024 at 15:39:46

* INTERF accumulator_out[0] accumulator_out[1] accumulator_out[2] 
* INTERF accumulator_out[3] accumulator_out[4] accumulator_out[5] 
* INTERF accumulator_out[6] accumulator_out[7] clk multiplicand[0] 
* INTERF multiplicand[1] multiplicand[2] multiplicand[3] multiplier[0] 
* INTERF multiplier[1] multiplier[2] multiplier[3] reset vdd vss 


.subckt mac_cts_r_ext_ihp 274 79 112 171 946 945 928 910 497 674 736 686 710 722 711 673 675 777 909 947 
* NET 15 = subckt_159_sff1_x4.sff_s
* NET 19 = subckt_159_sff1_x4.sff_m
* NET 21 = subckt_159_sff1_x4.ckr
* NET 22 = subckt_159_sff1_x4.nckr
* NET 26 = subckt_158_sff1_x4.sff_s
* NET 30 = subckt_158_sff1_x4.sff_m
* NET 31 = subckt_158_sff1_x4.ckr
* NET 33 = subckt_158_sff1_x4.nckr
* NET 44 = abc_567_auto_rtlil_cc_2608_muxgate_558
* NET 52 = subckt_157_sff1_x4.sff_s
* NET 55 = subckt_157_sff1_x4.sff_m
* NET 61 = subckt_157_sff1_x4.ckr
* NET 62 = subckt_157_sff1_x4.nckr
* NET 72 = abc_567_new_n148
* NET 76 = abc_567_new_n149
* NET 79 = accumulator_out[1]
* NET 83 = abc_567_new_n153
* NET 86 = abc_567_new_n157
* NET 93 = abc_567_auto_rtlil_cc_2608_muxgate_556
* NET 94 = abc_567_new_n151
* NET 99 = abc_567_new_n143
* NET 107 = abc_567_new_n156
* NET 112 = accumulator_out[2]
* NET 113 = abc_567_new_n142
* NET 114 = abc_567_new_n141
* NET 117 = abc_567_auto_rtlil_cc_2608_muxgate_554
* NET 118 = abc_567_new_n144
* NET 122 = spare_buffer_82.q
* NET 128 = spare_buffer_78.q
* NET 129 = spare_buffer_66.q
* NET 131 = spare_buffer_62.q
* NET 136 = spare_buffer_81.q
* NET 139 = abc_567_new_n147
* NET 140 = abc_567_new_n146
* NET 141 = abc_567_new_n150
* NET 143 = abc_567_new_n42
* NET 145 = spare_buffer_77.q
* NET 148 = abc_567_new_n138
* NET 149 = spare_buffer_65.q
* NET 152 = spare_buffer_61.q
* NET 154 = spare_buffer_60.q
* NET 171 = accumulator_out[3]
* NET 174 = subckt_149_sff1_x4.sff_s
* NET 177 = subckt_149_sff1_x4.sff_m
* NET 183 = subckt_149_sff1_x4.ckr
* NET 184 = subckt_149_sff1_x4.nckr
* NET 186 = subckt_156_sff1_x4.sff_s
* NET 189 = subckt_156_sff1_x4.sff_m
* NET 193 = subckt_156_sff1_x4.ckr
* NET 195 = clk_root_tl_tr_0
* NET 196 = subckt_156_sff1_x4.nckr
* NET 207 = partial_product[2]
* NET 210 = subckt_150_sff1_x4.sff_s
* NET 213 = abc_567_auto_rtlil_cc_2608_muxgate_540
* NET 215 = subckt_150_sff1_x4.sff_m
* NET 216 = clk_root_tr_tl_0
* NET 218 = subckt_150_sff1_x4.ckr
* NET 219 = subckt_150_sff1_x4.nckr
* NET 220 = abc_567_new_n43
* NET 221 = abc_567_auto_rtlil_cc_2608_muxgate_538
* NET 222 = partial_product[1]
* NET 227 = abc_567_auto_rtlil_cc_2608_muxgate_552
* NET 235 = partial_product[3]
* NET 236 = subckt_151_sff1_x4.sff_s
* NET 242 = subckt_151_sff1_x4.sff_m
* NET 244 = clk_root_tr_tr_0
* NET 245 = subckt_151_sff1_x4.ckr
* NET 247 = subckt_151_sff1_x4.nckr
* NET 248 = abc_567_new_n52
* NET 251 = abc_567_new_n160
* NET 252 = abc_567_new_n155
* NET 262 = abc_567_new_n65
* NET 266 = abc_567_auto_rtlil_cc_2608_muxgate_542
* NET 267 = abc_567_new_n159
* NET 269 = abc_567_new_n154
* NET 271 = abc_567_new_n139
* NET 274 = accumulator_out[0]
* NET 289 = abc_567_auto_rtlil_cc_2608_muxgate_536
* NET 291 = abc_567_new_n51
* NET 295 = subckt_148_sff1_x4.sff_s
* NET 296 = partial_product[0]
* NET 297 = subckt_148_sff1_x4.sff_m
* NET 303 = subckt_148_sff1_x4.ckr
* NET 304 = subckt_148_sff1_x4.nckr
* NET 313 = abc_567_new_n56
* NET 315 = abc_567_new_n47
* NET 319 = abc_567_new_n55
* NET 321 = abc_567_new_n50
* NET 325 = abc_567_new_n63
* NET 329 = abc_567_new_n161
* NET 334 = abc_567_new_n166
* NET 350 = abc_567_new_n91
* NET 354 = subckt_160_sff1_x4.sff_s
* NET 359 = abc_567_auto_rtlil_cc_2608_muxgate_560
* NET 361 = subckt_160_sff1_x4.sff_m
* NET 363 = subckt_160_sff1_x4.ckr
* NET 364 = subckt_160_sff1_x4.nckr
* NET 370 = abc_567_new_n59
* NET 372 = abc_567_new_n49
* NET 374 = abc_567_new_n60
* NET 375 = abc_567_new_n61
* NET 379 = abc_567_new_n164
* NET 386 = spare_buffer_74.q
* NET 388 = abc_567_new_n84
* NET 389 = abc_567_new_n62
* NET 390 = abc_567_new_n88
* NET 392 = spare_buffer_70.q
* NET 394 = spare_buffer_58.q
* NET 396 = spare_buffer_54.q
* NET 406 = subckt_152_sff1_x4.sff_m
* NET 407 = spare_buffer_73.q
* NET 409 = spare_buffer_72.q
* NET 411 = spare_buffer_69.q
* NET 413 = clk_root_tr_0
* NET 414 = spare_buffer_68.q
* NET 416 = subckt_152_sff1_x4.sff_s
* NET 421 = subckt_152_sff1_x4.ckr
* NET 422 = subckt_152_sff1_x4.nckr
* NET 423 = spare_buffer_57.q
* NET 425 = clk_root_tl_br_0
* NET 427 = spare_buffer_53.q
* NET 429 = spare_buffer_52.q
* NET 430 = clk_root_tl_0
* NET 439 = abc_567_new_n87
* NET 445 = abc_567_new_n58
* NET 449 = abc_567_new_n85
* NET 451 = abc_567_new_n89
* NET 463 = abc_567_new_n54
* NET 464 = abc_567_new_n86
* NET 467 = abc_567_new_n83
* NET 469 = abc_567_new_n113
* NET 470 = abc_567_new_n112
* NET 471 = abc_567_new_n93
* NET 472 = abc_567_auto_rtlil_cc_2608_muxgate_544
* NET 474 = abc_567_new_n100
* NET 477 = abc_567_new_n81
* NET 479 = abc_567_new_n82
* NET 482 = abc_567_new_n94
* NET 485 = abc_567_new_n110
* NET 493 = abc_567_new_n79
* NET 497 = clk
* NET 502 = abc_567_new_n57
* NET 506 = abc_567_new_n78
* NET 507 = abc_567_new_n67
* NET 513 = abc_567_new_n95
* NET 515 = abc_567_new_n108
* NET 521 = abc_567_new_n107
* NET 526 = abc_567_new_n101
* NET 535 = abc_567_new_n66
* NET 536 = abc_567_new_n80
* NET 540 = abc_567_new_n103
* NET 541 = abc_567_new_n104
* NET 543 = abc_567_new_n99
* NET 548 = abc_567_new_n74
* NET 552 = abc_567_new_n76
* NET 555 = abc_567_new_n90
* NET 556 = abc_567_new_n111
* NET 568 = abc_567_new_n75
* NET 569 = abc_567_new_n70
* NET 571 = abc_567_new_n77
* NET 572 = abc_567_new_n105
* NET 573 = abc_567_new_n106
* NET 576 = abc_567_new_n118
* NET 581 = spare_buffer_50.q
* NET 583 = abc_567_new_n97
* NET 586 = spare_buffer_46.q
* NET 588 = abc_567_new_n116
* NET 593 = spare_buffer_34.q
* NET 595 = spare_buffer_30.q
* NET 600 = spare_buffer_49.q
* NET 601 = spare_buffer_48.q
* NET 603 = abc_567_new_n109
* NET 606 = spare_buffer_45.q
* NET 609 = spare_buffer_44.q
* NET 610 = abc_567_new_n120
* NET 612 = spare_buffer_33.q
* NET 614 = spare_buffer_32.q
* NET 616 = spare_buffer_29.q
* NET 618 = spare_buffer_28.q
* NET 622 = abc_567_new_n72
* NET 625 = abc_567_new_n98
* NET 631 = abc_567_new_n124
* NET 632 = abc_567_new_n119
* NET 643 = abc_567_new_n68
* NET 645 = abc_567_new_n121
* NET 646 = abc_567_new_n117
* NET 647 = abc_567_new_n122
* NET 650 = abc_567_new_n69
* NET 660 = abc_567_new_n115
* NET 663 = abc_567_new_n123
* NET 673 = multiplier[2]
* NET 674 = multiplicand[0]
* NET 675 = multiplier[3]
* NET 676 = abc_567_new_n71
* NET 677 = abc_567_new_n127
* NET 679 = abc_567_new_n102
* NET 680 = abc_567_new_n44
* NET 681 = abc_567_new_n45
* NET 685 = abc_567_new_n73
* NET 686 = multiplicand[2]
* NET 688 = abc_567_new_n132
* NET 690 = abc_567_new_n129
* NET 691 = abc_567_new_n131
* NET 692 = abc_567_new_n130
* NET 694 = clk_root_0
* NET 702 = abc_567_new_n96
* NET 710 = multiplicand[3]
* NET 711 = multiplier[1]
* NET 715 = abc_567_new_n125
* NET 722 = multiplier[0]
* NET 726 = subckt_154_sff1_x4.sff_m
* NET 727 = abc_567_auto_rtlil_cc_2608_muxgate_548
* NET 728 = subckt_154_sff1_x4.ckr
* NET 733 = abc_567_auto_rtlil_cc_2608_muxgate_546
* NET 734 = subckt_153_sff1_x4.sff_m
* NET 735 = subckt_153_sff1_x4.ckr
* NET 736 = multiplicand[1]
* NET 742 = abc_567_new_n128
* NET 743 = abc_567_new_n133
* NET 744 = abc_567_new_n136
* NET 747 = subckt_154_sff1_x4.sff_s
* NET 750 = subckt_154_sff1_x4.nckr
* NET 753 = subckt_153_sff1_x4.sff_s
* NET 756 = subckt_153_sff1_x4.nckr
* NET 768 = subckt_155_sff1_x4.sff_s
* NET 772 = subckt_155_sff1_x4.sff_m
* NET 773 = abc_567_auto_rtlil_cc_2608_muxgate_550
* NET 775 = subckt_155_sff1_x4.ckr
* NET 776 = subckt_155_sff1_x4.nckr
* NET 777 = reset
* NET 778 = abc_567_new_n134
* NET 779 = abc_567_new_n163
* NET 792 = partial_product[7]
* NET 795 = partial_product[4]
* NET 798 = subckt_161_sff1_x4.sff_s
* NET 801 = subckt_161_sff1_x4.sff_m
* NET 803 = abc_567_auto_rtlil_cc_2608_muxgate_562
* NET 808 = subckt_161_sff1_x4.ckr
* NET 809 = subckt_161_sff1_x4.nckr
* NET 813 = spare_buffer_42.q
* NET 815 = abc_567_new_n162
* NET 816 = abc_567_new_n165
* NET 819 = spare_buffer_38.q
* NET 821 = abc_567_new_n168
* NET 822 = abc_567_new_n173
* NET 825 = spare_buffer_26.q
* NET 827 = spare_buffer_22.q
* NET 831 = spare_buffer_41.q
* NET 834 = abc_567_new_n175
* NET 837 = spare_buffer_37.q
* NET 839 = clk_root_br_0
* NET 841 = abc_567_new_n172
* NET 847 = spare_buffer_25.q
* NET 849 = clk_root_bl_br_0
* NET 851 = spare_buffer_21.q
* NET 853 = spare_buffer_20.q
* NET 854 = clk_root_bl_0
* NET 861 = abc_567_new_n171
* NET 865 = abc_567_new_n178
* NET 866 = abc_567_new_n185
* NET 867 = abc_567_new_n176
* NET 871 = abc_567_new_n181
* NET 872 = abc_567_new_n186
* NET 879 = abc_567_new_n180
* NET 880 = abc_567_new_n169
* NET 888 = abc_567_new_n187
* NET 889 = abc_567_new_n188
* NET 892 = abc_567_new_n179
* NET 897 = abc_567_new_n183
* NET 898 = abc_567_new_n182
* NET 899 = abc_567_new_n46
* NET 909 = vdd
* NET 910 = accumulator_out[7]
* NET 911 = subckt_163_sff1_x4.sff_s
* NET 914 = subckt_163_sff1_x4.sff_m
* NET 916 = abc_567_auto_rtlil_cc_2608_muxgate_566
* NET 921 = clk_root_br_br_0
* NET 922 = subckt_163_sff1_x4.ckr
* NET 923 = subckt_163_sff1_x4.nckr
* NET 924 = abc_567_new_n177
* NET 925 = partial_product[6]
* NET 928 = accumulator_out[6]
* NET 929 = subckt_162_sff1_x4.sff_s
* NET 933 = abc_567_auto_rtlil_cc_2608_muxgate_564
* NET 936 = subckt_162_sff1_x4.sff_m
* NET 938 = clk_root_br_bl_0
* NET 939 = subckt_162_sff1_x4.ckr
* NET 941 = subckt_162_sff1_x4.nckr
* NET 942 = abc_567_new_n170
* NET 943 = partial_product[5]
* NET 945 = accumulator_out[5]
* NET 946 = accumulator_out[4]
* NET 947 = vss
Mtr_02090 909 839 818 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02089 819 818 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02088 909 818 819 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02087 909 818 819 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02086 819 818 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02085 909 854 596 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02084 595 596 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02083 909 596 595 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02082 909 596 595 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02081 595 596 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02080 909 854 615 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02079 614 615 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02078 909 615 614 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02077 909 615 614 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02076 614 615 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02075 909 854 613 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02074 612 613 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02073 909 613 612 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02072 909 613 612 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02071 612 613 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02070 909 854 594 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02069 593 594 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02068 909 594 593 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02067 909 594 593 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02066 593 594 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02065 909 839 840 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02064 938 840 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02063 909 840 938 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02062 909 840 938 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02061 938 840 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02060 909 839 838 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02059 837 838 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02058 909 838 837 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02057 909 838 837 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02056 837 838 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02055 909 854 855 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02054 853 855 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02053 909 855 853 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02052 909 855 853 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02051 853 855 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02050 909 854 852 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02049 851 852 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02048 909 852 851 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02047 909 852 851 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02046 851 852 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02045 909 854 828 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02044 827 828 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02043 909 828 827 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02042 909 828 827 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02041 827 828 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02040 909 854 850 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02039 849 850 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02038 909 850 849 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02037 909 850 849 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02036 849 850 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02035 909 854 848 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02034 847 848 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02033 909 848 847 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02032 909 848 847 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02031 847 848 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02030 909 854 826 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02029 825 826 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02028 909 826 825 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02027 909 826 825 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02026 825 826 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02025 909 854 619 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02024 618 619 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02023 909 619 618 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02022 909 619 618 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02021 618 619 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02020 909 854 617 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02019 616 617 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02018 909 617 616 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02017 909 617 616 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02016 616 617 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02015 45 86 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02014 909 899 45 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02013 44 45 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02012 449 493 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02011 449 479 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02010 909 477 449 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_02009 909 694 305 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02008 430 305 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02007 909 305 430 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02006 909 305 430 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02005 430 305 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02004 909 694 292 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02003 413 292 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02002 909 292 413 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02001 909 292 413 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_02000 413 292 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01999 366 795 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01998 909 795 384 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01997 381 946 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01996 909 381 366 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01995 366 384 382 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01994 382 946 366 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01993 379 382 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01992 909 382 379 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01991 213 169 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01990 157 325 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01989 909 777 170 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01988 909 207 156 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01987 156 170 169 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01986 169 777 157 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01985 502 711 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01984 502 673 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01983 909 736 502 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01982 909 674 502 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01981 177 183 161 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01980 160 184 177 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01979 909 176 160 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01978 176 177 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01977 174 184 176 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01976 909 216 184 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01975 183 184 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01974 909 221 182 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01973 161 182 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01972 159 158 174 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01971 909 222 159 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01970 222 174 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01969 909 174 222 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01968 734 735 716 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01967 717 756 734 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01966 909 731 717 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01965 731 734 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01964 753 756 731 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01963 909 849 756 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01962 735 756 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01961 909 733 758 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01960 716 758 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01959 714 721 753 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01958 909 943 714 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01957 943 753 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01956 909 753 943 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01955 471 777 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01954 909 795 471 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01953 605 631 604 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01952 604 603 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01951 909 647 605 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01950 677 605 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01949 221 223 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01948 225 248 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01947 909 777 226 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01946 909 222 224 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01945 224 226 223 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01944 223 777 225 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01943 909 379 333 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01942 318 379 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01941 334 329 318 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01940 318 333 334 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01939 909 331 318 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01938 331 329 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01937 942 943 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01936 909 945 942 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01935 909 515 512 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01934 499 515 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01933 556 513 499 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01932 499 512 556 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01931 909 511 499 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01930 511 513 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01929 242 245 231 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01928 230 247 242 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01927 909 238 230 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01926 238 242 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01925 236 247 238 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01924 909 244 247 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01923 245 247 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01922 909 266 246 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01921 231 246 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01920 229 234 236 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01919 909 235 229 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01918 235 236 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01917 909 236 235 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01916 685 686 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01915 909 711 685 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01914 119 118 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01913 909 899 119 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01912 117 119 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01911 252 235 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01910 909 171 252 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01909 648 736 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01908 909 673 648 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01907 650 652 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01906 652 674 648 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01905 648 675 652 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01904 205 777 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01903 909 235 205 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01902 262 205 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01901 447 445 443 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01900 443 463 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01899 909 502 447 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01898 535 447 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01897 316 722 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01896 909 674 316 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01895 315 316 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01894 438 506 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01893 439 536 438 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01892 909 467 439 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01891 389 374 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01890 909 372 389 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01889 890 888 891 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01888 891 889 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01887 909 899 890 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01886 916 890 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01885 927 925 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01884 909 928 927 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01883 924 927 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01882 690 686 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01881 690 710 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01880 909 675 690 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01879 909 673 690 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01878 319 736 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01877 909 711 319 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01876 909 555 351 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01875 351 390 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01874 909 899 351 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01873 350 351 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01872 73 72 74 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01871 74 140 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01870 909 139 73 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01869 83 73 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01868 909 207 23 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01867 23 112 72 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01866 909 222 43 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01865 43 79 113 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01864 251 124 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01863 124 139 121 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01862 909 143 121 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01861 121 220 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01860 120 140 124 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01859 121 141 120 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01858 909 497 498 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01857 694 498 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01856 909 498 694 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01855 909 498 694 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01854 694 498 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01853 909 694 695 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01852 854 695 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01851 909 695 854 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01850 909 695 854 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01849 854 695 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01848 909 694 687 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01847 839 687 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01846 909 687 839 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01845 909 687 839 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01844 839 687 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01843 909 622 549 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01842 549 676 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01841 909 650 549 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01840 548 549 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01839 881 943 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01838 909 945 881 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01837 880 881 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01836 781 816 821 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01835 780 779 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01834 909 780 781 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01833 909 540 517 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01832 500 540 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01831 521 583 500 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01830 500 517 521 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01829 909 519 500 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01828 519 583 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01827 909 675 655 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01826 655 710 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01825 655 686 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01824 909 673 655 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01823 742 655 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01822 873 871 869 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01821 869 924 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01820 909 872 873 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01819 888 873 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01818 95 94 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01817 909 899 95 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01816 93 95 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01815 475 552 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01814 477 548 475 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01813 909 535 477 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01812 909 777 744 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01811 909 792 705 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01810 744 705 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01809 678 691 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01808 909 677 678 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01807 688 678 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01806 624 686 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01805 909 711 624 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01804 622 624 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01803 453 485 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01802 909 451 453 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01801 470 453 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01800 250 291 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01799 909 321 250 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01798 248 250 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01797 30 31 29 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01796 28 33 30 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01795 909 27 28 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01794 27 30 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01793 26 33 27 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01792 909 216 33 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01791 31 33 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01790 909 93 32 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01789 29 32 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01788 24 25 26 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01787 909 112 24 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01786 112 26 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01785 909 26 112 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01784 936 939 908 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01783 907 941 936 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01782 909 931 907 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01781 931 936 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01780 929 941 931 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01779 909 938 941 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01778 939 941 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01777 909 933 940 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01776 908 940 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01775 906 905 929 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01774 909 928 906 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01773 928 929 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01772 909 929 928 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01771 253 251 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01770 909 252 253 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01769 329 253 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01768 909 143 144 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01767 144 220 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01766 267 139 144 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01765 142 140 267 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01764 144 141 142 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01763 570 643 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01762 571 569 570 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01761 909 685 571 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01760 442 675 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01759 909 736 442 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01758 526 442 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01757 327 374 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01756 909 372 327 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01755 375 327 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01754 644 691 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01753 743 677 644 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01752 909 899 743 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01751 909 350 264 909 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_01750 266 265 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01749 264 263 265 909 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_01748 148 296 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01747 909 274 148 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01746 778 777 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01745 909 925 778 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01744 835 834 829 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01743 829 880 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01742 909 892 835 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01741 871 835 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01740 909 645 627 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01739 621 645 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01738 631 646 621 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01737 621 627 631 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01736 909 629 621 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01735 629 646 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01734 909 571 510 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01733 510 568 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01732 909 507 510 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01731 506 510 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01730 558 556 546 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01729 546 555 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01728 909 603 558 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01727 660 558 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01726 718 792 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01725 909 792 738 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01724 737 910 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01723 909 737 718 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01722 718 738 741 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01721 741 910 718 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01720 866 741 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01719 909 741 866 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01718 909 207 92 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01717 81 207 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01716 141 112 81 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01715 81 92 141 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01714 909 89 81 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01713 89 112 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01712 189 193 165 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01711 164 196 189 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01710 909 187 164 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01709 187 189 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01708 186 196 187 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01707 909 195 196 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01706 193 196 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01705 909 227 194 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01704 165 194 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01703 162 163 186 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01702 909 274 162 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01701 274 186 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01700 909 186 274 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01699 691 692 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01698 909 690 691 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01697 361 363 360 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01696 357 364 361 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01695 909 356 357 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01694 356 361 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01693 354 364 356 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01692 909 425 364 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01691 363 364 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01690 909 359 362 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01689 360 362 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01688 355 353 354 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01687 909 946 355 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01686 946 354 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01685 909 354 946 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01684 909 841 824 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01683 823 841 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01682 822 821 823 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01681 823 824 822 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01680 909 820 823 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01679 820 821 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01678 314 673 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01677 909 674 314 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01676 313 314 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01675 681 710 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01674 220 235 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01673 473 469 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01672 472 470 473 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01671 909 471 472 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01670 830 943 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01669 909 943 846 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01668 842 945 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01667 909 842 830 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01666 830 846 845 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01665 845 945 830 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01664 841 845 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01663 909 845 841 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01662 909 526 457 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01661 444 526 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01660 540 474 444 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01659 444 457 540 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01658 909 454 444 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01657 454 474 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01656 576 710 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01655 909 673 576 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01654 676 736 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01653 676 675 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01652 909 673 676 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01651 909 674 676 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01650 440 536 441 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01649 441 467 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01648 909 493 440 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01647 482 440 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01646 555 375 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01645 555 439 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01644 909 449 555 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01643 909 313 71 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01642 70 313 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01641 370 319 70 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01640 70 71 370 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01639 909 69 70 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01638 69 319 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01637 726 728 708 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01636 709 750 726 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01635 909 724 709 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01634 724 726 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01633 747 750 724 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01632 909 938 750 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01631 728 750 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01630 909 727 752 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01629 708 752 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01628 707 720 747 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01627 909 925 707 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01626 925 747 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01625 909 747 925 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01624 909 374 326 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01623 317 374 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01622 325 321 317 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01621 317 326 325 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01620 909 322 317 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01619 322 321 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01618 572 540 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01617 909 625 572 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01616 603 515 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01615 909 513 603 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01614 437 463 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01613 507 445 437 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01612 909 502 507 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01611 909 711 293 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01610 293 736 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01609 293 722 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01608 909 674 293 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01607 372 293 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01606 468 467 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01605 513 536 468 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01604 909 493 513 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01603 321 722 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01602 321 736 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01601 909 711 321 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01600 909 674 321 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01599 493 507 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01598 493 571 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01597 909 568 493 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01596 568 650 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01595 568 622 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01594 909 676 568 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01593 909 792 793 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01592 783 792 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01591 872 910 783 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01590 783 793 872 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01589 909 790 783 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01588 790 910 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01587 111 235 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01586 909 235 109 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01585 108 171 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01584 909 108 111 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01583 111 109 110 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01582 110 171 111 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01581 107 110 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01580 909 110 107 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01579 474 686 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01578 909 673 474 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01577 702 710 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01576 909 711 702 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01575 865 925 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01574 909 928 865 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01573 348 736 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01572 909 711 348 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01571 445 674 348 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01570 348 673 445 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01569 228 271 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01568 909 899 228 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01567 227 228 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01566 611 632 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01565 909 679 611 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01564 610 611 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01563 289 257 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01562 233 315 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01561 909 777 258 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01560 909 296 232 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01559 232 258 257 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01558 257 777 233 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01557 642 673 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01556 909 736 642 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01555 643 674 642 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01554 642 675 643 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01553 42 207 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01552 909 207 51 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01551 48 112 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01550 909 48 42 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01549 42 51 50 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01548 50 112 42 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01547 76 50 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01546 909 50 76 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01545 297 303 281 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01544 280 304 297 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01543 909 298 280 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01542 298 297 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01541 295 304 298 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01540 909 425 304 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01539 303 304 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01538 909 289 302 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01537 281 302 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01536 279 278 295 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01535 909 296 279 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01534 296 295 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01533 909 295 296 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01532 37 222 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01531 909 222 35 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01530 34 79 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01529 909 34 37 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01528 37 35 36 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01527 36 79 37 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01526 99 36 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01525 909 36 99 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01524 406 421 401 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01523 400 422 406 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01522 909 404 400 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01521 404 406 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01520 416 422 404 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01519 909 425 422 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01518 421 422 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01517 909 472 420 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01516 401 420 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01515 399 398 416 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01514 909 795 399 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01513 795 416 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01512 909 416 795 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01511 467 710 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01510 909 722 467 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01509 779 795 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01508 909 946 779 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01507 909 925 876 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01506 870 925 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01505 879 928 870 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01504 870 876 879 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01503 909 875 870 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01502 875 928 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01501 706 816 701 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01500 701 815 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01499 909 861 706 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01498 834 706 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01497 465 536 466 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01496 466 506 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01495 909 467 465 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01494 464 465 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01493 277 674 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01492 909 711 277 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01491 291 290 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01490 290 722 277 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01489 277 736 290 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01488 909 515 486 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01487 476 515 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01486 485 482 476 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01485 476 486 485 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01484 909 483 476 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01483 483 482 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01482 574 702 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01481 646 573 574 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01480 909 572 646 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01479 909 99 101 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01478 82 99 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01477 118 148 82 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01476 82 101 118 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01475 909 98 82 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01474 98 148 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01473 215 218 214 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01472 209 219 215 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01471 909 211 209 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01470 211 215 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01469 210 219 211 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01468 909 216 219 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01467 218 219 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01466 909 213 217 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01465 214 217 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01464 208 206 210 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01463 909 207 208 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01462 207 210 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01461 909 210 207 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01460 909 439 377 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01459 377 449 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01458 909 375 377 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01457 451 377 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01456 139 207 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01455 909 112 139 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01454 336 334 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01453 909 899 336 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01452 359 336 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01451 352 485 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01450 469 451 352 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01449 909 899 469 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01448 682 680 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01447 692 681 682 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01446 909 679 692 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01445 537 548 538 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01444 538 552 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01443 909 535 537 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01442 536 537 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01441 463 686 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01440 909 722 463 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01439 620 643 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01438 625 685 620 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01437 909 676 625 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01436 909 521 494 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01435 496 521 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01434 515 702 496 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01433 496 494 515 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01432 909 495 496 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01431 495 702 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01430 733 712 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01429 704 715 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01428 909 777 713 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01427 909 943 703 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01426 703 713 712 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01425 712 777 704 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01424 909 897 900 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01423 900 898 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01422 909 899 900 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01421 933 900 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01420 275 296 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01419 909 296 273 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01418 272 274 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01417 909 272 275 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01416 275 273 276 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01415 276 274 275 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01414 271 276 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01413 909 276 271 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01412 909 479 349 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01411 349 477 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01410 909 493 349 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01409 388 349 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01408 19 21 18 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01407 16 22 19 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01406 909 17 16 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01405 17 19 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01404 15 22 17 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01403 909 244 22 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01402 21 22 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01401 909 44 20 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01400 18 20 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01399 14 13 15 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01398 909 171 14 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01397 171 15 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01396 909 15 171 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01395 909 107 88 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01394 80 107 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01393 86 83 80 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01392 80 88 86 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01391 909 85 80 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01390 85 83 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01389 544 686 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01388 909 673 544 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01387 543 544 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01386 633 675 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01385 909 686 633 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01384 632 633 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01383 914 922 904 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01382 903 923 914 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01381 909 913 903 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01380 913 914 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01379 911 923 913 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01378 909 921 923 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01377 922 923 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01376 909 916 919 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01375 904 919 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01374 902 901 911 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01373 909 910 902 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01372 910 911 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01371 909 911 910 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01370 797 795 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01369 909 946 797 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01368 815 797 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01367 745 743 719 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01366 719 742 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01365 909 744 745 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01364 773 745 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01363 679 673 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01362 679 675 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01361 909 686 679 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01360 909 736 679 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01359 784 880 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01358 898 834 784 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01357 909 892 898 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01356 481 710 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01355 909 722 481 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01354 479 481 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01353 584 685 579 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01352 579 643 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01351 909 676 584 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01350 583 584 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01349 683 688 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01348 727 743 683 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01347 909 778 727 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01346 909 610 578 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01345 577 610 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01344 645 576 577 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01343 577 578 645 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01342 909 575 577 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01341 575 576 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01340 909 663 664 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01339 649 663 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01338 715 660 649 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01337 649 664 715 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01336 909 659 649 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01335 659 660 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01334 909 673 539 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01333 539 675 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01332 539 736 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01331 909 674 539 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01330 569 539 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01329 782 822 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01328 909 899 782 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01327 803 782 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01326 173 235 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01325 909 171 173 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01324 269 173 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01323 559 573 547 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01322 547 702 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01321 909 572 559 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01320 588 559 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01319 909 76 78 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01318 77 76 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01317 94 140 77 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01316 77 78 94 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01315 909 75 77 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01314 75 140 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01313 55 61 41 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01312 40 62 55 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01311 909 54 40 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01310 54 55 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01309 52 62 54 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01308 909 195 62 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01307 61 62 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01306 909 117 59 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01305 41 59 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01304 39 38 52 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01303 909 79 39 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01302 79 52 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01301 909 52 79 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01300 114 222 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01299 909 79 114 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01298 801 808 788 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01297 787 809 801 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01296 909 800 787 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01295 800 801 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01294 798 809 800 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01293 909 849 809 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01292 808 809 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01291 909 803 807 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01290 788 807 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01289 786 785 798 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01288 909 945 786 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01287 945 798 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01286 909 798 945 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01285 115 113 116 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01284 116 148 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01283 909 114 115 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01282 140 115 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01281 909 866 864 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01280 864 898 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01279 909 865 864 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01278 889 864 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01277 909 943 863 909 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_01276 861 868 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01275 863 862 868 909 sg13_lv_pmos L=0.13U W=2.27U AS=0.5448P AD=0.5448P PS=5.02U PD=5.02U 
Mtr_01274 268 267 270 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01273 270 269 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01272 909 379 268 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01271 816 268 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01270 553 569 545 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01269 545 643 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01268 909 685 553 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01267 552 553 909 909 sg13_lv_pmos L=0.13U W=2.34U AS=0.5616P AD=0.5616P PS=5.17U PD=5.17U 
Mtr_01266 391 464 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01265 390 388 391 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01264 909 389 390 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01263 897 942 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01262 897 879 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01261 909 867 897 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01260 909 526 523 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01259 501 526 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01258 541 543 501 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01257 501 523 541 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01256 909 522 501 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01255 522 543 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01254 647 645 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01253 909 646 647 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01252 817 815 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01251 867 816 817 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01250 909 861 867 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01249 542 541 909 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01248 909 583 542 909 sg13_lv_pmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_01247 573 542 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01246 909 645 591 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01245 580 645 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01244 663 588 580 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01243 580 591 663 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01242 909 589 580 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01241 589 588 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01240 899 777 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01239 680 675 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01238 143 171 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01237 895 925 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01236 909 925 894 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01235 893 928 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01234 909 893 895 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01233 895 894 896 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01232 896 928 895 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01231 892 896 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01230 909 896 892 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01229 909 370 371 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01228 365 370 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01227 374 463 365 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01226 365 371 374 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01225 909 367 365 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01224 367 463 909 909 sg13_lv_pmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_01223 772 775 770 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01222 771 776 772 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01221 909 769 771 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01220 769 772 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01219 768 776 769 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01218 909 921 776 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01217 775 776 909 909 sg13_lv_pmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_01216 909 773 774 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01215 770 774 909 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01214 767 766 768 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01213 909 792 767 909 sg13_lv_pmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01212 792 768 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01211 909 768 792 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01210 909 413 123 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01209 122 123 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01208 909 123 122 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01207 909 123 122 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01206 122 123 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01205 909 413 137 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01204 136 137 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01203 909 137 136 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01202 909 137 136 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01201 136 137 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01200 909 413 138 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01199 244 138 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01198 909 138 244 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01197 909 138 244 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01196 244 138 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01195 909 413 127 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01194 128 127 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01193 909 127 128 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01192 909 127 128 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01191 128 127 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01190 909 413 393 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01189 392 393 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01188 909 393 392 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01187 909 393 392 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01186 392 393 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01185 909 413 410 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01184 409 410 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01183 909 410 409 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01182 909 410 409 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01181 409 410 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01180 909 413 408 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01179 407 408 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01178 909 408 407 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01177 909 408 407 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01176 407 408 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01175 909 413 387 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01174 386 387 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01173 909 387 386 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01172 909 387 386 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01171 386 387 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01170 909 413 147 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01169 216 147 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01168 909 147 216 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01167 909 147 216 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01166 216 147 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01165 909 413 146 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01164 145 146 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01163 909 146 145 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01162 909 146 145 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01161 145 146 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01160 909 430 155 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01159 154 155 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01158 909 155 154 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01157 909 155 154 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01156 154 155 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01155 909 430 153 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01154 152 153 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01153 909 153 152 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01152 909 153 152 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01151 152 153 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01150 909 430 132 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01149 131 132 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01148 909 132 131 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01147 909 132 131 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01146 131 132 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01145 909 430 151 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01144 195 151 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01143 909 151 195 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01142 909 151 195 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01141 195 151 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01140 909 430 150 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01139 149 150 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01138 909 150 149 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01137 909 150 149 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01136 149 150 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01135 909 430 130 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01134 129 130 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01133 909 130 129 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01132 909 130 129 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01131 129 130 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01130 909 413 415 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01129 414 415 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01128 909 415 414 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01127 909 415 414 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01126 414 415 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01125 909 413 412 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01124 411 412 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01123 909 412 411 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01122 909 412 411 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01121 411 412 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01120 909 430 431 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01119 429 431 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01118 909 431 429 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01117 909 431 429 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01116 429 431 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01115 909 430 428 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01114 427 428 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01113 909 428 427 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01112 909 428 427 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01111 427 428 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01110 909 430 397 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01109 396 397 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01108 909 397 396 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01107 909 397 396 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01106 396 397 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01105 909 430 426 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01104 425 426 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01103 909 426 425 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01102 909 426 425 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01101 425 426 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01100 909 430 424 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01099 423 424 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01098 909 424 423 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01097 909 424 423 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01096 423 424 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01095 909 430 395 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01094 394 395 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01093 909 395 394 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01092 909 395 394 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01091 394 395 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01090 909 839 582 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01089 581 582 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01088 909 582 581 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01087 909 582 581 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01086 581 582 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01085 909 839 607 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01084 606 607 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01083 909 607 606 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01082 909 607 606 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01081 606 607 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01080 909 839 587 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01079 586 587 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01078 909 587 586 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01077 909 587 586 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01076 586 587 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01075 909 839 602 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01074 601 602 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01073 909 602 601 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01072 909 602 601 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01071 601 602 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01070 909 839 599 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01069 600 599 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01068 909 599 600 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01067 909 599 600 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01066 600 599 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01065 909 839 833 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01064 921 833 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01063 909 833 921 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01062 909 833 921 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01061 921 833 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01060 909 839 832 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01059 831 832 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01058 909 832 831 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01057 909 832 831 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01056 831 832 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01055 909 839 814 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01054 813 814 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01053 909 814 813 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01052 909 814 813 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01051 813 814 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01050 909 839 608 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01049 609 608 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01048 909 608 609 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01047 909 608 609 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01046 609 608 909 909 sg13_lv_pmos L=0.13U W=2.94U AS=0.7056P AD=0.7056P PS=6.37U PD=6.37U 
Mtr_01045 947 839 818 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01044 819 818 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01043 947 818 819 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01042 947 818 819 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01041 819 818 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01040 947 854 596 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01039 595 596 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01038 947 596 595 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01037 947 596 595 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01036 595 596 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01035 947 854 615 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01034 614 615 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01033 947 615 614 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01032 947 615 614 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01031 614 615 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01030 947 854 613 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01029 612 613 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01028 947 613 612 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01027 947 613 612 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01026 612 613 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01025 947 854 594 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01024 593 594 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01023 947 594 593 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01022 947 594 593 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01021 593 594 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01020 947 839 840 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01019 938 840 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01018 947 840 938 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01017 947 840 938 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01016 938 840 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01015 947 839 838 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01014 837 838 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01013 947 838 837 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01012 947 838 837 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01011 837 838 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01010 947 854 855 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01009 853 855 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01008 947 855 853 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01007 947 855 853 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01006 853 855 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01005 947 854 852 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01004 851 852 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01003 947 852 851 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01002 947 852 851 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01001 851 852 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_01000 947 854 828 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00999 827 828 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00998 947 828 827 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00997 947 828 827 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00996 827 828 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00995 947 854 850 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00994 849 850 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00993 947 850 849 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00992 947 850 849 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00991 849 850 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00990 947 854 848 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00989 847 848 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00988 947 848 847 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00987 947 848 847 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00986 847 848 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00985 947 854 826 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00984 825 826 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00983 947 826 825 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00982 947 826 825 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00981 825 826 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00980 947 854 619 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00979 618 619 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00978 947 619 618 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00977 947 619 618 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00976 618 619 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00975 947 854 617 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00974 616 617 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00973 947 617 616 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00972 947 617 616 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00971 616 617 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00970 947 899 46 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00969 46 86 45 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00968 44 45 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00967 448 477 450 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00966 450 479 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00965 449 493 448 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00964 947 694 305 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00963 430 305 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00962 947 305 430 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00961 947 305 430 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00960 430 305 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00959 947 694 292 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00958 413 292 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00957 947 292 413 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00956 947 292 413 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00955 413 292 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00954 383 795 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00953 947 795 384 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00952 947 946 380 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00951 382 381 383 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00950 380 384 382 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00949 379 382 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00948 947 382 379 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00947 381 946 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00946 213 169 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00945 947 777 170 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00944 168 325 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00943 169 170 168 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00942 167 777 169 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00941 947 207 167 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00940 504 736 505 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00939 505 673 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00938 503 711 504 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00937 502 674 503 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00936 176 177 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00935 947 176 178 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00934 178 183 177 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00933 177 184 181 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00932 947 216 184 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00931 183 184 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00930 947 179 182 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00929 181 180 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00928 174 183 176 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00927 175 184 174 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00926 947 222 175 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00925 222 174 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00924 947 174 222 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00923 731 734 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00922 947 731 732 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00921 732 735 734 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00920 734 756 755 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00919 947 849 756 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00918 735 756 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00917 947 757 758 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00916 755 754 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00915 753 735 731 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00914 730 756 753 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00913 947 943 730 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00912 943 753 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00911 947 753 943 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00910 435 777 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00909 471 795 435 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00908 605 603 597 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00907 597 631 605 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00906 947 647 597 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00905 677 605 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00904 221 223 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00903 947 777 226 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00902 203 248 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00901 223 226 203 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00900 202 777 223 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00899 947 222 202 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00898 332 379 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00897 947 379 333 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00896 334 331 332 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00895 330 333 334 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00894 947 329 330 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00893 331 329 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00892 944 943 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00891 942 945 944 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00890 516 515 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00889 947 515 512 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00888 556 511 516 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00887 514 512 556 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00886 947 513 514 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00885 511 513 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00884 238 242 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00883 947 238 239 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00882 239 245 242 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00881 242 247 243 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00880 947 244 247 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00879 245 247 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00878 947 240 246 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00877 243 241 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00876 236 245 238 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00875 237 247 236 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00874 947 235 237 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00873 235 236 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00872 947 236 235 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00871 684 686 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00870 685 711 684 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00869 947 899 105 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00868 105 118 119 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00867 117 119 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00866 166 235 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00865 252 171 166 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00864 650 652 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00863 651 673 652 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00862 947 736 651 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00861 653 674 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00860 652 675 653 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00859 947 235 197 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00858 197 777 205 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00857 262 205 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00856 447 463 446 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00855 446 445 447 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00854 947 502 446 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00853 535 447 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00852 947 674 312 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00851 312 722 316 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00850 315 316 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00849 439 506 433 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00848 433 536 439 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00847 947 467 433 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00846 373 374 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00845 389 372 373 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00844 890 889 883 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00843 883 888 890 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00842 947 899 883 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00841 916 890 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00840 947 928 926 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00839 926 925 927 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00838 924 927 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00837 666 675 667 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00836 667 710 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00835 665 686 666 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00834 690 673 665 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00833 320 736 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00832 319 711 320 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00831 341 390 342 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00830 342 555 351 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00829 947 899 341 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00828 350 351 947 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00827 73 140 65 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00826 65 72 73 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00825 947 139 65 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00824 83 73 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00823 72 112 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00822 947 207 72 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00821 113 79 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00820 947 222 113 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00819 251 124 947 947 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00818 125 139 124 947 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00817 124 220 126 947 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00816 126 143 947 947 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00815 947 140 125 947 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00814 125 141 947 947 sg13_lv_nmos L=0.13U W=2.12U AS=0.5088P AD=0.5088P PS=4.72U PD=4.72U 
Mtr_00813 947 497 498 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00812 694 498 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00811 947 498 694 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00810 947 498 694 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00809 694 498 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00808 947 694 695 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00807 854 695 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00806 947 695 854 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00805 947 695 854 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00804 854 695 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00803 947 694 687 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00802 839 687 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00801 947 687 839 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00800 947 687 839 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00799 839 687 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00798 551 676 550 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00797 550 622 549 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00796 947 650 551 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00795 548 549 947 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00794 947 945 882 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00793 882 943 881 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00792 880 881 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00791 947 780 821 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00790 780 779 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00789 821 816 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00788 520 540 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00787 947 540 517 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00786 521 519 520 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00785 518 517 521 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00784 947 583 518 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00783 519 583 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00782 657 675 658 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00781 658 710 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00780 656 686 657 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00779 742 655 947 947 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00778 655 654 656 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00777 873 924 874 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00776 874 871 873 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00775 947 872 874 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00774 888 873 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00773 947 899 96 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00772 96 94 95 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00771 93 95 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00770 477 552 478 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00769 478 548 477 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00768 947 535 478 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00767 744 777 699 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00766 947 792 705 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00765 699 705 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00764 947 677 671 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00763 671 691 678 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00762 688 678 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00761 947 711 623 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00760 623 686 624 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00759 622 624 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00758 947 451 452 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00757 452 485 453 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00756 470 453 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00755 947 321 249 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00754 249 291 250 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00753 248 250 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00752 27 30 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00751 947 27 7 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00750 7 31 30 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00749 30 33 6 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00748 947 216 33 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00747 31 33 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00746 947 8 32 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00745 6 12 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00744 26 31 27 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00743 5 33 26 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00742 947 112 5 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00741 112 26 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00740 947 26 112 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00739 931 936 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00738 947 931 932 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00737 932 939 936 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00736 936 941 937 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00735 947 938 941 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00734 939 941 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00733 947 934 940 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00732 937 935 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00731 929 939 931 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00730 930 941 929 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00729 947 928 930 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00728 928 929 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00727 947 929 928 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00726 947 252 254 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00725 254 251 253 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00724 329 253 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00723 134 143 947 947 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00722 267 220 134 947 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00721 133 139 267 947 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00720 947 140 133 947 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00719 133 141 947 947 sg13_lv_nmos L=0.13U W=1.97U AS=0.4728P AD=0.4728P PS=4.42U PD=4.42U 
Mtr_00718 571 643 564 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00717 564 569 571 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00716 947 685 564 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00715 947 736 436 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00714 436 675 442 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00713 526 442 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00712 947 372 328 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00711 328 374 327 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00710 375 327 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00709 743 691 637 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00708 637 677 743 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00707 947 899 637 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00706 266 265 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00705 265 263 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00704 947 350 265 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00703 135 296 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00702 148 274 135 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00701 763 777 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00700 778 925 763 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00699 835 880 836 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00698 836 834 835 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00697 947 892 836 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00696 871 835 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00695 630 645 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00694 947 645 627 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00693 631 629 630 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00692 628 627 631 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00691 947 646 628 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00690 629 646 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00689 508 568 509 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00688 509 571 510 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00687 947 507 508 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00686 506 510 947 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00685 558 555 557 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00684 557 556 558 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00683 947 603 557 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00682 660 558 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00681 740 792 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00680 947 792 738 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00679 947 910 739 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00678 741 737 740 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00677 739 738 741 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00676 866 741 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00675 947 741 866 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00674 737 910 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00673 91 207 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00672 947 207 92 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00671 141 89 91 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00670 90 92 141 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00669 947 112 90 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00668 89 112 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00667 187 189 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00666 947 187 190 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00665 190 193 189 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00664 189 196 191 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00663 947 195 196 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00662 193 196 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00661 947 192 194 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00660 191 188 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00659 186 193 187 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00658 185 196 186 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00657 947 274 185 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00656 274 186 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00655 947 186 274 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00654 693 692 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00653 691 690 693 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00652 356 361 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00651 947 356 345 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00650 345 363 361 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00649 361 364 347 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00648 947 425 364 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00647 363 364 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00646 947 346 362 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00645 347 358 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00644 354 363 356 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00643 344 364 354 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00642 947 946 344 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00641 946 354 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00640 947 354 946 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00639 812 841 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00638 947 841 824 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00637 822 820 812 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00636 811 824 822 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00635 947 821 811 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00634 820 821 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00633 947 674 306 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00632 306 673 314 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00631 313 314 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00630 681 710 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00629 220 235 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00628 472 469 461 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00627 461 470 472 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00626 947 471 461 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00625 844 943 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00624 947 943 846 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00623 947 945 843 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00622 845 842 844 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00621 843 846 845 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00620 841 845 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00619 947 845 841 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00618 842 945 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00617 456 526 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00616 947 526 457 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00615 540 454 456 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00614 455 457 540 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00613 947 474 455 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00612 454 474 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00611 561 710 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00610 576 673 561 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00609 669 673 670 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00608 670 675 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00607 668 736 669 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00606 676 674 668 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00605 440 467 434 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00604 434 536 440 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00603 947 493 434 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00602 482 440 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00601 310 449 311 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00600 311 439 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00599 555 375 310 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00598 64 313 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00597 947 313 71 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00596 370 69 64 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00595 63 71 370 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00594 947 319 63 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00593 69 319 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00592 724 726 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00591 947 724 725 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00590 725 728 726 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00589 726 750 749 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00588 947 938 750 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00587 728 750 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00586 947 751 752 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00585 749 748 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00584 747 728 724 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00583 723 750 747 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00582 947 925 723 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00581 925 747 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00580 947 747 925 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00579 324 374 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00578 947 374 326 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00577 325 322 324 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00576 323 326 325 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00575 947 321 323 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00574 322 321 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00573 532 540 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00572 572 625 532 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00571 492 515 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00570 603 513 492 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00569 507 463 432 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00568 432 445 507 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00567 947 502 432 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00566 285 711 286 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00565 286 736 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00564 284 722 285 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00563 372 293 947 947 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00562 293 294 284 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00561 513 467 460 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00560 460 536 513 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00559 947 493 460 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00558 309 711 308 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00557 308 736 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00556 307 722 309 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00555 321 674 307 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00554 488 568 489 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00553 489 571 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00552 493 507 488 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00551 562 676 563 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00550 563 622 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00549 568 650 562 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00548 791 792 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00547 947 792 793 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00546 872 790 791 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00545 789 793 872 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00544 947 910 789 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00543 790 910 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00542 103 235 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00541 947 235 109 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00540 947 171 102 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00539 110 108 103 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00538 102 109 110 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00537 107 110 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00536 947 110 107 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00535 108 171 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00534 462 686 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00533 474 673 462 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00532 700 710 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00531 702 711 700 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00530 860 925 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00529 865 928 860 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00528 947 736 337 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00527 337 711 445 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00526 338 674 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00525 445 673 338 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00524 947 899 204 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00523 204 271 228 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00522 227 228 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00521 947 679 598 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00520 598 632 611 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00519 610 611 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00518 289 257 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00517 947 777 258 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00516 256 315 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00515 257 258 256 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00514 255 777 257 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00513 947 296 255 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00512 947 673 635 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00511 635 736 643 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00510 636 674 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00509 643 675 636 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00508 49 207 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00507 947 207 51 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00506 947 112 47 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00505 50 48 49 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00504 47 51 50 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00503 76 50 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00502 947 50 76 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00501 48 112 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00500 298 297 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00499 947 298 288 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00498 288 303 297 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00497 297 304 299 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00496 947 425 304 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00495 303 304 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00494 947 300 302 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00493 299 301 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00492 295 303 298 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00491 287 304 295 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00490 947 296 287 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00489 296 295 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00488 947 295 296 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00487 10 222 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00486 947 222 35 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00485 947 79 9 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00484 36 34 10 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00483 9 35 36 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00482 99 36 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00481 947 36 99 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00480 34 79 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00479 404 406 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00478 947 404 405 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00477 405 421 406 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00476 406 422 418 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00475 947 425 422 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00474 421 422 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00473 947 419 420 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00472 418 417 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00471 416 421 404 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00470 403 422 416 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00469 947 795 403 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00468 795 416 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00467 947 416 795 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00466 402 710 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00465 467 722 402 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00464 729 795 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00463 779 946 729 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00462 878 925 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00461 947 925 876 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00460 879 875 878 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00459 877 876 879 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00458 947 928 877 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00457 875 928 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00456 706 815 696 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00455 696 816 706 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00454 947 861 696 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00453 834 706 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00452 465 506 459 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00451 459 536 465 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00450 947 467 459 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00449 464 465 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00448 291 290 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00447 282 711 290 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00446 947 674 282 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00445 283 722 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00444 290 736 283 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00443 487 515 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00442 947 515 486 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00441 485 483 487 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00440 484 486 485 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00439 947 482 484 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00438 483 482 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00437 646 702 565 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00436 565 573 646 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00435 947 572 565 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00434 100 99 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00433 947 99 101 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00432 118 98 100 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00431 97 101 118 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00430 947 148 97 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00429 98 148 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00428 211 215 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00427 947 211 199 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00426 199 218 215 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00425 215 219 201 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00424 947 216 219 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00423 218 219 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00422 947 200 217 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00421 201 212 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00420 210 218 211 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00419 198 219 210 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00418 947 207 198 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00417 207 210 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00416 947 210 207 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00415 376 449 378 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00414 378 439 377 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00413 947 375 376 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00412 451 377 947 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00411 106 207 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00410 139 112 106 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00409 947 899 335 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00408 335 334 336 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00407 359 336 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00406 469 485 343 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00405 343 451 469 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00404 947 899 343 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00403 692 680 672 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00402 672 681 692 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00401 947 679 672 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00400 537 552 527 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00399 527 548 537 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00398 947 535 527 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00397 536 537 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00396 458 686 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00395 463 722 458 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00394 625 643 626 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00393 626 685 625 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00392 947 676 626 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00391 491 521 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00390 947 521 494 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00389 515 495 491 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00388 490 494 515 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00387 947 702 490 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00386 495 702 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00385 733 712 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00384 947 777 713 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00383 698 715 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00382 712 713 698 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00381 697 777 712 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00380 947 943 697 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00379 886 898 887 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00378 887 897 900 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00377 947 899 886 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00376 933 900 947 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00375 261 296 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00374 947 296 273 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00373 947 274 260 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00372 276 272 261 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00371 260 273 276 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00370 271 276 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00369 947 276 271 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00368 272 274 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00367 339 477 340 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00366 340 479 349 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00365 947 493 339 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00364 388 349 947 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00363 17 19 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00362 947 17 2 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00361 2 21 19 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00360 19 22 4 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00359 947 244 22 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00358 21 22 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00357 947 3 20 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00356 4 11 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00355 15 21 17 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00354 1 22 15 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00353 947 171 1 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00352 171 15 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00351 947 15 171 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00350 87 107 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00349 947 107 88 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00348 86 85 87 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00347 84 88 86 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00346 947 83 84 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00345 85 83 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00344 947 673 534 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00343 534 686 544 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00342 543 544 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00341 947 686 634 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00340 634 675 633 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00339 632 633 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00338 913 914 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00337 947 913 915 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00336 915 922 914 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00335 914 923 920 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00334 947 921 923 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00333 922 923 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00332 947 917 919 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00331 920 918 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00330 911 922 913 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00329 912 923 911 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00328 947 910 912 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00327 910 911 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00326 947 911 910 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00325 947 946 796 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00324 796 795 797 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00323 815 797 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00322 745 742 746 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00321 746 743 745 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00320 947 744 746 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00319 773 745 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00318 641 686 640 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00317 640 675 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00316 639 673 641 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00315 679 736 639 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00314 898 880 794 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00313 794 834 898 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00312 947 892 794 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00311 947 722 480 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00310 480 710 481 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00309 479 481 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00308 584 643 585 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00307 585 685 584 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00306 947 676 585 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00305 583 584 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00304 727 688 689 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00303 689 743 727 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00302 947 778 689 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00301 567 610 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00300 947 610 578 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00299 645 575 567 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00298 566 578 645 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00297 947 576 566 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00296 575 576 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00295 662 663 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00294 947 663 664 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00293 715 659 662 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00292 661 664 715 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00291 947 660 661 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00290 659 660 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00289 530 673 531 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00288 531 675 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00287 529 736 530 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00286 569 539 947 947 sg13_lv_nmos L=0.13U W=1.89U AS=0.4536P AD=0.4536P PS=4.27U PD=4.27U 
Mtr_00285 539 528 529 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00284 947 899 764 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00283 764 822 782 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00282 803 782 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00281 947 171 172 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00280 172 235 173 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00279 269 173 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00278 559 702 560 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00277 560 573 559 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00276 947 572 560 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00275 588 559 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00274 67 76 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00273 947 76 78 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00272 94 75 67 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00271 66 78 94 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00270 947 140 66 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00269 75 140 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00268 54 55 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00267 947 54 56 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00266 56 61 55 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00265 55 62 60 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00264 947 195 62 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00263 61 62 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00262 947 57 59 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00261 60 58 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00260 52 61 54 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00259 53 62 52 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00258 947 79 53 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00257 79 52 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00256 947 52 79 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00255 68 222 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00254 114 79 68 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00253 800 801 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00252 947 800 802 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00251 802 808 801 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00250 801 809 806 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00249 947 849 809 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00248 808 809 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00247 947 804 807 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00246 806 805 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00245 798 808 800 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00244 799 809 798 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00243 947 945 799 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00242 945 798 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00241 947 798 945 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00240 115 148 104 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00239 104 113 115 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00238 947 114 104 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00237 140 115 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00236 859 898 858 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00235 858 866 864 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00234 947 865 859 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00233 889 864 947 947 sg13_lv_nmos L=0.13U W=2.19U AS=0.5256P AD=0.5256P PS=4.87U PD=4.87U 
Mtr_00232 861 868 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00231 868 862 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00230 947 943 868 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00229 268 269 259 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00228 259 267 268 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00227 947 379 259 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00226 816 268 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00225 553 643 554 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00224 554 569 553 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00223 947 685 554 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00222 552 553 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00221 390 464 385 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00220 385 388 390 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00219 947 389 385 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00218 857 867 856 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00217 856 879 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00216 897 942 857 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00215 525 526 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00214 947 526 523 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00213 541 522 525 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00212 524 523 541 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00211 947 543 524 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00210 522 543 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00209 638 645 947 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00208 647 646 638 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00207 867 815 810 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00206 810 816 867 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00205 947 861 810 947 sg13_lv_nmos L=0.13U W=1.52U AS=0.3648P AD=0.3648P PS=3.52U PD=3.52U 
Mtr_00204 947 583 533 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00203 533 541 542 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00202 573 542 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00201 592 645 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00200 947 645 591 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00199 663 589 592 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00198 590 591 663 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00197 947 588 590 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00196 589 588 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00195 899 777 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00194 680 675 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00193 143 171 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00192 884 925 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00191 947 925 894 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00190 947 928 885 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00189 896 893 884 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00188 885 894 896 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00187 892 896 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00186 947 896 892 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00185 893 928 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00184 369 370 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00183 947 370 371 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00182 374 367 369 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00181 368 371 374 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00180 947 463 368 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00179 367 463 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00178 769 772 947 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00177 947 769 761 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00176 761 775 772 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00175 772 776 760 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00174 947 921 776 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00173 775 776 947 947 sg13_lv_nmos L=0.13U W=1.07U AS=0.2568P AD=0.2568P PS=2.62U PD=2.62U 
Mtr_00172 947 762 774 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00171 760 765 947 947 sg13_lv_nmos L=0.13U W=1.37U AS=0.3288P AD=0.3288P PS=3.22U PD=3.22U 
Mtr_00170 768 775 769 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00169 759 776 768 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00168 947 792 759 947 sg13_lv_nmos L=0.13U W=0.77U AS=0.1848P AD=0.1848P PS=2.02U PD=2.02U 
Mtr_00167 792 768 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00166 947 768 792 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00165 947 413 123 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00164 122 123 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00163 947 123 122 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00162 947 123 122 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00161 122 123 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00160 947 413 137 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00159 136 137 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00158 947 137 136 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00157 947 137 136 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00156 136 137 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00155 947 413 138 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00154 244 138 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00153 947 138 244 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00152 947 138 244 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00151 244 138 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00150 947 413 127 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00149 128 127 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00148 947 127 128 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00147 947 127 128 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00146 128 127 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00145 947 413 393 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00144 392 393 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00143 947 393 392 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00142 947 393 392 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00141 392 393 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00140 947 413 410 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00139 409 410 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00138 947 410 409 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00137 947 410 409 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00136 409 410 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00135 947 413 408 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00134 407 408 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00133 947 408 407 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00132 947 408 407 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00131 407 408 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00130 947 413 387 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00129 386 387 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00128 947 387 386 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00127 947 387 386 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00126 386 387 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00125 947 413 147 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00124 216 147 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00123 947 147 216 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00122 947 147 216 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00121 216 147 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00120 947 413 146 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00119 145 146 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00118 947 146 145 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00117 947 146 145 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00116 145 146 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00115 947 430 155 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00114 154 155 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00113 947 155 154 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00112 947 155 154 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00111 154 155 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00110 947 430 153 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00109 152 153 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00108 947 153 152 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00107 947 153 152 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00106 152 153 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00105 947 430 132 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00104 131 132 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00103 947 132 131 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00102 947 132 131 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00101 131 132 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00100 947 430 151 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00099 195 151 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00098 947 151 195 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00097 947 151 195 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00096 195 151 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00095 947 430 150 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00094 149 150 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00093 947 150 149 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00092 947 150 149 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00091 149 150 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00090 947 430 130 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00089 129 130 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00088 947 130 129 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00087 947 130 129 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00086 129 130 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00085 947 413 415 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00084 414 415 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00083 947 415 414 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00082 947 415 414 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00081 414 415 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00080 947 413 412 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00079 411 412 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00078 947 412 411 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00077 947 412 411 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00076 411 412 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00075 947 430 431 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00074 429 431 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00073 947 431 429 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00072 947 431 429 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00071 429 431 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00070 947 430 428 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00069 427 428 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00068 947 428 427 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00067 947 428 427 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00066 427 428 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00065 947 430 397 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00064 396 397 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00063 947 397 396 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00062 947 397 396 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00061 396 397 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00060 947 430 426 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00059 425 426 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00058 947 426 425 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00057 947 426 425 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00056 425 426 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00055 947 430 424 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00054 423 424 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00053 947 424 423 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00052 947 424 423 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00051 423 424 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00050 947 430 395 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00049 394 395 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00048 947 395 394 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00047 947 395 394 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00046 394 395 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00045 947 839 582 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00044 581 582 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00043 947 582 581 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00042 947 582 581 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00041 581 582 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00040 947 839 607 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00039 606 607 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00038 947 607 606 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00037 947 607 606 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00036 606 607 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00035 947 839 587 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00034 586 587 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00033 947 587 586 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00032 947 587 586 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00031 586 587 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00030 947 839 602 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00029 601 602 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00028 947 602 601 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00027 947 602 601 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00026 601 602 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00025 947 839 599 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00024 600 599 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00023 947 599 600 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00022 947 599 600 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00021 600 599 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00020 947 839 833 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00019 921 833 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00018 947 833 921 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00017 947 833 921 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00016 921 833 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00015 947 839 832 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00014 831 832 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00013 947 832 831 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00012 947 832 831 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00011 831 832 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00010 947 839 814 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00009 813 814 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00008 947 814 813 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00007 947 814 813 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00006 813 814 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00005 947 839 608 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00004 609 608 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00003 947 608 609 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00002 947 608 609 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00001 609 608 947 947 sg13_lv_nmos L=0.13U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C988 3 947 2.46362e-15
C983 8 947 2.46362e-15
C979 11 947 9.91138e-15
C978 12 947 9.91138e-15
C977 13 947 5.27918e-15
C975 15 947 3.38702e-14
C973 17 947 2.08974e-14
C971 19 947 1.89138e-14
C970 20 947 1.54958e-14
C969 21 947 6.90483e-14
C968 22 947 9.52956e-14
C965 25 947 5.27918e-15
C964 26 947 3.38702e-14
C963 27 947 2.08974e-14
C960 30 947 1.89138e-14
C959 31 947 6.90483e-14
C958 32 947 1.54958e-14
C957 33 947 9.52956e-14
C956 34 947 3.09307e-14
C955 35 947 2.81118e-14
C954 36 947 3.4793e-14
C953 37 947 1.14176e-15
C952 38 947 5.27918e-15
C948 42 947 1.14176e-15
C945 44 947 1.50518e-14
C944 45 947 2.16616e-14
C941 48 947 3.09307e-14
C939 50 947 3.4793e-14
C938 51 947 2.81118e-14
C937 52 947 3.38702e-14
C935 54 947 2.08974e-14
C934 55 947 1.89138e-14
C932 57 947 2.46362e-15
C931 58 947 9.91138e-15
C930 59 947 1.54958e-14
C928 61 947 6.90483e-14
C927 62 947 9.52956e-14
C924 65 947 4.17738e-16
C919 69 947 2.7614e-14
C918 70 947 8.63047e-16
C917 71 947 2.86016e-14
C916 72 947 2.24388e-14
C915 73 947 3.01232e-14
C913 75 947 2.7614e-14
C912 76 947 3.2062e-14
C911 77 947 8.63047e-16
C910 78 947 2.86016e-14
C909 79 947 1.13069e-13
C908 80 947 8.63047e-16
C907 81 947 8.63047e-16
C906 82 947 8.63047e-16
C904 83 947 4.19639e-14
C902 85 947 2.7614e-14
C901 86 947 2.51577e-14
C899 88 947 2.86016e-14
C898 89 947 2.7614e-14
C895 92 947 2.86016e-14
C894 93 947 1.73203e-14
C893 94 947 2.42991e-14
C892 95 947 2.16616e-14
C889 98 947 2.7614e-14
C888 99 947 3.31691e-14
C886 101 947 2.86016e-14
C883 104 947 4.17738e-16
C879 107 947 3.10163e-14
C878 108 947 3.09307e-14
C877 109 947 2.81118e-14
C876 110 947 3.4793e-14
C875 111 947 1.14176e-15
C874 112 947 1.47551e-13
C873 113 947 2.39129e-14
C872 114 947 2.67162e-14
C871 115 947 3.01232e-14
C869 117 947 1.73203e-14
C868 118 947 2.54386e-14
C867 119 947 2.16616e-14
C865 121 947 9.28968e-16
C863 122 947 3.29763e-15
C862 123 947 8.3284e-14
C861 124 947 1.20682e-14
C860 125 947 4.45309e-16
C858 127 947 8.3284e-14
C857 128 947 3.29763e-15
C856 129 947 3.29763e-15
C855 130 947 8.3284e-14
C854 131 947 3.29763e-15
C853 132 947 8.3284e-14
C852 133 947 4.45309e-16
C848 136 947 3.29763e-15
C847 137 947 8.3284e-14
C846 138 947 8.3284e-14
C845 139 947 6.5526e-14
C844 140 947 1.08872e-13
C843 141 947 4.12192e-14
C841 143 947 3.38749e-14
C840 144 947 9.70324e-16
C839 145 947 3.29763e-15
C838 146 947 8.3284e-14
C837 147 947 8.3284e-14
C836 148 947 6.05503e-14
C835 149 947 3.29763e-15
C834 150 947 8.3284e-14
C833 151 947 8.3284e-14
C832 152 947 3.29763e-15
C831 153 947 8.3284e-14
C830 154 947 3.29763e-15
C829 155 947 8.3284e-14
C826 158 947 5.27918e-15
C821 163 947 5.27918e-15
C814 169 947 2.45636e-14
C813 170 947 1.82808e-14
C812 171 947 1.51371e-13
C810 173 947 2.16616e-14
C809 174 947 3.38702e-14
C807 176 947 2.08974e-14
C806 177 947 1.89138e-14
C804 179 947 2.46362e-15
C803 180 947 9.91138e-15
C801 182 947 1.54958e-14
C800 183 947 6.90483e-14
C799 184 947 9.52956e-14
C797 186 947 3.38702e-14
C796 187 947 2.08974e-14
C795 188 947 9.91138e-15
C794 189 947 1.89138e-14
C791 192 947 2.46362e-15
C790 193 947 6.90483e-14
C789 194 947 1.54958e-14
C788 195 947 4.21121e-14
C787 196 947 9.52956e-14
C783 200 947 2.46362e-15
C777 205 947 2.16616e-14
C776 206 947 5.27918e-15
C775 207 947 1.59704e-13
C772 210 947 3.38702e-14
C771 211 947 2.08974e-14
C770 212 947 9.91138e-15
C769 213 947 1.56996e-14
C767 215 947 1.89138e-14
C766 216 947 7.44141e-14
C765 217 947 1.54958e-14
C764 218 947 6.90483e-14
C763 219 947 9.52956e-14
C762 220 947 3.94905e-14
C761 221 947 1.55543e-14
C760 222 947 1.3363e-13
C759 223 947 2.45636e-14
C756 226 947 1.82808e-14
C755 227 947 1.50518e-14
C754 228 947 2.16616e-14
C748 234 947 5.27918e-15
C746 235 947 1.54329e-13
C745 236 947 3.38702e-14
C743 238 947 2.08974e-14
C741 240 947 2.46362e-15
C740 241 947 9.91138e-15
C739 242 947 1.89138e-14
C737 244 947 4.54013e-14
C736 245 947 6.90483e-14
C735 246 947 1.54958e-14
C734 247 947 9.52956e-14
C733 248 947 3.75825e-14
C731 250 947 2.16616e-14
C730 251 947 2.95166e-14
C729 252 947 3.48864e-14
C728 253 947 2.16616e-14
C724 257 947 2.45636e-14
C723 258 947 1.82808e-14
C722 259 947 4.17738e-16
C718 262 947 1.34751e-14
C717 263 947 1.09103e-14
C715 265 947 2.09836e-14
C714 266 947 1.5107e-14
C713 267 947 2.70926e-14
C712 268 947 3.01232e-14
C711 269 947 2.51078e-14
C709 271 947 2.48955e-14
C708 272 947 3.09307e-14
C707 273 947 2.81118e-14
C706 274 947 1.03766e-13
C705 275 947 1.14176e-15
C704 276 947 3.4793e-14
C703 277 947 8.87611e-16
C702 278 947 5.27918e-15
C690 289 947 1.75671e-14
C689 290 947 2.06663e-14
C688 291 947 2.7303e-14
C687 292 947 8.3284e-14
C686 293 947 1.80612e-14
C685 294 947 2.11167e-15
C684 295 947 3.38702e-14
C683 296 947 1.03956e-13
C682 297 947 1.89138e-14
C681 298 947 2.08974e-14
C679 300 947 2.46362e-15
C678 301 947 9.91138e-15
C677 302 947 1.54958e-14
C676 303 947 6.90483e-14
C675 304 947 9.52956e-14
C674 305 947 8.3284e-14
C665 313 947 4.05664e-14
C664 314 947 2.16616e-14
C663 315 947 2.91428e-14
C662 316 947 2.16616e-14
C661 317 947 8.63047e-16
C660 318 947 8.63047e-16
C658 319 947 4.57429e-14
C656 321 947 5.56891e-14
C655 322 947 2.7614e-14
C652 325 947 2.90183e-14
C651 326 947 2.86016e-14
C650 327 947 2.16616e-14
C648 329 947 4.46532e-14
C646 331 947 2.7614e-14
C644 333 947 2.86016e-14
C643 334 947 3.03745e-14
C641 336 947 2.16616e-14
C634 343 947 3.90167e-16
C631 346 947 2.46362e-15
C628 348 947 8.6004e-16
C627 349 947 1.44675e-14
C626 350 947 3.67578e-14
C625 351 947 1.44675e-14
C623 353 947 5.27918e-15
C622 354 947 3.38702e-14
C620 356 947 2.08974e-14
C618 358 947 9.91138e-15
C617 359 947 1.50518e-14
C615 361 947 1.89138e-14
C614 362 947 1.54958e-14
C613 363 947 6.90483e-14
C612 364 947 9.52956e-14
C611 365 947 8.63047e-16
C610 366 947 1.14176e-15
C608 367 947 2.7614e-14
C605 370 947 4.40448e-14
C604 371 947 2.86016e-14
C603 372 947 5.36932e-14
C601 374 947 9.19237e-14
C600 375 947 4.30792e-14
C598 377 947 1.44675e-14
C596 379 947 6.25406e-14
C594 381 947 3.09307e-14
C593 382 947 3.4793e-14
C591 384 947 2.81118e-14
C590 385 947 3.90167e-16
C588 386 947 3.29763e-15
C587 387 947 8.3284e-14
C586 388 947 2.16395e-14
C585 389 947 2.57931e-14
C584 390 947 2.77074e-14
C582 392 947 3.29763e-15
C581 393 947 8.3284e-14
C580 394 947 3.29763e-15
C579 395 947 8.3284e-14
C578 396 947 3.29763e-15
C577 397 947 8.3284e-14
C576 398 947 5.27918e-15
C569 404 947 2.08974e-14
C567 406 947 1.89138e-14
C566 407 947 3.29763e-15
C565 408 947 8.3284e-14
C564 409 947 3.29763e-15
C563 410 947 8.3284e-14
C562 411 947 3.29763e-15
C561 412 947 8.3284e-14
C560 413 947 2.96515e-13
C559 414 947 3.29763e-15
C558 415 947 8.3284e-14
C557 416 947 3.38702e-14
C556 417 947 9.91138e-15
C554 419 947 2.46362e-15
C553 420 947 1.54958e-14
C552 421 947 6.90483e-14
C551 422 947 9.52956e-14
C550 423 947 3.29763e-15
C549 424 947 8.3284e-14
C548 425 947 6.66248e-14
C547 426 947 8.3284e-14
C546 427 947 3.29763e-15
C545 428 947 8.3284e-14
C544 429 947 3.29763e-15
C543 430 947 2.96515e-13
C542 431 947 8.3284e-14
C541 432 947 3.90167e-16
C540 433 947 3.90167e-16
C539 434 947 4.17738e-16
C533 439 947 5.31374e-14
C532 440 947 3.01232e-14
C530 442 947 2.16616e-14
C528 444 947 8.63047e-16
C526 445 947 4.23983e-14
C525 446 947 4.17738e-16
C524 447 947 3.01232e-14
C522 449 947 5.38504e-14
C520 451 947 4.75727e-14
C518 453 947 2.16616e-14
C517 454 947 2.7614e-14
C514 457 947 2.86016e-14
C512 459 947 4.17738e-16
C511 460 947 3.90167e-16
C510 461 947 3.90167e-16
C507 463 947 7.34498e-14
C506 464 947 2.32971e-14
C505 465 947 3.01232e-14
C503 467 947 9.39746e-14
C501 469 947 2.43005e-14
C500 470 947 1.92332e-14
C499 471 947 2.7186e-14
C498 472 947 1.89001e-14
C496 474 947 3.51442e-14
C494 476 947 8.63047e-16
C492 477 947 5.80619e-14
C491 478 947 3.90167e-16
C490 479 947 4.68075e-14
C488 481 947 2.16616e-14
C487 482 947 4.16363e-14
C486 483 947 2.7614e-14
C484 485 947 4.98947e-14
C483 486 947 2.86016e-14
C475 493 947 1.02718e-13
C474 494 947 2.86016e-14
C473 495 947 2.7614e-14
C472 496 947 8.63047e-16
C471 497 947 6.29609e-14
C470 498 947 8.3284e-14
C469 499 947 8.63047e-16
C468 500 947 8.63047e-16
C467 501 947 8.63047e-16
C465 502 947 5.44453e-14
C461 506 947 4.1961e-14
C460 507 947 5.14842e-14
C457 510 947 1.44675e-14
C456 511 947 2.7614e-14
C455 512 947 2.86016e-14
C454 513 947 6.20098e-14
C452 515 947 8.86749e-14
C450 517 947 2.86016e-14
C448 519 947 2.7614e-14
C446 521 947 3.14281e-14
C445 522 947 2.7614e-14
C444 523 947 2.86016e-14
C441 526 947 6.23462e-14
C440 527 947 4.17738e-16
C439 528 947 2.11167e-15
C431 535 947 5.33812e-14
C430 536 947 9.36486e-14
C429 537 947 3.01232e-14
C427 539 947 1.80612e-14
C426 540 947 7.13107e-14
C425 541 947 3.01512e-14
C424 542 947 2.16616e-14
C423 543 947 3.54752e-14
C422 544 947 2.16616e-14
C417 548 947 4.19791e-14
C416 549 947 1.44675e-14
C413 552 947 4.60242e-14
C412 553 947 3.01232e-14
C411 554 947 4.17738e-16
C410 555 947 5.09564e-14
C409 556 947 2.18774e-14
C408 557 947 4.17738e-16
C407 558 947 3.01232e-14
C406 559 947 3.01232e-14
C405 560 947 4.17738e-16
C401 564 947 3.90167e-16
C400 565 947 3.90167e-16
C396 568 947 5.14589e-14
C395 569 947 3.8891e-14
C393 571 947 4.27053e-14
C392 572 947 5.45125e-14
C391 573 947 3.99692e-14
C389 575 947 2.7614e-14
C388 576 947 3.59142e-14
C387 577 947 8.63047e-16
C386 578 947 2.86016e-14
C384 580 947 8.63047e-16
C382 581 947 3.29763e-15
C381 582 947 8.3284e-14
C380 583 947 6.883e-14
C379 584 947 3.01232e-14
C378 585 947 4.17738e-16
C377 586 947 3.29763e-15
C376 587 947 8.3284e-14
C375 588 947 3.65764e-14
C374 589 947 2.7614e-14
C372 591 947 2.86016e-14
C370 593 947 3.29763e-15
C369 594 947 8.3284e-14
C368 595 947 3.29763e-15
C367 596 947 8.3284e-14
C366 597 947 4.17738e-16
C363 599 947 8.3284e-14
C362 600 947 3.29763e-15
C361 601 947 3.29763e-15
C360 602 947 8.3284e-14
C359 603 947 4.92824e-14
C357 605 947 3.01232e-14
C356 606 947 3.29763e-15
C355 607 947 8.3284e-14
C354 608 947 8.3284e-14
C353 609 947 3.29763e-15
C352 610 947 3.16229e-14
C351 611 947 2.16616e-14
C350 612 947 3.29763e-15
C349 613 947 8.3284e-14
C348 614 947 3.29763e-15
C347 615 947 8.3284e-14
C346 616 947 3.29763e-15
C345 617 947 8.3284e-14
C344 618 947 3.29763e-15
C343 619 947 8.3284e-14
C341 621 947 8.63047e-16
C339 622 947 4.12707e-14
C337 624 947 2.16616e-14
C336 625 947 3.81612e-14
C335 626 947 3.90167e-16
C334 627 947 2.86016e-14
C332 629 947 2.7614e-14
C330 631 947 2.84837e-14
C329 632 947 2.37061e-14
C328 633 947 2.16616e-14
C324 637 947 3.90167e-16
C318 642 947 8.6004e-16
C317 643 947 7.96787e-14
C315 645 947 9.18419e-14
C314 646 947 6.20532e-14
C313 647 947 3.2977e-14
C312 648 947 8.87611e-16
C311 649 947 8.63047e-16
C309 650 947 4.5463e-14
C307 652 947 2.06663e-14
C305 654 947 2.11167e-15
C304 655 947 1.80612e-14
C300 659 947 2.7614e-14
C299 660 947 4.16351e-14
C296 663 947 3.99518e-14
C295 664 947 2.86016e-14
C287 672 947 3.90167e-16
C285 673 947 3.41716e-13
C284 674 947 2.79812e-13
C283 675 947 2.79202e-13
C282 676 947 1.0251e-13
C281 677 947 4.22667e-14
C280 678 947 2.16616e-14
C279 679 947 4.63057e-14
C278 680 947 1.96687e-14
C277 681 947 2.63181e-14
C272 685 947 9.45275e-14
C271 686 947 2.67781e-13
C270 687 947 8.3284e-14
C269 688 947 1.80608e-14
C268 689 947 3.90167e-16
C267 690 947 2.81736e-14
C266 691 947 5.10565e-14
C265 692 947 3.05164e-14
C263 694 947 1.57555e-13
C262 695 947 8.3284e-14
C261 696 947 4.17738e-16
C254 702 947 8.26615e-14
C251 705 947 2.0721e-14
C250 706 947 3.01232e-14
C246 710 947 2.36525e-13
C245 711 947 2.60655e-13
C244 712 947 2.45636e-14
C243 713 947 1.82808e-14
C241 715 947 3.81028e-14
C238 718 947 1.14176e-15
C236 720 947 5.27918e-15
C235 721 947 5.27918e-15
C233 722 947 2.09984e-13
C231 724 947 2.08974e-14
C229 726 947 1.89138e-14
C228 727 947 1.72441e-14
C227 728 947 6.90483e-14
C224 731 947 2.08974e-14
C222 733 947 1.65463e-14
C221 734 947 1.89138e-14
C220 735 947 6.90483e-14
C219 736 947 3.51036e-13
C218 737 947 3.09307e-14
C217 738 947 2.81118e-14
C214 741 947 3.4793e-14
C213 742 947 2.46171e-14
C212 743 947 4.95701e-14
C211 744 947 2.54997e-14
C210 745 947 3.01232e-14
C209 746 947 4.17738e-16
C208 747 947 3.38702e-14
C207 748 947 9.91138e-15
C205 750 947 9.52956e-14
C204 751 947 2.46362e-15
C203 752 947 1.54958e-14
C202 753 947 3.38702e-14
C201 754 947 9.91138e-15
C199 756 947 9.52956e-14
C198 757 947 2.46362e-15
C197 758 947 1.54958e-14
C193 762 947 2.46362e-15
C189 765 947 9.91138e-15
C188 766 947 5.27918e-15
C186 768 947 3.38702e-14
C185 769 947 2.08974e-14
C182 772 947 1.89138e-14
C181 773 947 1.58442e-14
C180 774 947 1.54958e-14
C179 775 947 6.90483e-14
C178 776 947 9.52956e-14
C177 777 947 4.87759e-13
C176 778 947 2.88397e-14
C175 779 947 1.82049e-14
C174 780 947 2.12482e-14
C172 782 947 2.16616e-14
C171 783 947 8.63047e-16
C169 785 947 5.27918e-15
C163 790 947 2.7614e-14
C161 792 947 1.01618e-13
C160 793 947 2.86016e-14
C159 794 947 3.90167e-16
C158 795 947 1.44867e-13
C156 797 947 2.16616e-14
C155 798 947 3.38702e-14
C153 800 947 2.08974e-14
C152 801 947 1.89138e-14
C150 803 947 1.50518e-14
C149 804 947 2.46362e-15
C148 805 947 9.91138e-15
C146 807 947 1.54958e-14
C145 808 947 6.90483e-14
C144 809 947 9.52956e-14
C143 810 947 3.90167e-16
C139 813 947 3.29763e-15
C138 814 947 8.3284e-14
C137 815 947 4.8422e-14
C136 816 947 9.55827e-14
C134 818 947 8.3284e-14
C133 819 947 3.29763e-15
C132 820 947 2.7614e-14
C131 821 947 3.98933e-14
C130 822 947 2.73746e-14
C129 823 947 8.63047e-16
C128 824 947 2.86016e-14
C127 825 947 3.29763e-15
C126 826 947 8.3284e-14
C125 827 947 3.29763e-15
C124 828 947 8.3284e-14
C122 830 947 1.14176e-15
C120 831 947 3.29763e-15
C119 832 947 8.3284e-14
C118 833 947 8.3284e-14
C117 834 947 4.16108e-14
C116 835 947 3.01232e-14
C115 836 947 4.17738e-16
C114 837 947 3.29763e-15
C113 838 947 8.3284e-14
C112 839 947 2.96515e-13
C111 840 947 8.3284e-14
C110 841 947 3.00265e-14
C109 842 947 3.09307e-14
C106 845 947 3.4793e-14
C105 846 947 2.81118e-14
C104 847 947 3.29763e-15
C103 848 947 8.3284e-14
C102 849 947 3.95849e-14
C101 850 947 8.3284e-14
C100 851 947 3.29763e-15
C99 852 947 8.3284e-14
C98 853 947 3.29763e-15
C97 854 947 2.96515e-13
C96 855 947 8.3284e-14
C89 861 947 6.26155e-14
C88 862 947 1.09103e-14
C86 864 947 1.44675e-14
C85 865 947 2.45462e-14
C84 866 947 2.42101e-14
C83 867 947 2.75058e-14
C82 868 947 2.09836e-14
C80 870 947 8.63047e-16
C78 871 947 2.76492e-14
C77 872 947 2.83173e-14
C76 873 947 3.01232e-14
C75 874 947 4.17738e-16
C74 875 947 2.7614e-14
C73 876 947 2.86016e-14
C70 879 947 2.44873e-14
C69 880 947 4.93034e-14
C68 881 947 2.16616e-14
C66 883 947 4.17738e-16
C60 888 947 2.73747e-14
C59 889 947 2.23168e-14
C58 890 947 3.01232e-14
C56 892 947 5.73118e-14
C55 893 947 3.09307e-14
C54 894 947 2.81118e-14
C53 895 947 1.14176e-15
C52 896 947 3.4793e-14
C51 897 947 2.01557e-14
C50 898 947 5.4229e-14
C49 899 947 3.16939e-13
C48 900 947 1.44675e-14
C47 901 947 5.27918e-15
C43 905 947 5.27918e-15
C39 909 947 1.87176e-11
C38 910 947 1.07568e-13
C37 911 947 3.38702e-14
C35 913 947 2.08974e-14
C34 914 947 1.89138e-14
C32 916 947 1.5113e-14
C31 917 947 2.46362e-15
C30 918 947 9.91138e-15
C29 919 947 1.54958e-14
C27 921 947 4.90349e-14
C26 922 947 6.90483e-14
C25 923 947 9.52956e-14
C24 924 947 2.29153e-14
C23 925 947 1.61541e-13
C21 927 947 2.16616e-14
C20 928 947 1.42401e-13
C19 929 947 3.38702e-14
C17 931 947 2.08974e-14
C15 933 947 1.50518e-14
C14 934 947 2.46362e-15
C13 935 947 9.91138e-15
C12 936 947 1.89138e-14
C10 938 947 4.42848e-14
C9 939 947 6.90483e-14
C8 940 947 1.54958e-14
C7 941 947 9.52956e-14
C6 942 947 3.35086e-14
C5 943 947 1.44415e-13
C3 945 947 1.20544e-13
C2 946 947 1.51947e-13
C1 947 947 1.69239e-11
.ends mac_cts_r_ext_ihp

