../cpu.vhdl