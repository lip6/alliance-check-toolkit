* Spice description of na3_x1
* Spice driver version 235355931
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:50

* INTERF i0 i1 i2 nq vdd vss 


.subckt na3_x1 4 5 2 3 1 8 
* NET 1 = vdd
* NET 2 = i2
* NET 3 = nq
* NET 4 = i0
* NET 5 = i1
* NET 8 = vss
Mtr_00006 1 5 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00005 3 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00004 3 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00003 3 2 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 6 4 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 7 5 6 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C8 1 8 1.93752e-15
C7 2 8 1.54941e-15
C6 3 8 2.85687e-15
C5 4 8 2.12096e-15
C4 5 8 1.81693e-15
C1 8 8 1.41822e-15
.ends na3_x1

