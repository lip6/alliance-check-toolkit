-- no model for diode_w1
