* Spice description of noa2ao222_x1
* Spice driver version 1804295963
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:13

* INTERF i0 i1 i2 i3 i4 nq vdd vss 


.subckt noa2ao222_x1 10 7 5 4 6 8 3 12 
* NET 3 = vdd
* NET 4 = i3
* NET 5 = i2
* NET 6 = i4
* NET 7 = i1
* NET 8 = nq
* NET 10 = i0
* NET 12 = vss
Mtr_00010 2 4 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 1 5 8 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 8 6 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 2 7 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 3 10 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 9 4 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.21U AS=0.5304P AD=0.5304P PS=4.9U PD=4.9U 
Mtr_00004 12 5 9 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.21U AS=0.5304P AD=0.5304P PS=4.9U PD=4.9U 
Mtr_00003 9 6 8 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.21U AS=0.5304P AD=0.5304P PS=4.9U PD=4.9U 
Mtr_00002 8 7 11 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.21U AS=0.5304P AD=0.5304P PS=4.9U PD=4.9U 
Mtr_00001 11 10 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.21U AS=0.5304P AD=0.5304P PS=4.9U PD=4.9U 
C11 2 12 1.03614e-15
C10 3 12 1.95945e-15
C9 4 12 1.65532e-15
C8 5 12 1.67465e-15
C7 6 12 1.37008e-15
C6 7 12 1.67411e-15
C5 8 12 1.86634e-15
C4 9 12 4.67807e-16
C3 10 12 1.61613e-15
C1 12 12 2.26122e-15
.ends noa2ao222_x1

