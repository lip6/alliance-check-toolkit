*
* 

*****************

.TEMP 25

******************
* BSIM4 transistor model parameters for ngspice
*.lib /users/soft/analogdesign/scalable/techno/sky130_models_20220217/C4M.Sky130_all_lib.spice logic_tt 

*******************************
*Simulation conditions

Vground evss 0 0
Vsupply evdd 0 DC 1.8
*gfoncd evdd 0 evdd 0 1.0e-15

******************
* circuit model
* include circuit netlist
.include picorv32_cts_r.spi
*****************

*****************
* Circuit Instantiation
*.subckt inv_x2 vdd vss i nq


Xc 29046 59800 59787 59785 59775 59782 59774 59786 59762 59751 59760 59745 59761 59734 59724 59732 59713 59709 59712 59699 59694 59697 59698 59684 59672 59666 59663 59655 59652 59648 59639 59637 59636 59635 59623 59618 59613 59607 59599 59592 59589 59579 59574 59567 59562 59555 59546 59541 59534 59528 59523 59514 59508 59503 59495 59487 59482 59481 59471 59465 59460 59453 59452 59451 59449 10344 91 90 48122 46977 56766 56782 57428 53693 56151 55030 56133 55027 55024 53671 55021 53036 51222 53032 49277 53690 46981 48118 49257 45603 49904 49274 51778 50609 45618 46234 46229 48112 9238 51219 49888 51206 51761 50587 51203 49871 49866 55555 54372 55017 50576 51200 55004 56113 56119 58162 56778 55542 57423 58771 58775 51183 51740 52361 53685 53024 53652 52368 58764 58768 51746 15005 44234 14291 14458 13919 59251 59242 59238 59228 58597 58605 57778 57233 57096 56042 55376 54776 54283 53964 53342 52686 52050 51433 51123 50509 50166 49567 48511 47936 48577 49147 49146 48576 46894 47470 46128 44895 6527 9103 59441 59436 59428 59424 59415 59410 59409 59403 59398 59388 59384 59375 59373 59392 59360 59353 59438 59339 59335 59334 59425 59322 59315 59307 59300 59296 59288 59282 59275 59411 59262 59254 16114 15465 14671 14215 28223 27583 26416 25242 24081 23579 22934 22368 21751 21609 21177 20345 19912 19088 18586 17936 17491 16868 16277 16278 15623 15031 15622 14380 14379 13214 12637 12638 10766 10611 10221 9552 31325 8541 44871 41853 43768 42446 44861 46884 59031 59030 58413 57251 56542 55978 55377 54843 54658 54028 53495 53492 52220 52045 51428 50445 50162 49540 48900 48368 48365 47215 46681 46068 28657 28060 27449 26867 33763 32083 31441 27153 32692 29634 33253 31429 30186 26630 21280 21284 20707 19245 18621 18585 22076 17332 17592 18782 5997 28434 324 692 323 691 322 321 320 310 676 309 303 671 665 293 291 281 279 1039 270 268 259 258 257 256 246 245 244 234 232 231 230 229 218 216 215 564 7546 14438 evdd evss picorv32_cts_r 
.end

