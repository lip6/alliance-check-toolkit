* Spice description of oa2ao222_x2
* Spice driver version -462962917
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:33

* INTERF i0 i1 i2 i3 i4 q vdd vss 


.subckt oa2ao222_x2 11 8 6 4 7 5 3 13 
* NET 3 = vdd
* NET 4 = i3
* NET 5 = q
* NET 6 = i2
* NET 7 = i4
* NET 8 = i1
* NET 11 = i0
* NET 13 = vss
Mtr_00012 5 9 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 3 11 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 2 8 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 9 7 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 1 6 9 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 2 4 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 10 4 13 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00005 13 6 10 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00004 5 9 13 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00003 12 11 13 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00002 10 7 9 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00001 9 8 12 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
C12 2 13 1.02094e-15
C11 3 13 2.65269e-15
C10 4 13 1.49761e-15
C9 5 13 2.20321e-15
C8 6 13 1.35774e-15
C7 7 13 1.33872e-15
C6 8 13 1.64275e-15
C5 9 13 2.07157e-15
C4 10 13 5.43814e-16
C3 11 13 1.9559e-15
C1 13 13 2.85619e-15
.ends oa2ao222_x2

