* GuardRing_P418W1550HFF
* GuardRing_P418W1550HFF
.subckt GuardRing_P418W1550HFF conn

.ends GuardRing_P418W1550HFF
