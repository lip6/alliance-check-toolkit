* Spice description of sff1_x4
* Spice driver version 1835101979
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:40

* INTERF ck i q vdd vss 


.subckt sff1_x4 15 12 5 4 17 
* NET 4 = vdd
* NET 5 = q
* NET 7 = sff_s
* NET 8 = y
* NET 9 = sff_m
* NET 12 = i
* NET 13 = ckr
* NET 14 = u
* NET 15 = ck
* NET 16 = nckr
* NET 17 = vss
Mtr_00026 5 7 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00025 4 7 5 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00024 7 16 8 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00023 8 9 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00022 4 8 3 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00021 3 16 9 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00020 9 13 2 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00019 4 12 14 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00018 4 15 16 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00017 13 16 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.38U AS=0.5712P AD=0.5712P PS=5.24U PD=5.24U 
Mtr_00016 4 5 1 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00015 1 13 7 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00014 2 14 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00013 17 7 5 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00012 5 7 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00011 7 13 8 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00010 17 8 11 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00009 8 9 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00008 9 16 10 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00007 17 12 14 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00006 13 16 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00005 17 15 16 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00004 17 5 6 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00003 6 16 7 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 11 13 9 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 10 14 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
C14 4 17 5.8351e-15
C13 5 17 3.29526e-15
C11 7 17 2.21812e-15
C10 8 17 1.99446e-15
C9 9 17 2.3045e-15
C6 12 17 2.91895e-15
C5 13 17 3.90607e-15
C4 14 17 2.21801e-15
C3 15 17 1.94911e-15
C2 16 17 3.95204e-15
C1 17 17 5.66544e-15
.ends sff1_x4

