-- no model for or21nand_x0
