picorv32_m_hitas
*
* sta compatible ngspice
* taking into account modified library

*****************

.TEMP 25

******************
******************
*Technology is loaded in the db_ng.tcl file
*******************************

*******************************
*Simulation conditions

Vground evss 0 0
Vsupply evdd 0 DC 1.8
*gfoncd evdd 0 evdd 0 1.0e-15

******************
* circuit model
* include circuit netlist
.INCLUDE /users/cao/mariem/coriolis-2.x/src/alliance-check-toolkit/benchs/picorv32/skyWater130/timing/sta/picorv32_m.spi
*****************

*****************
* Circuit Instantiation
*.subckt picorv32_m VGND VPWR clk eoi[0] eoi[15] eoi[1] eoi[2] eoi[3] eoi[4] eoi[5] irq[0]
*+ irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[16] irq[17] irq[18] irq[19]
*+ irq[1] irq[20] irq[21] irq[22] irq[23] irq[24] irq[25] irq[26] irq[27] irq[28] irq[29]
*+ irq[2] irq[30] irq[31] irq[3] irq[4] irq[5] irq[6] irq[7] irq[8] irq[9] mem_addr[10]
*+ mem_addr[11] mem_addr[12] mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[16] mem_addr[17]
*+ mem_addr[18] mem_addr[19] mem_addr[20] mem_addr[21] mem_addr[22] mem_addr[23] mem_addr[24]
*+ mem_addr[25] mem_addr[26] mem_addr[27] mem_addr[28] mem_addr[29] mem_addr[2] mem_addr[30]
*+ mem_addr[31] mem_addr[3] mem_addr[4] mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8]
*+ mem_addr[9] mem_instr mem_la_addr[0] mem_la_addr[10] mem_la_addr[11] mem_la_addr[12]
*+ mem_la_addr[13] mem_la_addr[14] mem_la_addr[15] mem_la_addr[16] mem_la_addr[17]
*+ mem_la_addr[18] mem_la_addr[19] mem_la_addr[1] mem_la_addr[20] mem_la_addr[21] mem_la_addr[22]
*+ mem_la_addr[23] mem_la_addr[24] mem_la_addr[25] mem_la_addr[26] mem_la_addr[27]
*+ mem_la_addr[28] mem_la_addr[29] mem_la_addr[2] mem_la_addr[30] mem_la_addr[31] mem_la_addr[3]
*+ mem_la_addr[4] mem_la_addr[5] mem_la_addr[6] mem_la_addr[7] mem_la_addr[8] mem_la_addr[9]
*+ mem_la_read mem_la_wdata[0] mem_la_wdata[10] mem_la_wdata[11] mem_la_wdata[12] mem_la_wdata[13]
*+ mem_la_wdata[14] mem_la_wdata[15] mem_la_wdata[16] mem_la_wdata[17] mem_la_wdata[18]
*+ mem_la_wdata[19] mem_la_wdata[1] mem_la_wdata[20] mem_la_wdata[21] mem_la_wdata[22]
*+ mem_la_wdata[23] mem_la_wdata[24] mem_la_wdata[25] mem_la_wdata[26] mem_la_wdata[27]
*+ mem_la_wdata[28] mem_la_wdata[29] mem_la_wdata[2] mem_la_wdata[30] mem_la_wdata[31]
*+ mem_la_wdata[3] mem_la_wdata[4] mem_la_wdata[5] mem_la_wdata[6] mem_la_wdata[7]
*+ mem_la_wdata[8] mem_la_wdata[9] mem_la_write mem_la_wstrb[0] mem_la_wstrb[1] mem_la_wstrb[2]
*+ mem_la_wstrb[3] mem_rdata[0] mem_rdata[10] mem_rdata[11] mem_rdata[12] mem_rdata[13]
*+ mem_rdata[14] mem_rdata[15] mem_rdata[16] mem_rdata[17] mem_rdata[18] mem_rdata[19]
*+ mem_rdata[1] mem_rdata[20] mem_rdata[21] mem_rdata[22] mem_rdata[23] mem_rdata[24]
*+ mem_rdata[25] mem_rdata[26] mem_rdata[27] mem_rdata[28] mem_rdata[29] mem_rdata[2]
*+ mem_rdata[30] mem_rdata[31] mem_rdata[3] mem_rdata[4] mem_rdata[5] mem_rdata[6]
*+ mem_rdata[7] mem_rdata[8] mem_rdata[9] mem_ready mem_valid mem_wdata[0] mem_wdata[10]
*+ mem_wdata[11] mem_wdata[12] mem_wdata[13] mem_wdata[14] mem_wdata[15] mem_wdata[16]
*+ mem_wdata[17] mem_wdata[18] mem_wdata[19] mem_wdata[1] mem_wdata[20] mem_wdata[21]
*+ mem_wdata[22] mem_wdata[23] mem_wdata[24] mem_wdata[25] mem_wdata[26] mem_wdata[27]
*+ mem_wdata[28] mem_wdata[29] mem_wdata[2] mem_wdata[30] mem_wdata[31] mem_wdata[3]
*+ mem_wdata[4] mem_wdata[5] mem_wdata[6] mem_wdata[7] mem_wdata[8] mem_wdata[9] mem_wstrb[0]
*+ mem_wstrb[1] mem_wstrb[2] mem_wstrb[3] pcpi_insn[0] pcpi_insn[10] pcpi_insn[11]
*+ pcpi_insn[12] pcpi_insn[13] pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17]
*+ pcpi_insn[18] pcpi_insn[19] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[28]
*+ pcpi_insn[29] pcpi_insn[30] pcpi_insn[31] pcpi_insn[9] pcpi_rd[0] pcpi_rd[10] pcpi_rd[11]
*+ pcpi_rd[12] pcpi_rd[13] pcpi_rd[14] pcpi_rd[15] pcpi_rd[16] pcpi_rd[17] pcpi_rd[18]
*+ pcpi_rd[19] pcpi_rd[1] pcpi_rd[20] pcpi_rd[21] pcpi_rd[22] pcpi_rd[23] pcpi_rd[24]
*+ pcpi_rd[25] pcpi_rd[26] pcpi_rd[27] pcpi_rd[28] pcpi_rd[29] pcpi_rd[2] pcpi_rd[30]
*+ pcpi_rd[31] pcpi_rd[3] pcpi_rd[4] pcpi_rd[5] pcpi_rd[6] pcpi_rd[7] pcpi_rd[8] pcpi_rd[9]
*+ pcpi_ready pcpi_rs1[0] pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14]
*+ pcpi_rs1[15] pcpi_rs1[16] pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20]
*+ pcpi_rs1[21] pcpi_rs1[22] pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27]
*+ pcpi_rs1[28] pcpi_rs1[29] pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4]
*+ pcpi_rs1[5] pcpi_rs1[6] pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10]
*+ pcpi_rs2[11] pcpi_rs2[12] pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17]
*+ pcpi_rs2[18] pcpi_rs2[19] pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23]
*+ pcpi_rs2[24] pcpi_rs2[25] pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2]
*+ pcpi_rs2[30] pcpi_rs2[31] pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7]
*+ pcpi_rs2[8] pcpi_rs2[9] pcpi_wait pcpi_wr resetn trace_data[0] trace_data[15] trace_data[16]
*+ trace_data[1] trace_data[20] trace_data[21] trace_data[22] trace_data[23] trace_data[24]
*+ trace_data[25] trace_data[26] trace_data[27] trace_data[28] trace_data[29] trace_data[2]
*+ trace_data[35] trace_data[3] trace_data[4] trace_data[5] trace_data[6] trace_data[7]
*+ trace_data[8] trace_data[9] trace_valid trap pcpi_insn[27] pcpi_insn[26] trace_data[14]
*+ pcpi_insn[25] trace_data[13] pcpi_insn[24] trace_data[12] trace_data[34] pcpi_insn[23]
*+ trace_data[33] trace_data[11] trace_data[32] trace_data[10] pcpi_valid trace_data[31]
*+ trace_data[30] trace_data[19] trace_data[18] trace_data[17] eoi[14] eoi[25] eoi[24]
*+ eoi[13] eoi[23] eoi[12] mem_addr[1] pcpi_insn[8] eoi[11] eoi[22] pcpi_insn[7] mem_addr[0]
*+ eoi[21] eoi[10] pcpi_insn[6] eoi[31] eoi[9] eoi[20] pcpi_insn[5] eoi[30] eoi[19]
*+ eoi[8] eoi[18] eoi[29] pcpi_insn[4] eoi[7] eoi[28] eoi[17] pcpi_insn[3] eoi[6] eoi[27]
*+ pcpi_insn[2] eoi[16] pcpi_insn[1] eoi[26]




Xpicorv32_m evss evdd clk eoi[0] eoi[15] eoi[1] eoi[2] eoi[3] eoi[4] eoi[5] irq[0]
+ irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[16] irq[17] irq[18] irq[19]
+ irq[1] irq[20] irq[21] irq[22] irq[23] irq[24] irq[25] irq[26] irq[27] irq[28] irq[29]
+ irq[2] irq[30] irq[31] irq[3] irq[4] irq[5] irq[6] irq[7] irq[8] irq[9] mem_addr[10]
+ mem_addr[11] mem_addr[12] mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[16] mem_addr[17]
+ mem_addr[18] mem_addr[19] mem_addr[20] mem_addr[21] mem_addr[22] mem_addr[23] mem_addr[24]
+ mem_addr[25] mem_addr[26] mem_addr[27] mem_addr[28] mem_addr[29] mem_addr[2] mem_addr[30]
+ mem_addr[31] mem_addr[3] mem_addr[4] mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8]
+ mem_addr[9] mem_instr mem_la_addr[0] mem_la_addr[10] mem_la_addr[11] mem_la_addr[12]
+ mem_la_addr[13] mem_la_addr[14] mem_la_addr[15] mem_la_addr[16] mem_la_addr[17]
+ mem_la_addr[18] mem_la_addr[19] mem_la_addr[1] mem_la_addr[20] mem_la_addr[21] mem_la_addr[22]
+ mem_la_addr[23] mem_la_addr[24] mem_la_addr[25] mem_la_addr[26] mem_la_addr[27]
+ mem_la_addr[28] mem_la_addr[29] mem_la_addr[2] mem_la_addr[30] mem_la_addr[31] mem_la_addr[3]
+ mem_la_addr[4] mem_la_addr[5] mem_la_addr[6] mem_la_addr[7] mem_la_addr[8] mem_la_addr[9]
+ mem_la_read mem_la_wdata[0] mem_la_wdata[10] mem_la_wdata[11] mem_la_wdata[12] mem_la_wdata[13]
+ mem_la_wdata[14] mem_la_wdata[15] mem_la_wdata[16] mem_la_wdata[17] mem_la_wdata[18]
+ mem_la_wdata[19] mem_la_wdata[1] mem_la_wdata[20] mem_la_wdata[21] mem_la_wdata[22]
+ mem_la_wdata[23] mem_la_wdata[24] mem_la_wdata[25] mem_la_wdata[26] mem_la_wdata[27]
+ mem_la_wdata[28] mem_la_wdata[29] mem_la_wdata[2] mem_la_wdata[30] mem_la_wdata[31]
+ mem_la_wdata[3] mem_la_wdata[4] mem_la_wdata[5] mem_la_wdata[6] mem_la_wdata[7]
+ mem_la_wdata[8] mem_la_wdata[9] mem_la_write mem_la_wstrb[0] mem_la_wstrb[1] mem_la_wstrb[2]
+ mem_la_wstrb[3] mem_rdata[0] mem_rdata[10] mem_rdata[11] mem_rdata[12] mem_rdata[13]
+ mem_rdata[14] mem_rdata[15] mem_rdata[16] mem_rdata[17] mem_rdata[18] mem_rdata[19]
+ mem_rdata[1] mem_rdata[20] mem_rdata[21] mem_rdata[22] mem_rdata[23] mem_rdata[24]
+ mem_rdata[25] mem_rdata[26] mem_rdata[27] mem_rdata[28] mem_rdata[29] mem_rdata[2]
+ mem_rdata[30] mem_rdata[31] mem_rdata[3] mem_rdata[4] mem_rdata[5] mem_rdata[6]
+ mem_rdata[7] mem_rdata[8] mem_rdata[9] mem_ready mem_valid mem_wdata[0] mem_wdata[10]
+ mem_wdata[11] mem_wdata[12] mem_wdata[13] mem_wdata[14] mem_wdata[15] mem_wdata[16]
+ mem_wdata[17] mem_wdata[18] mem_wdata[19] mem_wdata[1] mem_wdata[20] mem_wdata[21]
+ mem_wdata[22] mem_wdata[23] mem_wdata[24] mem_wdata[25] mem_wdata[26] mem_wdata[27]
+ mem_wdata[28] mem_wdata[29] mem_wdata[2] mem_wdata[30] mem_wdata[31] mem_wdata[3]
+ mem_wdata[4] mem_wdata[5] mem_wdata[6] mem_wdata[7] mem_wdata[8] mem_wdata[9] mem_wstrb[0]
+ mem_wstrb[1] mem_wstrb[2] mem_wstrb[3] pcpi_insn[0] pcpi_insn[10] pcpi_insn[11]
+ pcpi_insn[12] pcpi_insn[13] pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17]
+ pcpi_insn[18] pcpi_insn[19] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[28]
+ pcpi_insn[29] pcpi_insn[30] pcpi_insn[31] pcpi_insn[9] pcpi_rd[0] pcpi_rd[10] pcpi_rd[11]
+ pcpi_rd[12] pcpi_rd[13] pcpi_rd[14] pcpi_rd[15] pcpi_rd[16] pcpi_rd[17] pcpi_rd[18]
+ pcpi_rd[19] pcpi_rd[1] pcpi_rd[20] pcpi_rd[21] pcpi_rd[22] pcpi_rd[23] pcpi_rd[24]
+ pcpi_rd[25] pcpi_rd[26] pcpi_rd[27] pcpi_rd[28] pcpi_rd[29] pcpi_rd[2] pcpi_rd[30]
+ pcpi_rd[31] pcpi_rd[3] pcpi_rd[4] pcpi_rd[5] pcpi_rd[6] pcpi_rd[7] pcpi_rd[8] pcpi_rd[9]
+ pcpi_ready pcpi_rs1[0] pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14]
+ pcpi_rs1[15] pcpi_rs1[16] pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20]
+ pcpi_rs1[21] pcpi_rs1[22] pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27]
+ pcpi_rs1[28] pcpi_rs1[29] pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4]
+ pcpi_rs1[5] pcpi_rs1[6] pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10]
+ pcpi_rs2[11] pcpi_rs2[12] pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17]
+ pcpi_rs2[18] pcpi_rs2[19] pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23]
+ pcpi_rs2[24] pcpi_rs2[25] pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2]
+ pcpi_rs2[30] pcpi_rs2[31] pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7]
+ pcpi_rs2[8] pcpi_rs2[9] pcpi_wait pcpi_wr resetn trace_data[0] trace_data[15] trace_data[16]
+ trace_data[1] trace_data[20] trace_data[21] trace_data[22] trace_data[23] trace_data[24]
+ trace_data[25] trace_data[26] trace_data[27] trace_data[28] trace_data[29] trace_data[2]
+ trace_data[35] trace_data[3] trace_data[4] trace_data[5] trace_data[6] trace_data[7]
+ trace_data[8] trace_data[9] trace_valid trap pcpi_insn[27] pcpi_insn[26] trace_data[14]
+ pcpi_insn[25] trace_data[13] pcpi_insn[24] trace_data[12] trace_data[34] pcpi_insn[23]
+ trace_data[33] trace_data[11] trace_data[32] trace_data[10] pcpi_valid trace_data[31]
+ trace_data[30] trace_data[19] trace_data[18] trace_data[17] eoi[14] eoi[25] eoi[24]
+ eoi[13] eoi[23] eoi[12] mem_addr[1] pcpi_insn[8] eoi[11] eoi[22] pcpi_insn[7] mem_addr[0]
+ eoi[21] eoi[10] pcpi_insn[6] eoi[31] eoi[9] eoi[20] pcpi_insn[5] eoi[30] eoi[19]
+ eoi[8] eoi[18] eoi[29] pcpi_insn[4] eoi[7] eoi[28] eoi[17] pcpi_insn[3] eoi[6] eoi[27]
+ pcpi_insn[2] eoi[16] pcpi_insn[1] eoi[26] picorv32_m

.end

