* Gallery
.subckt Gallery vss vdd
Xfill[0] vdd vss fill
Xdffnr_x1[1] vdd vss dffnr_x1[1].[_InstanceNet[i], 'Gallery'] dffnr_x1[1].[_InstanceNet[clk], 'Gallery'] dffnr_x1[1].[_InstanceNet[q], 'Gallery'] dffnr_x1[1].[_InstanceNet[nrst], 'Gallery'] dffnr_x1
Xdffnr_x1[2] vdd vss dffnr_x1[2].[_InstanceNet[i], 'Gallery'] dffnr_x1[2].[_InstanceNet[clk], 'Gallery'] dffnr_x1[2].[_InstanceNet[q], 'Gallery'] dffnr_x1[2].[_InstanceNet[nrst], 'Gallery'] dffnr_x1
Xtie[0] vdd vss tie
Xdff_x1[1] vdd vss dff_x1[1].[_InstanceNet[i], 'Gallery'] dff_x1[1].[_InstanceNet[clk], 'Gallery'] dff_x1[1].[_InstanceNet[q], 'Gallery'] dff_x1
Xfill[2] vdd vss fill
Xtie_diff[0] vdd vss tie_diff
Xnsnrlatch_x1[1] vdd vss nsnrlatch_x1[1].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x1[1].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x1[1].[_InstanceNet[q], 'Gallery'] nsnrlatch_x1[1].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x1
Xdff_x1[2] vdd vss dff_x1[2].[_InstanceNet[i], 'Gallery'] dff_x1[2].[_InstanceNet[clk], 'Gallery'] dff_x1[2].[_InstanceNet[q], 'Gallery'] dff_x1
Xtie_poly[0] vdd vss tie_poly
Xnsnrlatch_x0[1] vdd vss nsnrlatch_x0[1].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x0[1].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x0[1].[_InstanceNet[q], 'Gallery'] nsnrlatch_x0[1].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x0
Xtie[2] vdd vss tie
Xfill_w2[0] vdd vss fill_w2
Xnexor2_x0[1] vdd vss nexor2_x0[1].[_InstanceNet[i0], 'Gallery'] nexor2_x0[1].[_InstanceNet[i1], 'Gallery'] nexor2_x0[1].[_InstanceNet[nq], 'Gallery'] nexor2_x0
Xnsnrlatch_x1[2] vdd vss nsnrlatch_x1[2].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x1[2].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x1[2].[_InstanceNet[q], 'Gallery'] nsnrlatch_x1[2].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x1
Xtie_w2[0] vdd vss tie_w2
Xxor2_x0[1] vdd vss xor2_x0[1].[_InstanceNet[i0], 'Gallery'] xor2_x0[1].[_InstanceNet[i1], 'Gallery'] xor2_x0[1].[_InstanceNet[q], 'Gallery'] xor2_x0
Xtie_diff[2] vdd vss tie_diff
Xtie_diff_w2[0] vdd vss tie_diff_w2
Xor21nand_x1[1] vdd vss or21nand_x1[1].[_InstanceNet[nq], 'Gallery'] or21nand_x1[1].[_InstanceNet[i0], 'Gallery'] or21nand_x1[1].[_InstanceNet[i1], 'Gallery'] or21nand_x1[1].[_InstanceNet[i2], 'Gallery'] or21nand_x1
Xnsnrlatch_x0[2] vdd vss nsnrlatch_x0[2].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x0[2].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x0[2].[_InstanceNet[q], 'Gallery'] nsnrlatch_x0[2].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x0
Xtie_poly_w2[0] vdd vss tie_poly_w2
Xor21nand_x0[1] vdd vss or21nand_x0[1].[_InstanceNet[nq], 'Gallery'] or21nand_x0[1].[_InstanceNet[i0], 'Gallery'] or21nand_x0[1].[_InstanceNet[i1], 'Gallery'] or21nand_x0[1].[_InstanceNet[i2], 'Gallery'] or21nand_x0
Xtie_poly[2] vdd vss tie_poly
Xfill_w4[0] vdd vss fill_w4
Xand21nor_x1[1] vdd vss and21nor_x1[1].[_InstanceNet[nq], 'Gallery'] and21nor_x1[1].[_InstanceNet[i0], 'Gallery'] and21nor_x1[1].[_InstanceNet[i1], 'Gallery'] and21nor_x1[1].[_InstanceNet[i2], 'Gallery'] and21nor_x1
Xnexor2_x0[2] vdd vss nexor2_x0[2].[_InstanceNet[i0], 'Gallery'] nexor2_x0[2].[_InstanceNet[i1], 'Gallery'] nexor2_x0[2].[_InstanceNet[nq], 'Gallery'] nexor2_x0
Xtie_w4[0] vdd vss tie_w4
Xand21nor_x0[1] vdd vss and21nor_x0[1].[_InstanceNet[nq], 'Gallery'] and21nor_x0[1].[_InstanceNet[i0], 'Gallery'] and21nor_x0[1].[_InstanceNet[i1], 'Gallery'] and21nor_x0[1].[_InstanceNet[i2], 'Gallery'] and21nor_x0
Xfill_w2[2] vdd vss fill_w2
Xtie_diff_w4[0] vdd vss tie_diff_w4
Xmux2_x1[1] vdd vss mux2_x1[1].[_InstanceNet[i0], 'Gallery'] mux2_x1[1].[_InstanceNet[i1], 'Gallery'] mux2_x1[1].[_InstanceNet[cmd], 'Gallery'] mux2_x1[1].[_InstanceNet[q], 'Gallery'] mux2_x1
Xxor2_x0[2] vdd vss xor2_x0[2].[_InstanceNet[i0], 'Gallery'] xor2_x0[2].[_InstanceNet[i1], 'Gallery'] xor2_x0[2].[_InstanceNet[q], 'Gallery'] xor2_x0
Xtie_poly_w4[0] vdd vss tie_poly_w4
Xor4_x1[1] vdd vss or4_x1[1].[_InstanceNet[q], 'Gallery'] or4_x1[1].[_InstanceNet[i0], 'Gallery'] or4_x1[1].[_InstanceNet[i1], 'Gallery'] or4_x1[1].[_InstanceNet[i2], 'Gallery'] or4_x1[1].[_InstanceNet[i3], 'Gallery'] or4_x1
Xtie_w2[2] vdd vss tie_w2
Xdiode_w1[0] vdd vss diode_w1[0].[_InstanceNet[i], 'Gallery'] diode_w1
Xor3_x1[1] vdd vss or3_x1[1].[_InstanceNet[q], 'Gallery'] or3_x1[1].[_InstanceNet[i0], 'Gallery'] or3_x1[1].[_InstanceNet[i1], 'Gallery'] or3_x1[1].[_InstanceNet[i2], 'Gallery'] or3_x1
Xor21nand_x1[2] vdd vss or21nand_x1[2].[_InstanceNet[nq], 'Gallery'] or21nand_x1[2].[_InstanceNet[i0], 'Gallery'] or21nand_x1[2].[_InstanceNet[i1], 'Gallery'] or21nand_x1[2].[_InstanceNet[i2], 'Gallery'] or21nand_x1
Xzero_x1[0] vdd vss zero_x1[0].[_InstanceNet[zero], 'Gallery'] zero_x1
Xor2_x1[1] vdd vss or2_x1[1].[_InstanceNet[q], 'Gallery'] or2_x1[1].[_InstanceNet[i0], 'Gallery'] or2_x1[1].[_InstanceNet[i1], 'Gallery'] or2_x1
Xtie_diff_w2[2] vdd vss tie_diff_w2
Xone_x1[0] vdd vss one_x1[0].[_InstanceNet[one], 'Gallery'] one_x1
Xnor4_x1[1] vdd vss nor4_x1[1].[_InstanceNet[nq], 'Gallery'] nor4_x1[1].[_InstanceNet[i0], 'Gallery'] nor4_x1[1].[_InstanceNet[i1], 'Gallery'] nor4_x1[1].[_InstanceNet[i2], 'Gallery'] nor4_x1[1].[_InstanceNet[i3], 'Gallery'] nor4_x1
Xor21nand_x0[2] vdd vss or21nand_x0[2].[_InstanceNet[nq], 'Gallery'] or21nand_x0[2].[_InstanceNet[i0], 'Gallery'] or21nand_x0[2].[_InstanceNet[i1], 'Gallery'] or21nand_x0[2].[_InstanceNet[i2], 'Gallery'] or21nand_x0
Xzeroone_x1[0] vdd vss zeroone_x1[0].[_InstanceNet[one], 'Gallery'] zeroone_x1[0].[_InstanceNet[zero], 'Gallery'] zeroone_x1
Xnor4_x0[1] vdd vss nor4_x0[1].[_InstanceNet[nq], 'Gallery'] nor4_x0[1].[_InstanceNet[i0], 'Gallery'] nor4_x0[1].[_InstanceNet[i1], 'Gallery'] nor4_x0[1].[_InstanceNet[i2], 'Gallery'] nor4_x0[1].[_InstanceNet[i3], 'Gallery'] nor4_x0
Xtie_poly_w2[2] vdd vss tie_poly_w2
Xdecap_w0[0] vdd vss decap_w0
Xnor3_x1[1] vdd vss nor3_x1[1].[_InstanceNet[nq], 'Gallery'] nor3_x1[1].[_InstanceNet[i0], 'Gallery'] nor3_x1[1].[_InstanceNet[i1], 'Gallery'] nor3_x1[1].[_InstanceNet[i2], 'Gallery'] nor3_x1
Xand21nor_x1[2] vdd vss and21nor_x1[2].[_InstanceNet[nq], 'Gallery'] and21nor_x1[2].[_InstanceNet[i0], 'Gallery'] and21nor_x1[2].[_InstanceNet[i1], 'Gallery'] and21nor_x1[2].[_InstanceNet[i2], 'Gallery'] and21nor_x1
Xinv_x0[0] vdd vss inv_x0[0].[_InstanceNet[i], 'Gallery'] inv_x0[0].[_InstanceNet[nq], 'Gallery'] inv_x0
Xnor3_x0[1] vdd vss nor3_x0[1].[_InstanceNet[nq], 'Gallery'] nor3_x0[1].[_InstanceNet[i0], 'Gallery'] nor3_x0[1].[_InstanceNet[i1], 'Gallery'] nor3_x0[1].[_InstanceNet[i2], 'Gallery'] nor3_x0
Xfill_w4[2] vdd vss fill_w4
Xinv_x1[0] vdd vss inv_x1[0].[_InstanceNet[i], 'Gallery'] inv_x1[0].[_InstanceNet[nq], 'Gallery'] inv_x1
Xnor2_x1[1] vdd vss nor2_x1[1].[_InstanceNet[nq], 'Gallery'] nor2_x1[1].[_InstanceNet[i0], 'Gallery'] nor2_x1[1].[_InstanceNet[i1], 'Gallery'] nor2_x1
Xand21nor_x0[2] vdd vss and21nor_x0[2].[_InstanceNet[nq], 'Gallery'] and21nor_x0[2].[_InstanceNet[i0], 'Gallery'] and21nor_x0[2].[_InstanceNet[i1], 'Gallery'] and21nor_x0[2].[_InstanceNet[i2], 'Gallery'] and21nor_x0
Xinv_x2[0] vdd vss inv_x2[0].[_InstanceNet[i], 'Gallery'] inv_x2[0].[_InstanceNet[nq], 'Gallery'] inv_x2
Xnor2_x0[1] vdd vss nor2_x0[1].[_InstanceNet[nq], 'Gallery'] nor2_x0[1].[_InstanceNet[i0], 'Gallery'] nor2_x0[1].[_InstanceNet[i1], 'Gallery'] nor2_x0
Xtie_w4[2] vdd vss tie_w4
Xinv_x4[0] vdd vss inv_x4[0].[_InstanceNet[i], 'Gallery'] inv_x4[0].[_InstanceNet[nq], 'Gallery'] inv_x4
Xand4_x1[1] vdd vss and4_x1[1].[_InstanceNet[q], 'Gallery'] and4_x1[1].[_InstanceNet[i0], 'Gallery'] and4_x1[1].[_InstanceNet[i1], 'Gallery'] and4_x1[1].[_InstanceNet[i2], 'Gallery'] and4_x1[1].[_InstanceNet[i3], 'Gallery'] and4_x1
Xmux2_x1[2] vdd vss mux2_x1[2].[_InstanceNet[i0], 'Gallery'] mux2_x1[2].[_InstanceNet[i1], 'Gallery'] mux2_x1[2].[_InstanceNet[cmd], 'Gallery'] mux2_x1[2].[_InstanceNet[q], 'Gallery'] mux2_x1
Xbuf_x1[0] vdd vss buf_x1[0].[_InstanceNet[i], 'Gallery'] buf_x1[0].[_InstanceNet[q], 'Gallery'] buf_x1
Xand3_x1[1] vdd vss and3_x1[1].[_InstanceNet[q], 'Gallery'] and3_x1[1].[_InstanceNet[i0], 'Gallery'] and3_x1[1].[_InstanceNet[i1], 'Gallery'] and3_x1[1].[_InstanceNet[i2], 'Gallery'] and3_x1
Xtie_diff_w4[2] vdd vss tie_diff_w4
Xbuf_x2[0] vdd vss buf_x2[0].[_InstanceNet[i], 'Gallery'] buf_x2[0].[_InstanceNet[q], 'Gallery'] buf_x2
Xand2_x1[1] vdd vss and2_x1[1].[_InstanceNet[q], 'Gallery'] and2_x1[1].[_InstanceNet[i0], 'Gallery'] and2_x1[1].[_InstanceNet[i1], 'Gallery'] and2_x1
Xor4_x1[2] vdd vss or4_x1[2].[_InstanceNet[q], 'Gallery'] or4_x1[2].[_InstanceNet[i0], 'Gallery'] or4_x1[2].[_InstanceNet[i1], 'Gallery'] or4_x1[2].[_InstanceNet[i2], 'Gallery'] or4_x1[2].[_InstanceNet[i3], 'Gallery'] or4_x1
Xbuf_x4[0] vdd vss buf_x4[0].[_InstanceNet[i], 'Gallery'] buf_x4[0].[_InstanceNet[q], 'Gallery'] buf_x4
Xnand4_x1[1] vdd vss nand4_x1[1].[_InstanceNet[nq], 'Gallery'] nand4_x1[1].[_InstanceNet[i0], 'Gallery'] nand4_x1[1].[_InstanceNet[i1], 'Gallery'] nand4_x1[1].[_InstanceNet[i2], 'Gallery'] nand4_x1[1].[_InstanceNet[i3], 'Gallery'] nand4_x1
Xtie_poly_w4[2] vdd vss tie_poly_w4
Xnand2_x0[0] vdd vss nand2_x0[0].[_InstanceNet[nq], 'Gallery'] nand2_x0[0].[_InstanceNet[i0], 'Gallery'] nand2_x0[0].[_InstanceNet[i1], 'Gallery'] nand2_x0
Xnand4_x0[1] vdd vss nand4_x0[1].[_InstanceNet[nq], 'Gallery'] nand4_x0[1].[_InstanceNet[i0], 'Gallery'] nand4_x0[1].[_InstanceNet[i1], 'Gallery'] nand4_x0[1].[_InstanceNet[i2], 'Gallery'] nand4_x0[1].[_InstanceNet[i3], 'Gallery'] nand4_x0
Xor3_x1[2] vdd vss or3_x1[2].[_InstanceNet[q], 'Gallery'] or3_x1[2].[_InstanceNet[i0], 'Gallery'] or3_x1[2].[_InstanceNet[i1], 'Gallery'] or3_x1[2].[_InstanceNet[i2], 'Gallery'] or3_x1
Xnand2_x1[0] vdd vss nand2_x1[0].[_InstanceNet[nq], 'Gallery'] nand2_x1[0].[_InstanceNet[i0], 'Gallery'] nand2_x1[0].[_InstanceNet[i1], 'Gallery'] nand2_x1
Xnand3_x1[1] vdd vss nand3_x1[1].[_InstanceNet[nq], 'Gallery'] nand3_x1[1].[_InstanceNet[i0], 'Gallery'] nand3_x1[1].[_InstanceNet[i1], 'Gallery'] nand3_x1[1].[_InstanceNet[i2], 'Gallery'] nand3_x1
Xdiode_w1[2] vdd vss diode_w1[2].[_InstanceNet[i], 'Gallery'] diode_w1
Xnand3_x0[0] vdd vss nand3_x0[0].[_InstanceNet[nq], 'Gallery'] nand3_x0[0].[_InstanceNet[i0], 'Gallery'] nand3_x0[0].[_InstanceNet[i1], 'Gallery'] nand3_x0[0].[_InstanceNet[i2], 'Gallery'] nand3_x0
Xnand3_x0[1] vdd vss nand3_x0[1].[_InstanceNet[nq], 'Gallery'] nand3_x0[1].[_InstanceNet[i0], 'Gallery'] nand3_x0[1].[_InstanceNet[i1], 'Gallery'] nand3_x0[1].[_InstanceNet[i2], 'Gallery'] nand3_x0
Xor2_x1[2] vdd vss or2_x1[2].[_InstanceNet[q], 'Gallery'] or2_x1[2].[_InstanceNet[i0], 'Gallery'] or2_x1[2].[_InstanceNet[i1], 'Gallery'] or2_x1
Xnand3_x1[0] vdd vss nand3_x1[0].[_InstanceNet[nq], 'Gallery'] nand3_x1[0].[_InstanceNet[i0], 'Gallery'] nand3_x1[0].[_InstanceNet[i1], 'Gallery'] nand3_x1[0].[_InstanceNet[i2], 'Gallery'] nand3_x1
Xnand2_x1[1] vdd vss nand2_x1[1].[_InstanceNet[nq], 'Gallery'] nand2_x1[1].[_InstanceNet[i0], 'Gallery'] nand2_x1[1].[_InstanceNet[i1], 'Gallery'] nand2_x1
Xzero_x1[2] vdd vss zero_x1[2].[_InstanceNet[zero], 'Gallery'] zero_x1
Xnand4_x0[0] vdd vss nand4_x0[0].[_InstanceNet[nq], 'Gallery'] nand4_x0[0].[_InstanceNet[i0], 'Gallery'] nand4_x0[0].[_InstanceNet[i1], 'Gallery'] nand4_x0[0].[_InstanceNet[i2], 'Gallery'] nand4_x0[0].[_InstanceNet[i3], 'Gallery'] nand4_x0
Xnand2_x0[1] vdd vss nand2_x0[1].[_InstanceNet[nq], 'Gallery'] nand2_x0[1].[_InstanceNet[i0], 'Gallery'] nand2_x0[1].[_InstanceNet[i1], 'Gallery'] nand2_x0
Xnor4_x1[2] vdd vss nor4_x1[2].[_InstanceNet[nq], 'Gallery'] nor4_x1[2].[_InstanceNet[i0], 'Gallery'] nor4_x1[2].[_InstanceNet[i1], 'Gallery'] nor4_x1[2].[_InstanceNet[i2], 'Gallery'] nor4_x1[2].[_InstanceNet[i3], 'Gallery'] nor4_x1
Xnand4_x1[0] vdd vss nand4_x1[0].[_InstanceNet[nq], 'Gallery'] nand4_x1[0].[_InstanceNet[i0], 'Gallery'] nand4_x1[0].[_InstanceNet[i1], 'Gallery'] nand4_x1[0].[_InstanceNet[i2], 'Gallery'] nand4_x1[0].[_InstanceNet[i3], 'Gallery'] nand4_x1
Xbuf_x4[1] vdd vss buf_x4[1].[_InstanceNet[i], 'Gallery'] buf_x4[1].[_InstanceNet[q], 'Gallery'] buf_x4
Xone_x1[2] vdd vss one_x1[2].[_InstanceNet[one], 'Gallery'] one_x1
Xand2_x1[0] vdd vss and2_x1[0].[_InstanceNet[q], 'Gallery'] and2_x1[0].[_InstanceNet[i0], 'Gallery'] and2_x1[0].[_InstanceNet[i1], 'Gallery'] and2_x1
Xbuf_x2[1] vdd vss buf_x2[1].[_InstanceNet[i], 'Gallery'] buf_x2[1].[_InstanceNet[q], 'Gallery'] buf_x2
Xnor4_x0[2] vdd vss nor4_x0[2].[_InstanceNet[nq], 'Gallery'] nor4_x0[2].[_InstanceNet[i0], 'Gallery'] nor4_x0[2].[_InstanceNet[i1], 'Gallery'] nor4_x0[2].[_InstanceNet[i2], 'Gallery'] nor4_x0[2].[_InstanceNet[i3], 'Gallery'] nor4_x0
Xand3_x1[0] vdd vss and3_x1[0].[_InstanceNet[q], 'Gallery'] and3_x1[0].[_InstanceNet[i0], 'Gallery'] and3_x1[0].[_InstanceNet[i1], 'Gallery'] and3_x1[0].[_InstanceNet[i2], 'Gallery'] and3_x1
Xbuf_x1[1] vdd vss buf_x1[1].[_InstanceNet[i], 'Gallery'] buf_x1[1].[_InstanceNet[q], 'Gallery'] buf_x1
Xzeroone_x1[2] vdd vss zeroone_x1[2].[_InstanceNet[one], 'Gallery'] zeroone_x1[2].[_InstanceNet[zero], 'Gallery'] zeroone_x1
Xand4_x1[0] vdd vss and4_x1[0].[_InstanceNet[q], 'Gallery'] and4_x1[0].[_InstanceNet[i0], 'Gallery'] and4_x1[0].[_InstanceNet[i1], 'Gallery'] and4_x1[0].[_InstanceNet[i2], 'Gallery'] and4_x1[0].[_InstanceNet[i3], 'Gallery'] and4_x1
Xinv_x4[1] vdd vss inv_x4[1].[_InstanceNet[i], 'Gallery'] inv_x4[1].[_InstanceNet[nq], 'Gallery'] inv_x4
Xnor3_x1[2] vdd vss nor3_x1[2].[_InstanceNet[nq], 'Gallery'] nor3_x1[2].[_InstanceNet[i0], 'Gallery'] nor3_x1[2].[_InstanceNet[i1], 'Gallery'] nor3_x1[2].[_InstanceNet[i2], 'Gallery'] nor3_x1
Xnor2_x0[0] vdd vss nor2_x0[0].[_InstanceNet[nq], 'Gallery'] nor2_x0[0].[_InstanceNet[i0], 'Gallery'] nor2_x0[0].[_InstanceNet[i1], 'Gallery'] nor2_x0
Xinv_x2[1] vdd vss inv_x2[1].[_InstanceNet[i], 'Gallery'] inv_x2[1].[_InstanceNet[nq], 'Gallery'] inv_x2
Xdecap_w0[2] vdd vss decap_w0
Xnor2_x1[0] vdd vss nor2_x1[0].[_InstanceNet[nq], 'Gallery'] nor2_x1[0].[_InstanceNet[i0], 'Gallery'] nor2_x1[0].[_InstanceNet[i1], 'Gallery'] nor2_x1
Xinv_x1[1] vdd vss inv_x1[1].[_InstanceNet[i], 'Gallery'] inv_x1[1].[_InstanceNet[nq], 'Gallery'] inv_x1
Xnor3_x0[2] vdd vss nor3_x0[2].[_InstanceNet[nq], 'Gallery'] nor3_x0[2].[_InstanceNet[i0], 'Gallery'] nor3_x0[2].[_InstanceNet[i1], 'Gallery'] nor3_x0[2].[_InstanceNet[i2], 'Gallery'] nor3_x0
Xnor3_x0[0] vdd vss nor3_x0[0].[_InstanceNet[nq], 'Gallery'] nor3_x0[0].[_InstanceNet[i0], 'Gallery'] nor3_x0[0].[_InstanceNet[i1], 'Gallery'] nor3_x0[0].[_InstanceNet[i2], 'Gallery'] nor3_x0
Xinv_x0[1] vdd vss inv_x0[1].[_InstanceNet[i], 'Gallery'] inv_x0[1].[_InstanceNet[nq], 'Gallery'] inv_x0
Xinv_x0[2] vdd vss inv_x0[2].[_InstanceNet[i], 'Gallery'] inv_x0[2].[_InstanceNet[nq], 'Gallery'] inv_x0
Xnor3_x1[0] vdd vss nor3_x1[0].[_InstanceNet[nq], 'Gallery'] nor3_x1[0].[_InstanceNet[i0], 'Gallery'] nor3_x1[0].[_InstanceNet[i1], 'Gallery'] nor3_x1[0].[_InstanceNet[i2], 'Gallery'] nor3_x1
Xdecap_w0[1] vdd vss decap_w0
Xnor2_x1[2] vdd vss nor2_x1[2].[_InstanceNet[nq], 'Gallery'] nor2_x1[2].[_InstanceNet[i0], 'Gallery'] nor2_x1[2].[_InstanceNet[i1], 'Gallery'] nor2_x1
Xnor4_x0[0] vdd vss nor4_x0[0].[_InstanceNet[nq], 'Gallery'] nor4_x0[0].[_InstanceNet[i0], 'Gallery'] nor4_x0[0].[_InstanceNet[i1], 'Gallery'] nor4_x0[0].[_InstanceNet[i2], 'Gallery'] nor4_x0[0].[_InstanceNet[i3], 'Gallery'] nor4_x0
Xzeroone_x1[1] vdd vss zeroone_x1[1].[_InstanceNet[one], 'Gallery'] zeroone_x1[1].[_InstanceNet[zero], 'Gallery'] zeroone_x1
Xinv_x1[2] vdd vss inv_x1[2].[_InstanceNet[i], 'Gallery'] inv_x1[2].[_InstanceNet[nq], 'Gallery'] inv_x1
Xnor4_x1[0] vdd vss nor4_x1[0].[_InstanceNet[nq], 'Gallery'] nor4_x1[0].[_InstanceNet[i0], 'Gallery'] nor4_x1[0].[_InstanceNet[i1], 'Gallery'] nor4_x1[0].[_InstanceNet[i2], 'Gallery'] nor4_x1[0].[_InstanceNet[i3], 'Gallery'] nor4_x1
Xone_x1[1] vdd vss one_x1[1].[_InstanceNet[one], 'Gallery'] one_x1
Xnor2_x0[2] vdd vss nor2_x0[2].[_InstanceNet[nq], 'Gallery'] nor2_x0[2].[_InstanceNet[i0], 'Gallery'] nor2_x0[2].[_InstanceNet[i1], 'Gallery'] nor2_x0
Xor2_x1[0] vdd vss or2_x1[0].[_InstanceNet[q], 'Gallery'] or2_x1[0].[_InstanceNet[i0], 'Gallery'] or2_x1[0].[_InstanceNet[i1], 'Gallery'] or2_x1
Xzero_x1[1] vdd vss zero_x1[1].[_InstanceNet[zero], 'Gallery'] zero_x1
Xinv_x2[2] vdd vss inv_x2[2].[_InstanceNet[i], 'Gallery'] inv_x2[2].[_InstanceNet[nq], 'Gallery'] inv_x2
Xor3_x1[0] vdd vss or3_x1[0].[_InstanceNet[q], 'Gallery'] or3_x1[0].[_InstanceNet[i0], 'Gallery'] or3_x1[0].[_InstanceNet[i1], 'Gallery'] or3_x1[0].[_InstanceNet[i2], 'Gallery'] or3_x1
Xdiode_w1[1] vdd vss diode_w1[1].[_InstanceNet[i], 'Gallery'] diode_w1
Xand4_x1[2] vdd vss and4_x1[2].[_InstanceNet[q], 'Gallery'] and4_x1[2].[_InstanceNet[i0], 'Gallery'] and4_x1[2].[_InstanceNet[i1], 'Gallery'] and4_x1[2].[_InstanceNet[i2], 'Gallery'] and4_x1[2].[_InstanceNet[i3], 'Gallery'] and4_x1
Xor4_x1[0] vdd vss or4_x1[0].[_InstanceNet[q], 'Gallery'] or4_x1[0].[_InstanceNet[i0], 'Gallery'] or4_x1[0].[_InstanceNet[i1], 'Gallery'] or4_x1[0].[_InstanceNet[i2], 'Gallery'] or4_x1[0].[_InstanceNet[i3], 'Gallery'] or4_x1
Xtie_poly_w4[1] vdd vss tie_poly_w4
Xinv_x4[2] vdd vss inv_x4[2].[_InstanceNet[i], 'Gallery'] inv_x4[2].[_InstanceNet[nq], 'Gallery'] inv_x4
Xmux2_x1[0] vdd vss mux2_x1[0].[_InstanceNet[i0], 'Gallery'] mux2_x1[0].[_InstanceNet[i1], 'Gallery'] mux2_x1[0].[_InstanceNet[cmd], 'Gallery'] mux2_x1[0].[_InstanceNet[q], 'Gallery'] mux2_x1
Xtie_diff_w4[1] vdd vss tie_diff_w4
Xand3_x1[2] vdd vss and3_x1[2].[_InstanceNet[q], 'Gallery'] and3_x1[2].[_InstanceNet[i0], 'Gallery'] and3_x1[2].[_InstanceNet[i1], 'Gallery'] and3_x1[2].[_InstanceNet[i2], 'Gallery'] and3_x1
Xand21nor_x0[0] vdd vss and21nor_x0[0].[_InstanceNet[nq], 'Gallery'] and21nor_x0[0].[_InstanceNet[i0], 'Gallery'] and21nor_x0[0].[_InstanceNet[i1], 'Gallery'] and21nor_x0[0].[_InstanceNet[i2], 'Gallery'] and21nor_x0
Xtie_w4[1] vdd vss tie_w4
Xbuf_x1[2] vdd vss buf_x1[2].[_InstanceNet[i], 'Gallery'] buf_x1[2].[_InstanceNet[q], 'Gallery'] buf_x1
Xand21nor_x1[0] vdd vss and21nor_x1[0].[_InstanceNet[nq], 'Gallery'] and21nor_x1[0].[_InstanceNet[i0], 'Gallery'] and21nor_x1[0].[_InstanceNet[i1], 'Gallery'] and21nor_x1[0].[_InstanceNet[i2], 'Gallery'] and21nor_x1
Xfill_w4[1] vdd vss fill_w4
Xand2_x1[2] vdd vss and2_x1[2].[_InstanceNet[q], 'Gallery'] and2_x1[2].[_InstanceNet[i0], 'Gallery'] and2_x1[2].[_InstanceNet[i1], 'Gallery'] and2_x1
Xor21nand_x0[0] vdd vss or21nand_x0[0].[_InstanceNet[nq], 'Gallery'] or21nand_x0[0].[_InstanceNet[i0], 'Gallery'] or21nand_x0[0].[_InstanceNet[i1], 'Gallery'] or21nand_x0[0].[_InstanceNet[i2], 'Gallery'] or21nand_x0
Xtie_poly_w2[1] vdd vss tie_poly_w2
Xbuf_x2[2] vdd vss buf_x2[2].[_InstanceNet[i], 'Gallery'] buf_x2[2].[_InstanceNet[q], 'Gallery'] buf_x2
Xor21nand_x1[0] vdd vss or21nand_x1[0].[_InstanceNet[nq], 'Gallery'] or21nand_x1[0].[_InstanceNet[i0], 'Gallery'] or21nand_x1[0].[_InstanceNet[i1], 'Gallery'] or21nand_x1[0].[_InstanceNet[i2], 'Gallery'] or21nand_x1
Xtie_diff_w2[1] vdd vss tie_diff_w2
Xnand4_x1[2] vdd vss nand4_x1[2].[_InstanceNet[nq], 'Gallery'] nand4_x1[2].[_InstanceNet[i0], 'Gallery'] nand4_x1[2].[_InstanceNet[i1], 'Gallery'] nand4_x1[2].[_InstanceNet[i2], 'Gallery'] nand4_x1[2].[_InstanceNet[i3], 'Gallery'] nand4_x1
Xxor2_x0[0] vdd vss xor2_x0[0].[_InstanceNet[i0], 'Gallery'] xor2_x0[0].[_InstanceNet[i1], 'Gallery'] xor2_x0[0].[_InstanceNet[q], 'Gallery'] xor2_x0
Xtie_w2[1] vdd vss tie_w2
Xbuf_x4[2] vdd vss buf_x4[2].[_InstanceNet[i], 'Gallery'] buf_x4[2].[_InstanceNet[q], 'Gallery'] buf_x4
Xnexor2_x0[0] vdd vss nexor2_x0[0].[_InstanceNet[i0], 'Gallery'] nexor2_x0[0].[_InstanceNet[i1], 'Gallery'] nexor2_x0[0].[_InstanceNet[nq], 'Gallery'] nexor2_x0
Xfill_w2[1] vdd vss fill_w2
Xnand4_x0[2] vdd vss nand4_x0[2].[_InstanceNet[nq], 'Gallery'] nand4_x0[2].[_InstanceNet[i0], 'Gallery'] nand4_x0[2].[_InstanceNet[i1], 'Gallery'] nand4_x0[2].[_InstanceNet[i2], 'Gallery'] nand4_x0[2].[_InstanceNet[i3], 'Gallery'] nand4_x0
Xnsnrlatch_x0[0] vdd vss nsnrlatch_x0[0].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x0[0].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x0[0].[_InstanceNet[q], 'Gallery'] nsnrlatch_x0[0].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x0
Xtie_poly[1] vdd vss tie_poly
Xnand2_x0[2] vdd vss nand2_x0[2].[_InstanceNet[nq], 'Gallery'] nand2_x0[2].[_InstanceNet[i0], 'Gallery'] nand2_x0[2].[_InstanceNet[i1], 'Gallery'] nand2_x0
Xnsnrlatch_x1[0] vdd vss nsnrlatch_x1[0].[_InstanceNet[nset], 'Gallery'] nsnrlatch_x1[0].[_InstanceNet[nrst], 'Gallery'] nsnrlatch_x1[0].[_InstanceNet[q], 'Gallery'] nsnrlatch_x1[0].[_InstanceNet[nq], 'Gallery'] nsnrlatch_x1
Xtie_diff[1] vdd vss tie_diff
Xnand3_x1[2] vdd vss nand3_x1[2].[_InstanceNet[nq], 'Gallery'] nand3_x1[2].[_InstanceNet[i0], 'Gallery'] nand3_x1[2].[_InstanceNet[i1], 'Gallery'] nand3_x1[2].[_InstanceNet[i2], 'Gallery'] nand3_x1
Xdff_x1[0] vdd vss dff_x1[0].[_InstanceNet[i], 'Gallery'] dff_x1[0].[_InstanceNet[clk], 'Gallery'] dff_x1[0].[_InstanceNet[q], 'Gallery'] dff_x1
Xtie[1] vdd vss tie
Xnand2_x1[2] vdd vss nand2_x1[2].[_InstanceNet[nq], 'Gallery'] nand2_x1[2].[_InstanceNet[i0], 'Gallery'] nand2_x1[2].[_InstanceNet[i1], 'Gallery'] nand2_x1
Xdffnr_x1[0] vdd vss dffnr_x1[0].[_InstanceNet[i], 'Gallery'] dffnr_x1[0].[_InstanceNet[clk], 'Gallery'] dffnr_x1[0].[_InstanceNet[q], 'Gallery'] dffnr_x1[0].[_InstanceNet[nrst], 'Gallery'] dffnr_x1
Xfill[1] vdd vss fill
Xnand3_x0[2] vdd vss nand3_x0[2].[_InstanceNet[nq], 'Gallery'] nand3_x0[2].[_InstanceNet[i0], 'Gallery'] nand3_x0[2].[_InstanceNet[i1], 'Gallery'] nand3_x0[2].[_InstanceNet[i2], 'Gallery'] nand3_x0
.ends Gallery
