* BulkConn_200WNoUp
.subckt BulkConn_200WNoUp vdd vss iovdd iovss

.ends BulkConn_200WNoUp
