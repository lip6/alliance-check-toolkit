********************************************************************************
* sram2bw2r2.cir
* ngspice simulation
* lsxram
********************************************************************************

.option  nopage nomod
+        newtol numdgt=7 ingold=2 gmindc=1e-18
.option DOTNODE
.option MSGNODE = 0

********************************************************************************
* BSIM4 transistor model parameters for ngspice and simulation conditions
********************************************************************************

.lib _TECHNO _MODEL
.TEMP _TEMP
Vground vss 0 0
Vsupply vdd 0 DC _VDD
gfoncd vdd 0 vdd 0 1.0e-15

********************************************************************************
* Circuit Instantiation with loading output
********************************************************************************
.INCLUDE ../spi/sram2bw2r2.spi
*.subckt sram2bw2r2 at0 at1 ax ay az0 az1 ck it iz nqx nqy vdd vss 

Xa at0 at1 ax ay az0 az1 ck it iz nqx nqy vdd vss sram2bw2r2 
*Cload q vss 0.0020pF

********************************************************************************
* input stimluli and transient analysis
********************************************************************************

vck  ck  vss dc 0.8 pulse (0 _VDD 1000ps 30ps 30ps 970ps 2000ps)
vit  it  vss dc 0.8 pulse (0 _VDD 500ps 30ps 30ps 1970ps 4000ps)
viz  iz  vss dc 0

vat0 at0 vss dc _VDD
vaz0 az0 vss dc 0

vat1 at1 vss dc 0
vaz1 az1 vss dc 0

vax  ax  vss dc 0
vay  ay  vss dc 0

.control
TRAN 1ps 24ns 0 

set width=110

meas tran proptimeRF TRIG v(ck) val=0.9 RISE=1 TARG v(q) VAL=0.9 FALL=1
meas tran proptimeFR TRIG v(ck) val=0.9 FALL=1 TARG v(q) VAL=0.9 RISE=1

gnuplot sram2bw2r2/sram2bw2r2._MODEL v(ck) v(it) v(nqx)
+ title 'input and output of the sff1_x4'
+ xlabel 'time / s' ylabel 'Voltage / V' 

.endc

.end
