* pnp_f
.param
+ dkispp=1.1857e+00 dkbfpp=1.4174e+00 dknfpp=1.000
+ dkispp5x=1.2104e+00 dkbfpp5x=1.7922e+00 dknfpp5x=1.0009e+00 dkisepp5x=6.4618e-01
