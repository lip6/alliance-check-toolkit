* or21nand_x1
* or21nand_x1
.subckt or21nand_x1 vdd vss nq i0 i1 i2
Mi0_nmos _net0 i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi0_pmos vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
Mi1_nmos vss i1 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi1_pmos _net1 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
Mi2_nmos _net0 i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi2_pmos nq i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
.ends or21nand_x1
