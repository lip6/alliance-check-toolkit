* diode_tt
.param
+ sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult=9.8286e-01 
+ sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult=9.8954e-01 
+ sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult=1.0116e+0 
+ sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult=9.8200e-01 
+ sky130_fd_pr__nfet_01v8__ajunction_mult=9.9543e-1
+ sky130_fd_pr__nfet_01v8__pjunction_mult=1.0204e+0
+ sky130_fd_pr__pfet_01v8__ajunction_mult=9.9626e-1
+ sky130_fd_pr__pfet_01v8__pjunction_mult=1.0009e+0
