* DP8TBlock_512x64_8WE
.subckt DP8TBlock_512x64_8WE clk1 clk2 a1[0] a2[0] a1[1] a2[1] a1[2] a2[2] a1[3] a2[3] a1[4] a2[4] a1[5] a2[5] a1[6] a2[6] a1[7] a2[7] a1[8] a2[8] vss vdd q1[0] q1[1] q1[2] q1[3] q1[4] q1[5] q1[6] q1[7] q1[8] q1[9] q1[10] q1[11] q1[12] q1[13] q1[14] q1[15] q1[16] q1[17] q1[18] q1[19] q1[20] q1[21] q1[22] q1[23] q1[24] q1[25] q1[26] q1[27] q1[28] q1[29] q1[30] q1[31] q1[32] q1[33] q1[34] q1[35] q1[36] q1[37] q1[38] q1[39] q1[40] q1[41] q1[42] q1[43] q1[44] q1[45] q1[46] q1[47] q1[48] q1[49] q1[50] q1[51] q1[52] q1[53] q1[54] q1[55] q1[56] q1[57] q1[58] q1[59] q1[60] q1[61] q1[62] q1[63] q2[0] q2[1] q2[2] q2[3] q2[4] q2[5] q2[6] q2[7] q2[8] q2[9] q2[10] q2[11] q2[12] q2[13] q2[14] q2[15] q2[16] q2[17] q2[18] q2[19] q2[20] q2[21] q2[22] q2[23] q2[24] q2[25] q2[26] q2[27] q2[28] q2[29] q2[30] q2[31] q2[32] q2[33] q2[34] q2[35] q2[36] q2[37] q2[38] q2[39] q2[40] q2[41] q2[42] q2[43] q2[44] q2[45] q2[46] q2[47] q2[48] q2[49] q2[50] q2[51] q2[52] q2[53] q2[54] q2[55] q2[56] q2[57] q2[58] q2[59] q2[60] q2[61] q2[62] q2[63] d1[0] d1[1] d1[2] d1[3] d1[4] d1[5] d1[6] d1[7] d1[8] d1[9] d1[10] d1[11] d1[12] d1[13] d1[14] d1[15] d1[16] d1[17] d1[18] d1[19] d1[20] d1[21] d1[22] d1[23] d1[24] d1[25] d1[26] d1[27] d1[28] d1[29] d1[30] d1[31] d1[32] d1[33] d1[34] d1[35] d1[36] d1[37] d1[38] d1[39] d1[40] d1[41] d1[42] d1[43] d1[44] d1[45] d1[46] d1[47] d1[48] d1[49] d1[50] d1[51] d1[52] d1[53] d1[54] d1[55] d1[56] d1[57] d1[58] d1[59] d1[60] d1[61] d1[62] d1[63] d2[0] d2[1] d2[2] d2[3] d2[4] d2[5] d2[6] d2[7] d2[8] d2[9] d2[10] d2[11] d2[12] d2[13] d2[14] d2[15] d2[16] d2[17] d2[18] d2[19] d2[20] d2[21] d2[22] d2[23] d2[24] d2[25] d2[26] d2[27] d2[28] d2[29] d2[30] d2[31] d2[32] d2[33] d2[34] d2[35] d2[36] d2[37] d2[38] d2[39] d2[40] d2[41] d2[42] d2[43] d2[44] d2[45] d2[46] d2[47] d2[48] d2[49] d2[50] d2[51] d2[52] d2[53] d2[54] d2[55] d2[56] d2[57] d2[58] d2[59] d2[60] d2[61] d2[62] d2[63] we1[0] we1[1] we1[2] we1[3] we1[4] we1[5] we1[6] we1[7] we2[0] we2[1] we2[2] we2[3] we2[4] we2[5] we2[6] we2[7]
Xrowperiph1 vss vdd clk1 a1[0] a1[1] a1[2] a1[3] a1[4] a1[5] a1[6] a1[7] a1[8] wl1[0] wl1[1] wl1[2] wl1[3] wl1[4] wl1[5] wl1[6] wl1[7] wl1[8] wl1[9] wl1[10] wl1[11] wl1[12] wl1[13] wl1[14] wl1[15] wl1[16] wl1[17] wl1[18] wl1[19] wl1[20] wl1[21] wl1[22] wl1[23] wl1[24] wl1[25] wl1[26] wl1[27] wl1[28] wl1[29] wl1[30] wl1[31] wl1[32] wl1[33] wl1[34] wl1[35] wl1[36] wl1[37] wl1[38] wl1[39] wl1[40] wl1[41] wl1[42] wl1[43] wl1[44] wl1[45] wl1[46] wl1[47] wl1[48] wl1[49] wl1[50] wl1[51] wl1[52] wl1[53] wl1[54] wl1[55] wl1[56] wl1[57] wl1[58] wl1[59] wl1[60] wl1[61] wl1[62] wl1[63] wl1[64] wl1[65] wl1[66] wl1[67] wl1[68] wl1[69] wl1[70] wl1[71] wl1[72] wl1[73] wl1[74] wl1[75] wl1[76] wl1[77] wl1[78] wl1[79] wl1[80] wl1[81] wl1[82] wl1[83] wl1[84] wl1[85] wl1[86] wl1[87] wl1[88] wl1[89] wl1[90] wl1[91] wl1[92] wl1[93] wl1[94] wl1[95] wl1[96] wl1[97] wl1[98] wl1[99] wl1[100] wl1[101] wl1[102] wl1[103] wl1[104] wl1[105] wl1[106] wl1[107] wl1[108] wl1[109] wl1[110] wl1[111] wl1[112] wl1[113] wl1[114] wl1[115] wl1[116] wl1[117] wl1[118] wl1[119] wl1[120] wl1[121] wl1[122] wl1[123] wl1[124] wl1[125] wl1[126] wl1[127] mux1[0] mux1[1] mux1[2] mux1[3] columnclk1 precharge1_n we_en1 DP8TRowPeriphery_3_4_2_wl1
Xrowperiph2 vss vdd clk2 a2[0] a2[1] a2[2] a2[3] a2[4] a2[5] a2[6] a2[7] a2[8] wl2[0] wl2[1] wl2[2] wl2[3] wl2[4] wl2[5] wl2[6] wl2[7] wl2[8] wl2[9] wl2[10] wl2[11] wl2[12] wl2[13] wl2[14] wl2[15] wl2[16] wl2[17] wl2[18] wl2[19] wl2[20] wl2[21] wl2[22] wl2[23] wl2[24] wl2[25] wl2[26] wl2[27] wl2[28] wl2[29] wl2[30] wl2[31] wl2[32] wl2[33] wl2[34] wl2[35] wl2[36] wl2[37] wl2[38] wl2[39] wl2[40] wl2[41] wl2[42] wl2[43] wl2[44] wl2[45] wl2[46] wl2[47] wl2[48] wl2[49] wl2[50] wl2[51] wl2[52] wl2[53] wl2[54] wl2[55] wl2[56] wl2[57] wl2[58] wl2[59] wl2[60] wl2[61] wl2[62] wl2[63] wl2[64] wl2[65] wl2[66] wl2[67] wl2[68] wl2[69] wl2[70] wl2[71] wl2[72] wl2[73] wl2[74] wl2[75] wl2[76] wl2[77] wl2[78] wl2[79] wl2[80] wl2[81] wl2[82] wl2[83] wl2[84] wl2[85] wl2[86] wl2[87] wl2[88] wl2[89] wl2[90] wl2[91] wl2[92] wl2[93] wl2[94] wl2[95] wl2[96] wl2[97] wl2[98] wl2[99] wl2[100] wl2[101] wl2[102] wl2[103] wl2[104] wl2[105] wl2[106] wl2[107] wl2[108] wl2[109] wl2[110] wl2[111] wl2[112] wl2[113] wl2[114] wl2[115] wl2[116] wl2[117] wl2[118] wl2[119] wl2[120] wl2[121] wl2[122] wl2[123] wl2[124] wl2[125] wl2[126] wl2[127] mux2[0] mux2[1] mux2[2] mux2[3] columnclk2 precharge2_n we_en2 DP8TRowPeriphery_3_4_2_wl2
Xcolumnblock vss vdd columnclk1 columnclk2 precharge1_n precharge2_n we_en1 we_en2 wl1[0] wl1[1] wl1[2] wl1[3] wl1[4] wl1[5] wl1[6] wl1[7] wl1[8] wl1[9] wl1[10] wl1[11] wl1[12] wl1[13] wl1[14] wl1[15] wl1[16] wl1[17] wl1[18] wl1[19] wl1[20] wl1[21] wl1[22] wl1[23] wl1[24] wl1[25] wl1[26] wl1[27] wl1[28] wl1[29] wl1[30] wl1[31] wl1[32] wl1[33] wl1[34] wl1[35] wl1[36] wl1[37] wl1[38] wl1[39] wl1[40] wl1[41] wl1[42] wl1[43] wl1[44] wl1[45] wl1[46] wl1[47] wl1[48] wl1[49] wl1[50] wl1[51] wl1[52] wl1[53] wl1[54] wl1[55] wl1[56] wl1[57] wl1[58] wl1[59] wl1[60] wl1[61] wl1[62] wl1[63] wl1[64] wl1[65] wl1[66] wl1[67] wl1[68] wl1[69] wl1[70] wl1[71] wl1[72] wl1[73] wl1[74] wl1[75] wl1[76] wl1[77] wl1[78] wl1[79] wl1[80] wl1[81] wl1[82] wl1[83] wl1[84] wl1[85] wl1[86] wl1[87] wl1[88] wl1[89] wl1[90] wl1[91] wl1[92] wl1[93] wl1[94] wl1[95] wl1[96] wl1[97] wl1[98] wl1[99] wl1[100] wl1[101] wl1[102] wl1[103] wl1[104] wl1[105] wl1[106] wl1[107] wl1[108] wl1[109] wl1[110] wl1[111] wl1[112] wl1[113] wl1[114] wl1[115] wl1[116] wl1[117] wl1[118] wl1[119] wl1[120] wl1[121] wl1[122] wl1[123] wl1[124] wl1[125] wl1[126] wl1[127] wl2[0] wl2[1] wl2[2] wl2[3] wl2[4] wl2[5] wl2[6] wl2[7] wl2[8] wl2[9] wl2[10] wl2[11] wl2[12] wl2[13] wl2[14] wl2[15] wl2[16] wl2[17] wl2[18] wl2[19] wl2[20] wl2[21] wl2[22] wl2[23] wl2[24] wl2[25] wl2[26] wl2[27] wl2[28] wl2[29] wl2[30] wl2[31] wl2[32] wl2[33] wl2[34] wl2[35] wl2[36] wl2[37] wl2[38] wl2[39] wl2[40] wl2[41] wl2[42] wl2[43] wl2[44] wl2[45] wl2[46] wl2[47] wl2[48] wl2[49] wl2[50] wl2[51] wl2[52] wl2[53] wl2[54] wl2[55] wl2[56] wl2[57] wl2[58] wl2[59] wl2[60] wl2[61] wl2[62] wl2[63] wl2[64] wl2[65] wl2[66] wl2[67] wl2[68] wl2[69] wl2[70] wl2[71] wl2[72] wl2[73] wl2[74] wl2[75] wl2[76] wl2[77] wl2[78] wl2[79] wl2[80] wl2[81] wl2[82] wl2[83] wl2[84] wl2[85] wl2[86] wl2[87] wl2[88] wl2[89] wl2[90] wl2[91] wl2[92] wl2[93] wl2[94] wl2[95] wl2[96] wl2[97] wl2[98] wl2[99] wl2[100] wl2[101] wl2[102] wl2[103] wl2[104] wl2[105] wl2[106] wl2[107] wl2[108] wl2[109] wl2[110] wl2[111] wl2[112] wl2[113] wl2[114] wl2[115] wl2[116] wl2[117] wl2[118] wl2[119] wl2[120] wl2[121] wl2[122] wl2[123] wl2[124] wl2[125] wl2[126] wl2[127] mux1[0] mux1[1] mux1[2] mux1[3] mux2[0] mux2[1] mux2[2] mux2[3] we1[0] we2[0] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1[1] we2[1] q1[8] q2[8] d1[8] d2[8] q1[9] q2[9] d1[9] d2[9] q1[10] q2[10] d1[10] d2[10] q1[11] q2[11] d1[11] d2[11] q1[12] q2[12] d1[12] d2[12] q1[13] q2[13] d1[13] d2[13] q1[14] q2[14] d1[14] d2[14] q1[15] q2[15] d1[15] d2[15] we1[2] we2[2] q1[16] q2[16] d1[16] d2[16] q1[17] q2[17] d1[17] d2[17] q1[18] q2[18] d1[18] d2[18] q1[19] q2[19] d1[19] d2[19] q1[20] q2[20] d1[20] d2[20] q1[21] q2[21] d1[21] d2[21] q1[22] q2[22] d1[22] d2[22] q1[23] q2[23] d1[23] d2[23] we1[3] we2[3] q1[24] q2[24] d1[24] d2[24] q1[25] q2[25] d1[25] d2[25] q1[26] q2[26] d1[26] d2[26] q1[27] q2[27] d1[27] d2[27] q1[28] q2[28] d1[28] d2[28] q1[29] q2[29] d1[29] d2[29] q1[30] q2[30] d1[30] d2[30] q1[31] q2[31] d1[31] d2[31] we1[4] we2[4] q1[32] q2[32] d1[32] d2[32] q1[33] q2[33] d1[33] d2[33] q1[34] q2[34] d1[34] d2[34] q1[35] q2[35] d1[35] d2[35] q1[36] q2[36] d1[36] d2[36] q1[37] q2[37] d1[37] d2[37] q1[38] q2[38] d1[38] d2[38] q1[39] q2[39] d1[39] d2[39] we1[5] we2[5] q1[40] q2[40] d1[40] d2[40] q1[41] q2[41] d1[41] d2[41] q1[42] q2[42] d1[42] d2[42] q1[43] q2[43] d1[43] d2[43] q1[44] q2[44] d1[44] d2[44] q1[45] q2[45] d1[45] d2[45] q1[46] q2[46] d1[46] d2[46] q1[47] q2[47] d1[47] d2[47] we1[6] we2[6] q1[48] q2[48] d1[48] d2[48] q1[49] q2[49] d1[49] d2[49] q1[50] q2[50] d1[50] d2[50] q1[51] q2[51] d1[51] d2[51] q1[52] q2[52] d1[52] d2[52] q1[53] q2[53] d1[53] d2[53] q1[54] q2[54] d1[54] d2[54] q1[55] q2[55] d1[55] d2[55] we1[7] we2[7] q1[56] q2[56] d1[56] d2[56] q1[57] q2[57] d1[57] d2[57] q1[58] q2[58] d1[58] d2[58] q1[59] q2[59] d1[59] d2[59] q1[60] q2[60] d1[60] d2[60] q1[61] q2[61] d1[61] d2[61] q1[62] q2[62] d1[62] d2[62] q1[63] q2[63] d1[63] d2[63] DP8TColumnBlock_128R64B4M8W
.ends DP8TBlock_512x64_8WE
