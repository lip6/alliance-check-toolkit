* Spice description of no2_x1
* Spice driver version -780419301
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:00

* INTERF i0 i1 nq vdd vss 


.subckt no2_x1 3 4 5 2 6 
* NET 2 = vdd
* NET 3 = i0
* NET 4 = i1
* NET 5 = nq
* NET 6 = vss
Mtr_00004 1 4 5 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00003 2 3 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00002 6 3 5 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00001 5 4 6 6 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
C5 2 6 1.17336e-15
C4 3 6 2.1784e-15
C3 4 6 2.10538e-15
C2 5 6 2.27334e-15
C1 6 6 1.40651e-15
.ends no2_x1

