* GuardRing_N1270W450HTF
* GuardRing_N1270W450HTF
.subckt GuardRing_N1270W450HTF conn

.ends GuardRing_N1270W450HTF
