* Gallery
* GuardRing_N1270W450HTF
.subckt GuardRing_N1270W450HTF conn

.ends GuardRing_N1270W450HTF
* GuardRing_P418W1550HFF
.subckt GuardRing_P418W1550HFF conn

.ends GuardRing_P418W1550HFF
* GuardRing_P632W1550HFF
.subckt GuardRing_P632W1550HFF conn

.ends GuardRing_P632W1550HFF
* GuardRing_N8666W2488HTT
.subckt GuardRing_N8666W2488HTT conn

.ends GuardRing_N8666W2488HTT
* GuardRing_P18000W3888HFT
.subckt GuardRing_P18000W3888HFT conn

.ends GuardRing_P18000W3888HFT
* nand2_x1
.subckt nand2_x1 vdd vss nq i0 i1
Mi0_nmos vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi0_pmos vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
Mi1_nmos _net0 i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi1_pmos nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
.ends nand2_x1
* LevelUp
.subckt LevelUp vdd iovdd vss i o
Mn_i_inv i_n i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.46um
Mp_i_inv i_n i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.56um
Mn_lvld_n vss i lvld_n vss sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=2.4um
Mn_lvld lvld i_n vss vss sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=2.4um
Mp_lvld_n iovdd lvld lvld_n iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=0.42um
Mp_lvld lvld lvld_n iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=0.42um
Mn_lvld_n_inv vss lvld_n o vss sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=2.4um
Mp_lvld_n_inv iovdd lvld_n o iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=4.4um
.ends LevelUp
* nor2_x1
.subckt nor2_x1 vdd vss nq i0 i1
Mi0_nmos vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi0_pmos vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
Mi1_nmos nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mi1_pmos _net0 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
.ends nor2_x1
* inv_x1
.subckt inv_x1 vdd vss i nq
Mnmos vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.535um
Mpmos vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.095um
.ends inv_x1
* tie
.subckt tie vdd vss

.ends tie
* LevelUpInv
.subckt LevelUpInv vdd iovdd vss i o
Mn_i_inv i_n i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.46um
Mp_i_inv i_n i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.56um
Mn_lvld_n vss i_n lvld_n vss sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=2.4um
Mn_lvld lvld i vss vss sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=2.4um
Mp_lvld_n iovdd lvld lvld_n iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=0.42um
Mp_lvld lvld lvld_n iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=0.42um
Mn_lvld_n_inv vss lvld_n o vss sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=2.4um
Mp_lvld_n_inv iovdd lvld_n o iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=4.4um
.ends LevelUpInv
* GuardRing_N17368W8096HTF
.subckt GuardRing_N17368W8096HTF conn

.ends GuardRing_N17368W8096HTF
* GuardRing_P18000W8728HFF
.subckt GuardRing_P18000W8728HFF conn

.ends GuardRing_P18000W8728HFF
* GuardRing_P17368W3836HFF
.subckt GuardRing_P17368W3836HFF conn

.ends GuardRing_P17368W3836HFF
* GuardRing_N18000W4468HFF
.subckt GuardRing_N18000W4468HFF conn

.ends GuardRing_N18000W4468HFF
* SecondaryProtection
.subckt SecondaryProtection iovdd iovss pad core
RR pad core 241.0
Xguard1 iovss GuardRing_P632W1550HFF
DDN iovss core sky130_fd_pr__diode_pw2nd_05v5 area=3.6875e-12 pj=13.68um
Xguard2 iovss GuardRing_P418W1550HFF
DDP core iovdd sky130_fd_pr__diode_pd2nw_05v5 area=3.6375000000000002e-12 pj=11.2um
Xguard3 iovdd GuardRing_N1270W450HTF
.ends SecondaryProtection
* Clamp_P12N0D
.subckt Clamp_P12N0D iovss iovdd pad
Mclamp_g0 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g1 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g2 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g3 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g4 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g5 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g6 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g7 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g8 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g9 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g10 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g11 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
XOuterRing iovss GuardRing_P18000W8728HFF
XInnerRing iovdd GuardRing_N17368W8096HTF
RRoff iovdd off 5502.103030303
.ends Clamp_P12N0D
* Clamp_N12N0D
.subckt Clamp_N12N0D iovss iovdd pad
Mclamp_g0 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g1 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g2 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g3 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g4 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g5 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g6 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g7 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g8 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g9 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g10 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g11 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
XOuterRing iovdd GuardRing_N18000W4468HFF
XInnerRing iovss GuardRing_P17368W3836HFF
RRoff iovss off 2391.0121212121
.ends Clamp_N12N0D
* RCClampInverter
.subckt RCClampInverter supply ground in out
Mcapmos0 ground in ground ground sky130_fd_pr__nfet_g5v0d10v5__model l=10.0um w=14.0um
Mcapmos1 ground in ground ground sky130_fd_pr__nfet_g5v0d10v5__model l=10.0um w=14.0um
Mcapmos2 ground in ground ground sky130_fd_pr__nfet_g5v0d10v5__model l=10.0um w=14.0um
Mcapmos3 ground in ground ground sky130_fd_pr__nfet_g5v0d10v5__model l=10.0um w=14.0um
Mcapmos4 ground in ground ground sky130_fd_pr__nfet_g5v0d10v5__model l=10.0um w=14.0um
Mnmos0 ground in out ground sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=14.0um
Mnmos1 out in ground ground sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=14.0um
Mnmos2 ground in out ground sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=14.0um
Mnmos3 out in ground ground sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=14.0um
Mnmos4 ground in out ground sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=14.0um
Mnmos5 out in ground ground sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=14.0um
Mnmos6 ground in out ground sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=14.0um
Xnmosguardring ground GuardRing_P18000W3888HFT
Mpmos0 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos1 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos2 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos3 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos4 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos5 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos6 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos7 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos8 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos9 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos10 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos11 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos12 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos13 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos14 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos15 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos16 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos17 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos18 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos19 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos20 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos21 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos22 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos23 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos24 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos25 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos26 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos27 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos28 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos29 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos30 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos31 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos32 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos33 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos34 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos35 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos36 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos37 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos38 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos39 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos40 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos41 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos42 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos43 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos44 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos45 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos46 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos47 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos48 supply in out supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Mpmos49 out in supply supply sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=7.0um
Xpmosguardring supply GuardRing_N8666W2488HTT
.ends RCClampInverter
* RCClampResistor
.subckt RCClampResistor pin1 pin2

.ends RCClampResistor
* Clamp_N32N32D
.subckt Clamp_N32N32D iovss iovdd pad gate
Mclamp_g0 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g1 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g2 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g3 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g4 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g5 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g6 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g7 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g8 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g9 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g10 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g11 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g12 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g13 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g14 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g15 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g16 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g17 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g18 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g19 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g20 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g21 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g22 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g23 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g24 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g25 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g26 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g27 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g28 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g29 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g30 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g31 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
XOuterRing iovdd GuardRing_N18000W4468HFF
XInnerRing iovss GuardRing_P17368W3836HFF
DDGATE iovss gate sky130_fd_pr__diode_pw2nd_05v5 area=1.875e-13 pj=2.0um
.ends Clamp_N32N32D
* GateDecode
.subckt GateDecode vdd vss iovdd core en ngate pgate
Xtieinst vdd vss tie
Xen_inv vdd vss en en_n inv_x1
Xngate_nor vdd vss ngate_core core en_n nor2_x1
Xngate_levelup vdd iovdd vss ngate_core ngate LevelUp
Xpgate_nand vdd vss pgate_core core en nand2_x1
Xpgate_levelup vdd iovdd vss pgate_core pgate LevelUp
.ends GateDecode
* GateLevelUpInv
.subckt GateLevelUpInv vdd vss iovdd core ngate pgate
Xngate_levelup vdd iovdd vss core ngate LevelUpInv
Xpgate_levelup vdd iovdd vss core pgate LevelUpInv
.ends GateLevelUpInv
* Clamp_P32N4D
.subckt Clamp_P32N4D iovss iovdd pad gate
Mclamp_g0 iovdd gate pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g1 pad gate iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g2 iovdd gate pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g3 pad gate iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g4 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g5 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g6 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g7 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g8 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g9 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g10 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g11 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g12 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g13 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g14 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g15 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g16 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g17 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g18 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g19 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g20 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g21 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g22 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g23 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g24 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g25 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g26 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g27 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g28 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g29 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g30 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g31 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
XOuterRing iovss GuardRing_P18000W8728HFF
XInnerRing iovdd GuardRing_N17368W8096HTF
DDGATE gate iovdd sky130_fd_pr__diode_pd2nw_05v5 area=1.875e-13 pj=2.0um
RRoff iovdd off 5502.103030303
.ends Clamp_P32N4D
* Clamp_N32N4D
.subckt Clamp_N32N4D iovss iovdd pad gate
Mclamp_g0 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g1 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g2 iovss gate pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g3 pad gate iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g4 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g5 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g6 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g7 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g8 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g9 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g10 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g11 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g12 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g13 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g14 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g15 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g16 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g17 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g18 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g19 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g20 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g21 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g22 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g23 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g24 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g25 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g26 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g27 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g28 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g29 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g30 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g31 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
XOuterRing iovdd GuardRing_N18000W4468HFF
XInnerRing iovss GuardRing_P17368W3836HFF
DDGATE iovss gate sky130_fd_pr__diode_pw2nd_05v5 area=1.875e-13 pj=2.0um
RRoff iovss off 2391.0121212121
.ends Clamp_N32N4D
* LevelDown
.subckt LevelDown vdd vss iovdd iovss pad core
Mn_hvinv vss padres padres_n vss sky130_fd_pr__nfet_g5v0d10v5__model l=0.5um w=1.35um
Mp_hvinv vdd padres padres_n vdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.5um w=2.45um
Mn_lvinv core padres_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.46um
Mp_lvinv core padres_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.56um
Xsecondprot iovdd iovss pad padres SecondaryProtection
.ends LevelDown
* GuardRing_N18000W13312HFF
.subckt GuardRing_N18000W13312HFF conn

.ends GuardRing_N18000W13312HFF
* Clamp_P32N0D
.subckt Clamp_P32N0D iovss iovdd pad
Mclamp_g0 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g1 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g2 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g3 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g4 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g5 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g6 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g7 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g8 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g9 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g10 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g11 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g12 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g13 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g14 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g15 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g16 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g17 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g18 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g19 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g20 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g21 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g22 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g23 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g24 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g25 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g26 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g27 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g28 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g29 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g30 iovdd off pad iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
Mclamp_g31 pad off iovdd iovdd sky130_fd_pr__pfet_g5v0d10v5__model l=0.6um w=38.2um
XOuterRing iovss GuardRing_P18000W8728HFF
XInnerRing iovdd GuardRing_N17368W8096HTF
RRoff iovdd off 5502.103030303
.ends Clamp_P32N0D
* Clamp_N32N0D
.subckt Clamp_N32N0D iovss iovdd pad
Mclamp_g0 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g1 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g2 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g3 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g4 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g5 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g6 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g7 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g8 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g9 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g10 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g11 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g12 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g13 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g14 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g15 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g16 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g17 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g18 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g19 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g20 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g21 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g22 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g23 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g24 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g25 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g26 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g27 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g28 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g29 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g30 iovss off pad iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
Mclamp_g31 pad off iovss iovss sky130_fd_pr__nfet_g5v0d10v5__model l=0.6um w=16.9um
XOuterRing iovdd GuardRing_N18000W4468HFF
XInnerRing iovss GuardRing_P17368W3836HFF
RRoff iovss off 2391.0121212121
.ends Clamp_N32N0D
* Pad_15800W12000H
.subckt Pad_15800W12000H pad

.ends Pad_15800W12000H
* IOPadAnalog
.subckt IOPadAnalog vss vdd iovss iovdd pad padres
Xpad pad Pad_15800W12000H
Xnclamp iovss iovdd pad Clamp_N12N0D
Xpclamp iovss iovdd pad Clamp_P12N0D
Xsecondprot iovdd iovss pad padres SecondaryProtection
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadAnalog
* IOPadIOVdd
.subckt IOPadIOVdd vss vdd iovss iovdd
Xpad iovdd Pad_15800W12000H
Xnclamp iovss iovdd iovdd ngate Clamp_N32N32D
Xrcres iovdd res_cap RCClampResistor
Xrcinv iovdd iovss res_cap ngate RCClampInverter
Xpad_guard iovss GuardRing_N18000W13312HFF
.ends IOPadIOVdd
* IOPadIOVss
.subckt IOPadIOVss vss vdd iovss iovdd
Xpad iovss Pad_15800W12000H
Xnclamp iovss iovdd iovss Clamp_N32N0D
Xpclamp iovss iovdd iovss Clamp_P32N0D
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadIOVss
* IOPadInOut
.subckt IOPadInOut vss vdd iovss iovdd p2c c2p c2p_en pad
Xpad pad Pad_15800W12000H
Xnclamp iovss iovdd pad ngate Clamp_N32N4D
Xpclamp iovss iovdd pad pgate Clamp_P32N4D
Xgatedec vdd vss iovdd c2p c2p_en ngate pgate GateDecode
Xleveldown vdd vss iovdd iovss pad p2c LevelDown
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadInOut
* IOPadTriOut
.subckt IOPadTriOut vss vdd iovss iovdd c2p c2p_en pad
Xpad pad Pad_15800W12000H
Xnclamp iovss iovdd pad ngate Clamp_N32N4D
Xpclamp iovss iovdd pad pgate Clamp_P32N4D
Xgatedec vdd vss iovdd c2p c2p_en ngate pgate GateDecode
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadTriOut
* IOPadOut
.subckt IOPadOut vss vdd iovss iovdd c2p pad
Xpad pad Pad_15800W12000H
Xnclamp iovss iovdd pad ngate Clamp_N32N4D
Xpclamp iovss iovdd pad pgate Clamp_P32N4D
Xgatelu vdd vss iovdd c2p ngate pgate GateLevelUpInv
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadOut
* IOPadIn
.subckt IOPadIn vss vdd iovss iovdd p2c pad
Xpad pad Pad_15800W12000H
Xnclamp iovss iovdd pad Clamp_N32N0D
Xpclamp iovss iovdd pad Clamp_P32N0D
Xleveldown vdd vss iovdd iovss pad p2c LevelDown
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadIn
* IOPadVdd
.subckt IOPadVdd vss vdd iovss iovdd
Xpad vdd Pad_15800W12000H
Xnclamp iovss iovdd vdd Clamp_N32N0D
Xpclamp iovss iovdd vdd Clamp_P32N0D
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadVdd
* IOPadVss
.subckt IOPadVss vss vdd iovss iovdd
Xpad vss Pad_15800W12000H
Xnclamp iovss iovdd vss Clamp_N32N0D
Xpclamp iovss iovdd vss Clamp_P32N0D
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadVss
* Filler10000
.subckt Filler10000 vss vdd iovss iovdd

.ends Filler10000
* Filler4000
.subckt Filler4000 vss vdd iovss iovdd

.ends Filler4000
* Filler2000
.subckt Filler2000 vss vdd iovss iovdd

.ends Filler2000
* Filler1000
.subckt Filler1000 vss vdd iovss iovdd

.ends Filler1000
* Filler400
.subckt Filler400 vss vdd iovss iovdd

.ends Filler400
* Filler200
.subckt Filler200 vss vdd iovss iovdd

.ends Filler200
* Corner
.subckt Corner vss vdd iovss iovdd

.ends Corner
* Gallery
.subckt Gallery vdd vss iovdd iopadin_pad iopadout_pad iopadtriout_pad iopadinout_pad iopadin_p2c iopadinout_p2c iopadout_c2p iopadtriout_c2p iopadinout_c2p iopadtriout_c2p_en iopadinout_c2p_en ana_out ana_outres
Xcorner vss vdd vss iovdd Corner
Xfiller200 vss vdd vss iovdd Filler200
Xfiller400 vss vdd vss iovdd Filler400
Xfiller1000 vss vdd vss iovdd Filler1000
Xfiller2000 vss vdd vss iovdd Filler2000
Xfiller4000 vss vdd vss iovdd Filler4000
Xfiller10000 vss vdd vss iovdd Filler10000
Xiopadvss vss vdd vss iovdd IOPadVss
Xiopadvdd vss vdd vss iovdd IOPadVdd
Xiopadin vss vdd vss iovdd iopadin_p2c iopadin_pad IOPadIn
Xiopadout vss vdd vss iovdd iopadout_c2p iopadout_pad IOPadOut
Xiopadtriout vss vdd vss iovdd iopadtriout_c2p iopadtriout_c2p_en iopadtriout_pad IOPadTriOut
Xiopadinout vss vdd vss iovdd iopadinout_p2c iopadinout_c2p iopadinout_c2p_en iopadinout_pad IOPadInOut
Xiopadiovss vss vdd vss iovdd IOPadIOVss
Xiopadiovdd vss vdd vss iovdd IOPadIOVdd
Xiopadanalog vss vdd vss iovdd ana_out ana_outres IOPadAnalog
Xcorner2 vss vdd vss iovdd Corner
.ends Gallery
