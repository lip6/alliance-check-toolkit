* Spice description of nao2o22_x1
* Spice driver version 486584091
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:55

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt nao2o22_x1 8 4 6 5 9 2 7 
* NET 2 = vdd
* NET 4 = i1
* NET 5 = i3
* NET 6 = i2
* NET 7 = vss
* NET 8 = i0
* NET 9 = nq
Mtr_00008 3 8 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.91U AS=0.9384P AD=0.9384P PS=8.3U PD=8.3U 
Mtr_00007 2 6 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.91U AS=0.9384P AD=0.9384P PS=8.3U PD=8.3U 
Mtr_00006 1 5 9 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.91U AS=0.9384P AD=0.9384P PS=8.3U PD=8.3U 
Mtr_00005 9 4 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.91U AS=0.9384P AD=0.9384P PS=8.3U PD=8.3U 
Mtr_00004 9 8 10 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 10 4 9 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 7 5 10 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 10 6 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C9 2 7 1.62372e-15
C7 4 7 1.777e-15
C6 5 7 2.07758e-15
C5 6 7 2.02358e-15
C4 7 7 1.57223e-15
C3 8 7 1.73781e-15
C2 9 7 2.24293e-15
C1 10 7 8.84127e-16
.ends nao2o22_x1

