* Spice description of na4_x1
* Spice driver version 963464987
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:52

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt na4_x1 6 7 3 2 5 1 10 
* NET 1 = vdd
* NET 2 = i3
* NET 3 = i2
* NET 5 = nq
* NET 6 = i0
* NET 7 = i1
* NET 10 = vss
Mtr_00008 1 2 5 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00007 1 7 5 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00006 5 6 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00005 5 3 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00004 5 2 4 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 4 3 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 8 6 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 9 7 8 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C10 1 10 1.96957e-15
C9 2 10 1.80781e-15
C8 3 10 2.10271e-15
C6 5 10 2.7235e-15
C5 6 10 2.09358e-15
C4 7 10 2.10271e-15
C1 10 10 1.66309e-15
.ends na4_x1

