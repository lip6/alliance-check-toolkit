* GuardRing_P632W1550HFF
* GuardRing_P632W1550HFF
.subckt GuardRing_P632W1550HFF conn

.ends GuardRing_P632W1550HFF
