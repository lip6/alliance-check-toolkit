-- no model for nor2_x1
