* Spice description of nao22_x1
* Spice driver version -970236133
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:53

* INTERF i0 i1 i2 nq vdd vss 


.subckt nao22_x1 6 5 3 7 2 4 
* NET 2 = vdd
* NET 3 = i2
* NET 4 = vss
* NET 5 = i1
* NET 6 = i0
* NET 7 = nq
Mtr_00006 2 3 7 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 7 5 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00004 1 6 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00003 4 3 8 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00002 8 5 7 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00001 7 6 8 4 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
C7 2 4 1.46971e-15
C6 3 4 2.39212e-15
C5 4 4 1.41822e-15
C4 5 4 1.68915e-15
C3 6 4 1.70741e-15
C2 7 4 2.18063e-15
C1 8 4 4.07001e-16
.ends nao22_x1

