* Spice description of noa2a22_x4
* Spice driver version 1232875291
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:08

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt noa2a22_x4 10 9 6 5 3 2 12 
* NET 2 = vdd
* NET 3 = nq
* NET 5 = i3
* NET 6 = i2
* NET 9 = i1
* NET 10 = i0
* NET 12 = vss
Mtr_00014 3 4 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 2 4 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 2 8 4 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00011 1 9 8 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00010 8 10 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00009 1 6 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00008 2 5 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 3 4 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00006 12 4 3 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 12 8 4 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00004 7 5 8 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00003 8 9 11 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 11 10 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 12 6 7 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C12 1 12 9.1453e-16
C11 2 12 3.98684e-15
C10 3 12 2.15173e-15
C9 4 12 1.77721e-15
C8 5 12 1.95384e-15
C7 6 12 1.86257e-15
C5 8 12 2.6497e-15
C4 9 12 1.83787e-15
C3 10 12 1.55511e-15
C1 12 12 3.82894e-15
.ends noa2a22_x4

