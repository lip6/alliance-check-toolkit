* DP8TRowDecoderDriverPage_2PD8R_wl2
* DP8TWLDrive_30LN100WN30LP200WP_wl2
.subckt DP8TWLDrive_30LN100WN30LP200WP_wl2 vss vdd wl_n wl_drive
Mnmos1 vss wl_n wl_drive vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.5um
Mnmos2 wl_drive wl_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.5um
Mpmos1 vdd wl_n wl_drive vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.0um
Mpmos2 wl_drive wl_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.0um
.ends DP8TWLDrive_30LN100WN30LP200WP_wl2
* DP8TRowDecoderNand3
.subckt DP8TRowDecoderNand3 vss vdd pd[0] pd[1] wl_en wl_n
Mnmos[0] vss pd[0] int[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.65um
Mnmos[1] int[0] pd[1] int[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.65um
Mnmos[2] int[1] wl_en wl_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.65um
Mpmos[0] vdd pd[0] wl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.65um
Mpmos[1] wl_n pd[1] vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.65um
Mpmos[2] vdd wl_en wl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.65um
.ends DP8TRowDecoderNand3
* DP8TRowDecoderDriverPage_2PD8R_wl2
.subckt DP8TRowDecoderDriverPage_2PD8R_wl2 vss vdd pd[0][0] wl[0] pd[0][1] wl[1] pd[0][2] wl[2] pd[0][3] wl[3] pd[0][4] wl[4] pd[0][5] wl[5] pd[0][6] wl[6] pd[0][7] wl[7] pd[1] wl_en
Xnand3[0] vss vdd pd[0][0] pd[1] wl_en wl_n[0] DP8TRowDecoderNand3
Xnand3[1] vss vdd pd[0][1] pd[1] wl_en wl_n[1] DP8TRowDecoderNand3
Xnand3[2] vss vdd pd[0][2] pd[1] wl_en wl_n[2] DP8TRowDecoderNand3
Xnand3[3] vss vdd pd[0][3] pd[1] wl_en wl_n[3] DP8TRowDecoderNand3
Xnand3[4] vss vdd pd[0][4] pd[1] wl_en wl_n[4] DP8TRowDecoderNand3
Xnand3[5] vss vdd pd[0][5] pd[1] wl_en wl_n[5] DP8TRowDecoderNand3
Xnand3[6] vss vdd pd[0][6] pd[1] wl_en wl_n[6] DP8TRowDecoderNand3
Xnand3[7] vss vdd pd[0][7] pd[1] wl_en wl_n[7] DP8TRowDecoderNand3
Xdrive[0] vss vdd wl_n[0] wl[0] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[1] vss vdd wl_n[1] wl[1] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[2] vss vdd wl_n[2] wl[2] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[3] vss vdd wl_n[3] wl[3] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[4] vss vdd wl_n[4] wl[4] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[5] vss vdd wl_n[5] wl[5] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[6] vss vdd wl_n[6] wl[6] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[7] vss vdd wl_n[7] wl[7] DP8TWLDrive_30LN100WN30LP200WP_wl2
.ends DP8TRowDecoderDriverPage_2PD8R_wl2
