*
* 

*****************

.TEMP 25

******************
* BSIM4 transistor model parameters for ngspice
*.lib /users/soft/analogdesign/scalable/techno/sky130_models_20220217/C4M.Sky130_all_lib.spice logic_tt 

*******************************
*Simulation conditions

Vground evss 0 0
Vsupply evdd 0 DC 1.8
*gfoncd evdd 0 evdd 0 1.0e-15

******************
* circuit model
* include circuit netlist
.include picorv32_cts_r.spi
*****************

*****************
* Circuit Instantiation
*.subckt inv_x2 vdd vss i nq


Xc 29279 59920 59919 59918 59917 59916 59915 59914 59913 59900 59899 59896 59898 59885 59884 59872 59870 59869 59868 59865 59867 59851 59850 59837 59836 59833 59826 59818 59815 59814 59812 59803 59799 59798 59797 59785 59784 59783 59782 59774 59768 59761 59755 59747 59742 59737 59728 59723 59716 59709 59705 59700 59693 59685 59680 59676 59667 59666 59657 59652 59646 59638 59632 59627 59618 7031 91 90 53734 58492 57807 58497 57800 59040 56056 56606 55560 54347 57170 54949 56589 57786 59017 59648 57782 52532 52538 51407 50133 59014 54320 54318 54939 52527 52512 53115 53112 53700 6016 56049 54933 56040 54310 55518 54923 55503 54916 58460 59002 57768 59612 58979 58448 57121 57126 58465 58471 58966 58424 58950 57153 57776 57770 57764 58429 57714 57103 57118 56531 58963 58441 12202 49429 10953 11859 10964 59414 59405 59397 59525 58818 58388 58025 57420 56422 55868 55448 54873 54565 54015 52926 52303 53108 51311 53097 50391 49342 49470 48323 48849 49461 47828 50027 49441 48282 47173 46607 47149 3873 6387 59609 59604 59633 59594 59621 59582 59572 59617 59561 59634 59596 59610 59583 59534 59526 59517 59513 59619 59570 59493 59535 59481 59476 59468 59460 59456 59549 59444 59436 59432 59558 59416 13415 12950 12205 11579 25294 24777 24165 24167 23610 24166 23006 23611 23007 19844 18780 18156 17618 17130 16618 16351 15363 14702 14127 13575 13031 12802 12361 11117 10543 10008 9512 9285 8291 7666 7130 6618 26326 5886 47825 44830 50041 47836 47391 52461 59250 58668 58098 57569 56795 56269 55761 55168 54606 54123 53373 52750 52169 51650 51036 50518 49767 49166 48556 48121 47596 47103 46336 45750 27360 26907 26187 25681 26480 25426 25436 23890 26494 24907 25946 24866 20500 20012 19217 18603 18008 17527 17001 16516 15788 16010 16700 16688 3011 28723 607 606 285 284 605 283 281 282 271 270 260 259 257 567 566 565 243 242 241 551 545 225 216 215 214 213 212 210 201 200 199 198 188 502 178 177 4827 10001 evdd evss picorv32_cts_r 
.end

